PK
     �8�ZuaKbH bH    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_7"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_4"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_1","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_1"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5":["pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_10"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6":["pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_0"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7":["pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_1"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8":["pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_2"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_5"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14":[],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15":["pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_4"],"pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0":[],"pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1":[],"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13"],"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1"],"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"],"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12"],"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2"],"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7"],"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11"],"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8"],"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3"],"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"],"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6"],"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10"],"pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15"],"pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"],"pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9"],"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_0":["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_14"],"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_1":["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_13"],"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_2":["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_12"],"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_3":["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_11"],"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_4":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3"],"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_5":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_3":[],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_4":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_5":[],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_6":[],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_7":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_9":[],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_10":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_11":["pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_3"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_12":["pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_2"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_13":["pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_1"],"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_14":["pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_0"],"pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"],"pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"]},"pin_to_color":{"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0":"#ff0000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1":"#ff0000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2":"#ff0000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3":"#ff0000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4":"#ff0000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5":"#98FF52","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6":"#0300b3","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7":"#0cdf2f","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8":"#b6c11a","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9":"#000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10":"#000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11":"#000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12":"#000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13":"#000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14":"#000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15":"#01FFFE","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0":"#000000","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1":"#000000","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0":"#000000","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1":"#ff0000","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2":"#98FF52","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0":"#000000","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1":"#ff0000","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2":"#0cdf2f","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0":"#000000","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1":"#b6c11a","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2":"#ff0000","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0":"#ff0000","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1":"#0300b3","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2":"#000000","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0":"#01FFFE","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_1":"#ff0000","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2":"#000000","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_0":"#968AE8","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_1":"#FF74A3","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_2":"#FF029D","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_3":"#683D3B","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_4":"#ff0000","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_5":"#000000","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_0":"#0300b3","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_1":"#0cdf2f","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_3":"#000000","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_2":"#b6c11a","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_4":"#01FFFE","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_5":"#000000","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_6":"#000000","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_7":"#ff0000","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8":"#000000","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_9":"#000000","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_10":"#98FF52","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_11":"#683D3B","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_12":"#FF029D","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_13":"#FF74A3","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_14":"#968AE8","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0":"#98FF52","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_1":"#ff0000"},"pin_to_state":{"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15":"neutral","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0":"neutral","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1":"neutral","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0":"neutral","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1":"neutral","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2":"neutral","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0":"neutral","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1":"neutral","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2":"neutral","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0":"neutral","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1":"neutral","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2":"neutral","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0":"neutral","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1":"neutral","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2":"neutral","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0":"neutral","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_1":"neutral","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2":"neutral","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_0":"neutral","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_1":"neutral","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_2":"neutral","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_3":"neutral","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_4":"neutral","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_5":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_0":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_1":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_3":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_2":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_4":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_5":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_6":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_7":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_9":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_10":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_11":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_12":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_13":"neutral","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_14":"neutral","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0":"neutral","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_1":"neutral"},"next_color_idx":22,"wires_placed_in_order":[["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_23","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_22"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_35"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21"],["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6"],["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_bd8b6d2d-60e6-4b66-abf0-62afb810491d_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_8"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_7"],["pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_4"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_2"],["pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_7","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_8"],["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_7"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8"],["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_12","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_2"],["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_11","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_3"],["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_13","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_1"],["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_14","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_4"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_5"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_1"],["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0"],["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0"],["pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_4"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_10"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_0"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_23","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_22"]]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_35"]]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21"]]],[[],[["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20"]]],[[["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21"]],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21"]],[]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20"]],[]],[[["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_22","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_23"]],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_35"]],[]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"]]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"]],[]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"]]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6"]]],[[],[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_bd8b6d2d-60e6-4b66-abf0-62afb810491d_0"]]],[[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_bd8b6d2d-60e6-4b66-abf0-62afb810491d_0"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2"]]],[[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]],[]],[[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]]],[[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2"]]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9"]],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0"]],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6"]],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7"]],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8"]],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_8"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_7"]]],[[],[["pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_4"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_2"]]],[[],[["pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_7","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_8"]]],[[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_0"]],[]],[[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_1"]],[]],[[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_2"]],[]],[[["pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_4"]],[]],[[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_7"],["pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_7","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_8"]],[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2"]]],[[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_5f38e467-a28b-4220-b03f-542b6f72ddb0_8"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_7"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8"]]],[[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8"]],[]],[[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8"]]],[[],[["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_12","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_2"]]],[[],[["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_11","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_3"]]],[[],[["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_13","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_1"]]],[[],[["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_14","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_4"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_5"]]],[[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_1"]]],[[],[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0"]]],[[],[]],[[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"]],[]],[[],[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"]]],[[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"]],[]],[[["pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0"]]],[[],[["pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_4"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_10"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_2"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_0"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0":"0000000000000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1":"0000000000000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2":"0000000000000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3":"0000000000000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4":"0000000000000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5":"0000000000000005","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6":"0000000000000004","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7":"0000000000000003","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8":"0000000000000002","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9":"0000000000000001","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10":"0000000000000001","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11":"0000000000000001","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12":"0000000000000001","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13":"0000000000000001","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14":"_","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15":"0000000000000010","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0":"_","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1":"_","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0":"0000000000000001","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1":"0000000000000000","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2":"0000000000000005","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0":"0000000000000001","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1":"0000000000000000","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2":"0000000000000003","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0":"0000000000000001","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1":"0000000000000002","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2":"0000000000000000","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0":"0000000000000000","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1":"0000000000000004","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2":"0000000000000001","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0":"0000000000000010","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_1":"0000000000000000","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2":"0000000000000001","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_0":"0000000000000009","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_1":"0000000000000008","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_2":"0000000000000006","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_3":"0000000000000007","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_4":"0000000000000000","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_5":"0000000000000001","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_0":"0000000000000004","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_1":"0000000000000003","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_3":"_","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_2":"0000000000000002","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_4":"0000000000000010","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_5":"_","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_6":"_","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_7":"0000000000000000","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8":"0000000000000001","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_9":"_","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_10":"0000000000000005","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_11":"0000000000000007","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_12":"0000000000000006","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_13":"0000000000000008","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_14":"0000000000000009","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0":"0000000000000005","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_1":"0000000000000000"},"component_id_to_pins":{"413adb9e-60b4-4310-bd72-e4e11d56ccb2":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"1cb3a49d-dc66-4fa6-8d47-aea3068df0b4":["0","1"],"7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c":["0","1","2"],"6709695f-c694-4d3b-8888-654e702eb44c":["0","1","2"],"ff0891dd-490d-4f7f-b028-abe315436194":["0","1","2"],"9160c2c5-ef89-4fab-911c-be70a3060d8a":["0","1","2"],"686232c8-bdc9-4b03-9791-f090cd6c7e85":[],"470753c0-2a44-41d6-b577-b515fa83a749":[],"17669cf5-00f7-487e-af61-6dc7cec32cac":[],"78042b3a-f2f8-4275-8b35-53f2a17714ef":[],"2efedb33-0a07-490d-b599-10accff66be5":["0","1","2"],"0cfff15f-c777-4f91-842e-b8dc1b9acc4a":["0","1","2","3","4","5"],"b9f30b96-c79a-461e-b5af-a20a819f12ff":["0","1","3","2","4","5","6","7","8","9","10","11","12","13","14"],"d5a8db9d-834a-4142-867c-6467eef2692c":[],"c7f861b9-9e3f-47e9-8093-8c86ac31e125":[],"05b878bc-14bf-43ae-b053-88be25e3fc2e":["0","1"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_4","pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_7","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2","pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_1"],"0000000000000002":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_2"],"0000000000000003":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_1"],"0000000000000004":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_0"],"0000000000000005":["pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_10"],"0000000000000001":["pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_5"],"0000000000000006":["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_12","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_2"],"0000000000000007":["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_11","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_3"],"0000000000000008":["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_13","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_1"],"0000000000000009":["pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_14","pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_0"],"0000000000000010":["pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15","pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_4"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000001":"Net 1","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000009":"Net 9","0000000000000010":"Net 10"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"4.7","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[528.299914926406,239.30827804023798],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"1cb3a49d-dc66-4fa6-8d47-aea3068df0b4","orientation":"up","circleData":[[512.5,260.00000000000006],[542.5,290.00000000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[318.2035,528.6544999999999],"typeId":"6500d8ea-11fe-42e2-8a9f-99be354012a7","componentVersion":1,"instanceId":"7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c","orientation":"up","circleData":[[212.5,560],[222.44650000000001,567.7579999999998],[240.05050000000006,567.1609999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[43.31500000000004,434.6300000000002],"typeId":"6d0c07c0-db0e-4413-b9a4-ee378c2ed587","componentVersion":1,"instanceId":"ff0891dd-490d-4f7f-b028-abe315436194","orientation":"up","circleData":[[-87.50000000000001,485],[-81.25249999999996,496.5335000000001],[-73.08349999999997,506.8655000000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Turbidity sensor","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[57.96696427243663,531.1244549982175],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"686232c8-bdc9-4b03-9791-f090cd6c7e85","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Temperature Sensor","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[292.2231314606828,614.5459012322258],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"470753c0-2a44-41d6-b577-b515fa83a749","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"PH SENSOR","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[550.8560026663338,727.7651803249732],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"17669cf5-00f7-487e-af61-6dc7cec32cac","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[570.165334,616.4889995],"typeId":"8e0ee0b2-778d-4065-bf79-38edea29856f","componentVersion":1,"instanceId":"6709695f-c694-4d3b-8888-654e702eb44c","orientation":"up","circleData":[[497.5,665],[507.055,672.077],[517.3165,677.7395]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[801.3969999999999,646.5035],"typeId":"1cec4e8a-72c2-4b6a-9a5c-b6be0dc427d1","componentVersion":1,"instanceId":"9160c2c5-ef89-4fab-911c-be70a3060d8a","orientation":"up","circleData":[[812.5,695],[820.9989999999998,687.0725],[829.7424999999998,679.31]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"TDS SENSOR","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[772.1681606443491,794.1359304792926],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"78042b3a-f2f8-4275-8b35-53f2a17714ef","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1198.4483395000002,676.7642555000003],"typeId":"fdbf9524-da67-4179-8c49-1739e12a7ba1","componentVersion":2,"instanceId":"2efedb33-0a07-490d-b599-10accff66be5","orientation":"down","circleData":[[1037.5,650],[1037.5,635],[1037.5,620]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1257.0931135,507.5196440000001],"typeId":"86f6860e-1b0a-4bec-9c42-62e574033eb9","componentVersion":1,"instanceId":"0cfff15f-c777-4f91-842e-b8dc1b9acc4a","orientation":"down","circleData":[[1157.5,470],[1157.5,485],[1157.5,500],[1157.5,515],[1157.5,530],[1157.5,545]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1074.185311,146.5564009999999],"typeId":"da94d5db-27d7-4cba-87e7-6294921d661c","componentVersion":3,"instanceId":"b9f30b96-c79a-461e-b5af-a20a819f12ff","orientation":"up","circleData":[[947.5,200],[947.5,214.99999999999994],[947.5,240.4999999999999],[947.5,226.99999999999994],[962.5,226.99999999999994],[962.5,214.99999999999994],[962.5,200],[947.5,132.5],[947.5,162.5],[947.5,117.5],[962.5,95],[1204.15,100.55000000000001],[1203.4,113.14999999999998],[1202.5,87.5],[1187.5,176]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"SD CARD MODULE","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1259.3707464064173,599.8893023249628],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"d5a8db9d-834a-4142-867c-6467eef2692c","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"PRESSURE SENSOR","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1256.9194702265036,770.2267710836668],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"c7f861b9-9e3f-47e9-8093-8c86ac31e125","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[511.8908200000001,204.4938005],"typeId":"a634ff83-abbb-414f-80bc-066b6f1a8bb9","componentVersion":1,"instanceId":"413adb9e-60b4-4310-bd72-e4e11d56ccb2","orientation":"up","circleData":[[602.5,215.00000000000003],[602.3500000000001,236.0000000000001],[601.9000000000001,259.33399999999995],[600.25,282.66650000000004],[603.6670000000001,306.0005],[532.1335000000001,306.0005],[509.16700000000014,306.0005],[487.0000000000001,306.0005],[464.83450000000005,307.1675],[602.5,143.834],[603.6670000000001,119.33449999999999],[602.5,98.33449999999999],[602.5,77.33449999999999],[601.3345000000002,52.833500000000015],[533.6671585000001,283.83383000000003],[580.3338265000001,304.83383000000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"4.7","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[504.9999999999998,245],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"05b878bc-14bf-43ae-b053-88be25e3fc2e","orientation":"up","circleData":[[467.49999999999994,245],[542.5,245]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-108.76672","left":"-101.68500","width":"1487.83881","height":"931.40265","x":"-101.68500","y":"-108.76672"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_215.0000000000\\\",\\\"602.5000000000_236.0000000000\\\",\\\"602.3500000000_236.0000000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.3500000000_236.0000000000\\\",\\\"602.5000000000_236.0000000000\\\",\\\"602.5000000000_259.3340000000\\\",\\\"601.9000000000_259.3340000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"601.9000000000_259.3340000000\\\",\\\"602.5000000000_259.3340000000\\\",\\\"602.5000000000_282.5000000000\\\",\\\"600.2500000000_282.5000000000\\\",\\\"600.2500000000_282.6665000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"600.2500000000_282.6665000000\\\",\\\"602.5000000000_282.6665000000\\\",\\\"602.5000000000_305.0000000000\\\",\\\"603.6670000000_305.0000000000\\\",\\\"603.6670000000_306.0005000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"endPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"rawEndPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.3500000000_236.0000000000\\\",\\\"580.0000000000_236.0000000000\\\",\\\"580.0000000000_170.0000000000\\\",\\\"227.5000000000_170.0000000000\\\",\\\"227.5000000000_567.7580000000\\\",\\\"222.4465000000_567.7580000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"endPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"rawEndPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"601.9000000000_259.3340000000\\\",\\\"572.5000000000_259.3340000000\\\",\\\"572.5000000000_177.5000000000\\\",\\\"445.0000000000_177.5000000000\\\",\\\"445.0000000000_680.0000000000\\\",\\\"507.0550000000_680.0000000000\\\",\\\"507.0550000000_672.0770000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"endPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"rawEndPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"600.2500000000_282.6665000000\\\",\\\"625.0000000000_282.6665000000\\\",\\\"625.0000000000_155.0000000000\\\",\\\"-117.5000000000_155.0000000000\\\",\\\"-117.5000000000_506.8655000000\\\",\\\"-73.0835000000_506.8655000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"endPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"rawEndPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"603.6670000000_306.0005000000\\\",\\\"655.0000000000_306.0005000000\\\",\\\"655.0000000000_755.0000000000\\\",\\\"812.5000000000_755.0000000000\\\",\\\"812.5000000000_695.0000000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_1\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"rawStartPinId\":\"pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_1\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1037.5000000000_635.0000000000\\\",\\\"992.5000000000_635.0000000000\\\",\\\"992.5000000000_462.5000000000\\\",\\\"603.6670000000_462.5000000000\\\",\\\"603.6670000000_306.0005000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_7\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_215.0000000000\\\",\\\"767.5000000000_215.0000000000\\\",\\\"767.5000000000_132.5000000000\\\",\\\"947.5000000000_132.5000000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_4\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"rawStartPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_4\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_530.0000000000\\\",\\\"752.5000000000_530.0000000000\\\",\\\"752.5000000000_282.6665000000\\\",\\\"600.2500000000_282.6665000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_1\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"rawStartPinId\":\"pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_1\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.5000000000_245.0000000000\\\",\\\"722.5000000000_245.0000000000\\\",\\\"722.5000000000_395.0000000000\\\",\\\"603.6670000000_395.0000000000\\\",\\\"603.6670000000_306.0005000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"603.6670000000_119.3345000000\\\",\\\"603.6670000000_117.5000000000\\\",\\\"602.5000000000_117.5000000000\\\",\\\"602.5000000000_143.8340000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"603.6670000000_119.3345000000\\\",\\\"602.5000000000_119.3345000000\\\",\\\"602.5000000000_98.3345000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_98.3345000000\\\",\\\"602.5000000000_77.3345000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_77.3345000000\\\",\\\"602.5000000000_52.8335000000\\\",\\\"601.3345000000_52.8335000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13\",\"endPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13\",\"rawEndPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"601.3345000000_52.8335000000\\\",\\\"601.3345000000_5.0000000000\\\",\\\"182.5000000000_5.0000000000\\\",\\\"182.5000000000_560.0000000000\\\",\\\"212.5000000000_560.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"endPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"rawEndPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_77.3345000000\\\",\\\"602.5000000000_80.0000000000\\\",\\\"302.5000000000_80.0000000000\\\",\\\"302.5000000000_447.5000000000\\\",\\\"430.0000000000_447.5000000000\\\",\\\"430.0000000000_665.0000000000\\\",\\\"497.5000000000_665.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"endPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"rawEndPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_98.3345000000\\\",\\\"602.5000000000_95.0000000000\\\",\\\"-102.5000000000_95.0000000000\\\",\\\"-102.5000000000_485.0000000000\\\",\\\"-87.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"endPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"rawEndPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"603.6670000000_119.3345000000\\\",\\\"603.6670000000_125.0000000000\\\",\\\"677.5000000000_125.0000000000\\\",\\\"677.5000000000_740.0000000000\\\",\\\"829.7425000000_740.0000000000\\\",\\\"829.7425000000_679.3100000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9\",\"rawStartPinId\":\"pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_2\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1037.5000000000_620.0000000000\\\",\\\"887.5000000000_620.0000000000\\\",\\\"887.5000000000_395.0000000000\\\",\\\"842.5000000000_395.0000000000\\\",\\\"842.5000000000_170.0000000000\\\",\\\"602.5000000000_170.0000000000\\\",\\\"602.5000000000_143.8340000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"601.3345000000_52.8335000000\\\",\\\"601.3345000000_50.0000000000\\\",\\\"947.5000000000_50.0000000000\\\",\\\"947.5000000000_162.5000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_5\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9\",\"rawStartPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_5\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_545.0000000000\\\",\\\"730.0000000000_545.0000000000\\\",\\\"730.0000000000_143.8340000000\\\",\\\"602.5000000000_143.8340000000\\\"]}\"}","{\"color\":\"#b6c11a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8\",\"endPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8\",\"rawEndPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"464.8345000000_307.1675000000\\\",\\\"464.8345000000_267.5000000000\\\",\\\"-80.0000000000_267.5000000000\\\",\\\"-80.0000000000_496.5335000000\\\",\\\"-81.2525000000_496.5335000000\\\"]}\"}","{\"color\":\"#b6c11a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"464.8345000000_307.1675000000\\\",\\\"464.8345000000_425.0000000000\\\",\\\"782.5000000000_425.0000000000\\\",\\\"782.5000000000_227.0000000000\\\",\\\"947.5000000000_227.0000000000\\\"]}\"}","{\"color\":\"#0cdf2f\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7\",\"endPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7\",\"rawEndPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"487.0000000000_306.0005000000\\\",\\\"487.0000000000_290.0000000000\\\",\\\"452.5000000000_290.0000000000\\\",\\\"452.5000000000_695.0000000000\\\",\\\"517.3165000000_695.0000000000\\\",\\\"517.3165000000_677.7395000000\\\"]}\"}","{\"color\":\"#0cdf2f\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"487.0000000000_306.0005000000\\\",\\\"487.0000000000_402.5000000000\\\",\\\"767.5000000000_402.5000000000\\\",\\\"767.5000000000_215.0000000000\\\",\\\"947.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#0300b3\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6\",\"endPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6\",\"rawEndPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"509.1670000000_306.0005000000\\\",\\\"509.1670000000_410.0000000000\\\",\\\"632.5000000000_410.0000000000\\\",\\\"632.5000000000_770.0000000000\\\",\\\"820.9990000000_770.0000000000\\\",\\\"820.9990000000_687.0725000000\\\"]}\"}","{\"color\":\"#0300b3\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_0\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"509.1670000000_306.0005000000\\\",\\\"509.1670000000_477.5000000000\\\",\\\"820.0000000000_477.5000000000\\\",\\\"820.0000000000_200.0000000000\\\",\\\"947.5000000000_200.0000000000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"endPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"rawEndPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"532.1335000000_306.0005000000\\\",\\\"532.1335000000_282.5000000000\\\",\\\"242.5000000000_282.5000000000\\\",\\\"242.5000000000_567.1610000000\\\",\\\"240.0505000000_567.1610000000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"rawStartPinId\":\"pin-type-component_05b878bc-14bf-43ae-b053-88be25e3fc2e_0\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"467.5000000000_245.0000000000\\\",\\\"467.5000000000_260.0000000000\\\",\\\"532.1335000000_260.0000000000\\\",\\\"532.1335000000_306.0005000000\\\"]}\"}","{\"color\":\"#98FF52\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_10\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"532.1335000000_306.0005000000\\\",\\\"532.1335000000_447.5000000000\\\",\\\"797.5000000000_447.5000000000\\\",\\\"797.5000000000_95.0000000000\\\",\\\"962.5000000000_95.0000000000\\\"]}\"}","{\"color\":\"#FF029D\",\"startPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_2\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_12\",\"rawStartPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_2\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_500.0000000000\\\",\\\"1127.5000000000_500.0000000000\\\",\\\"1127.5000000000_417.5000000000\\\",\\\"1367.5000000000_417.5000000000\\\",\\\"1367.5000000000_113.1500000000\\\",\\\"1203.4000000000_113.1500000000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_3\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_11\",\"rawStartPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_3\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_515.0000000000\\\",\\\"1112.5000000000_515.0000000000\\\",\\\"1112.5000000000_402.5000000000\\\",\\\"1345.0000000000_402.5000000000\\\",\\\"1345.0000000000_100.5500000000\\\",\\\"1204.1500000000_100.5500000000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_1\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_13\",\"rawStartPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_1\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_13\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_485.0000000000\\\",\\\"1090.0000000000_485.0000000000\\\",\\\"1090.0000000000_387.5000000000\\\",\\\"1330.0000000000_387.5000000000\\\",\\\"1330.0000000000_87.5000000000\\\",\\\"1202.5000000000_87.5000000000\\\"]}\"}","{\"color\":\"#968AE8\",\"startPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_0\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_14\",\"rawStartPinId\":\"pin-type-component_0cfff15f-c777-4f91-842e-b8dc1b9acc4a_0\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_14\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_470.0000000000\\\",\\\"1075.0000000000_470.0000000000\\\",\\\"1075.0000000000_372.5000000000\\\",\\\"1285.0000000000_372.5000000000\\\",\\\"1285.0000000000_176.0000000000\\\",\\\"1187.5000000000_176.0000000000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15\",\"rawStartPinId\":\"pin-type-component_2efedb33-0a07-490d-b599-10accff66be5_0\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1037.5000000000_650.0000000000\\\",\\\"1037.5000000000_507.5000000000\\\",\\\"580.3338265000_507.5000000000\\\",\\\"580.3338265000_304.8338300000\\\"]}\"}","{\"color\":\"#01FFFE\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15\",\"endPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_4\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15\",\"rawEndPinId\":\"pin-type-component_b9f30b96-c79a-461e-b5af-a20a819f12ff_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"580.3338265000_304.8338300000\\\",\\\"580.3338265000_305.0000000000\\\",\\\"962.5000000000_305.0000000000\\\",\\\"962.5000000000_227.0000000000\\\"]}\"}"],"projectDescription":""}PK
     �8�Z               jsons/PK
     �8�Z�֎�?  �?     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"TEMP","category":["User Defined"],"id":"6500d8ea-11fe-42e2-8a9f-99be354012a7","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"49baae61-cb81-429b-96a1-6cfb8f124b59.png","iconPic":"9c69fbd4-c376-47ca-8b4c-793dd402431a.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"15.00000","numDisplayRows":"15.00000","pins":[{"uniquePinIdString":"0","positionMil":"45.31000,541.03000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"111.62000,489.31000","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"228.98000,493.29000","isAnchorPin":false,"label":"A0"}],"pinType":"wired"},"properties":[]},{"subtypeName":"TURBI","category":["User Defined"],"id":"6d0c07c0-db0e-4413-b9a4-ee378c2ed587","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"a1588c66-a70c-44df-b30c-55fdbd854069.png","iconPic":"2dd92824-eee5-446a-82e5-cb3be823b6e8.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"18.00000","numDisplayRows":"15.00000","pins":[{"uniquePinIdString":"0","positionMil":"27.90000,414.20000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"69.55000,337.31000","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"2","positionMil":"124.01000,268.43000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"PH","category":["User Defined"],"id":"8e0ee0b2-778d-4065-bf79-38edea29856f","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"256658b1-ffe9-46c3-9f0b-70052a8fe00d.png","iconPic":"d18021d8-4522-4af4-a3c6-358ee97fa8ad.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"18.00000","numDisplayRows":"15.00000","pins":[{"uniquePinIdString":"0","positionMil":"415.56444,426.59333","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"479.26444,379.41333","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"547.67444,341.66333","isAnchorPin":false,"label":"A1"}],"pinType":"wired"},"properties":[]},{"subtypeName":"TDS","category":["User Defined"],"id":"1cec4e8a-72c2-4b6a-9a5c-b6be0dc427d1","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"a05d3615-68b8-4f26-98d6-1aedf7f6d878.png","iconPic":"b75f5fea-d559-4623-b1ce-f8cd504066c2.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"18.00000","numDisplayRows":"15.00000","pins":[{"uniquePinIdString":"0","positionMil":"974.02000,426.69000","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"1030.68000,479.54000","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"2","positionMil":"1088.97000,531.29000","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Gravity: Analog Water Pressure Sensor","category":["User Defined"],"id":"fdbf9524-da67-4179-8c49-1739e12a7ba1","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"00f35920-432a-4227-a0de-f9ff33566dcd.png","iconPic":"fce5a045-7211-4fa3-86b3-f57a3d8041ae.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"21.66377","numDisplayRows":"8.51543","pins":[{"uniquePinIdString":"0","positionMil":"2156.17743,247.34313","isAnchorPin":true,"label":"Signal"},{"uniquePinIdString":"1","positionMil":"2156.17743,147.34313","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"2156.17743,47.34313","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"SDmodule","category":["User Defined"],"id":"86f6860e-1b0a-4bec-9c42-62e574033eb9","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"91777b75-38f2-4118-94bc-a70a6868aa47.jpg","iconPic":"0b0a0ee7-c404-40e4-9217-cd21fece1ba1.jpg","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"15.87476","numDisplayRows":"8.45131","pins":[{"uniquePinIdString":"0","positionMil":"1457.69209,172.43454","isAnchorPin":true,"label":"CS"},{"uniquePinIdString":"1","positionMil":"1457.69209,272.43454","isAnchorPin":false,"label":"SCK"},{"uniquePinIdString":"2","positionMil":"1457.69209,372.43454","isAnchorPin":false,"label":"MOSI"},{"uniquePinIdString":"3","positionMil":"1457.69209,472.43454","isAnchorPin":false,"label":"MISO"},{"uniquePinIdString":"4","positionMil":"1457.69209,572.43454","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"5","positionMil":"1457.69209,672.43454","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Vega Aries IoT","category":["User Defined"],"id":"da94d5db-27d7-4cba-87e7-6294921d661c","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"ed998360-ed4f-472d-a3e6-52adfa722a6d.png","iconPic":"08988072-c7a8-475c-9331-8aa77c72a02a.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"37.49015","numDisplayRows":"32.70975","pins":[{"uniquePinIdString":"0","positionMil":"1029.93876,1279.19684","isAnchorPin":true,"label":"AO"},{"uniquePinIdString":"1","positionMil":"1029.93876,1179.19684","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"3","positionMil":"1029.93876,1009.19684","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"2","positionMil":"1029.93876,1099.19684","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"4","positionMil":"1129.93876,1099.19684","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"5","positionMil":"1129.93876,1179.19684","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"6","positionMil":"1129.93876,1279.19684","isAnchorPin":false,"label":"A6"},{"uniquePinIdString":"7","positionMil":"1029.93876,1729.19684","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"8","positionMil":"1029.93876,1529.19684","isAnchorPin":false,"label":""},{"uniquePinIdString":"9","positionMil":"1029.93876,1829.19684","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"10","positionMil":"1129.93876,1979.19684","isAnchorPin":false,"label":"GPIO30"},{"uniquePinIdString":"11","positionMil":"2740.93876,1942.19684","isAnchorPin":false,"label":"MISO"},{"uniquePinIdString":"12","positionMil":"2735.93876,1858.19684","isAnchorPin":false,"label":"MOSI"},{"uniquePinIdString":"13","positionMil":"2729.93876,2029.19684","isAnchorPin":false,"label":"SCLK"},{"uniquePinIdString":"14","positionMil":"2629.93876,1439.19684","isAnchorPin":false,"label":"GPIO10"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"PCB","category":["User Defined"],"id":"a634ff83-abbb-414f-80bc-066b6f1a8bb9","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"3281a32a-bb08-42cb-a591-9481e2c9eb0d.png","iconPic":"35c60fd9-1fb3-48b8-b3d7-7968b0279531.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"25.12926","numDisplayRows":"23.63459","pins":[{"uniquePinIdString":"0","positionMil":"1860.52420,1111.68817","isAnchorPin":true,"label":"5V"},{"uniquePinIdString":"1","positionMil":"1859.52420,971.68817","isAnchorPin":false,"label":"5V(PH)"},{"uniquePinIdString":"2","positionMil":"1856.52420,816.12817","isAnchorPin":false,"label":"5V TDS"},{"uniquePinIdString":"3","positionMil":"1845.52420,660.57817","isAnchorPin":false,"label":" 5V TURBI"},{"uniquePinIdString":"4","positionMil":"1868.30420,505.01817","isAnchorPin":false,"label":"5V TEMP"},{"uniquePinIdString":"5","positionMil":"1391.41420,505.01817","isAnchorPin":false,"label":"GPIO25  TEMP"},{"uniquePinIdString":"6","positionMil":"1238.30420,505.01817","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"7","positionMil":"1090.52420,505.01817","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"8","positionMil":"942.75420,497.23817","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"9","positionMil":"1860.52420,1586.12817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"10","positionMil":"1868.30420,1749.45817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"11","positionMil":"1860.52420,1889.45817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"12","positionMil":"1860.52420,2029.45817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"13","positionMil":"1852.75420,2192.79817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"14","positionMil":"1401.63859,652.79597","isAnchorPin":false,"label":""},{"uniquePinIdString":"15","positionMil":"1712.74971,512.79597","isAnchorPin":false,"label":""}],"pinType":"wired"},"properties":[]},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"}]}PK
     �8�Z               images/PK
     �8�Z	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     �8�Zd��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     �8�Z�Xw�s� s� /   images/49baae61-cb81-429b-96a1-6cfb8f124b59.png�PNG

   IHDR  7  �   �&�>   	pHYs  �  ��+  ��IDATx��	�Wu/^[�3ӳ�fӾ�F�-ll��1$��;�'���~�|$$�@H�%���9��`0��Ɩ�%[�-K#Y�G�f����ޗ��z�ܪS}�%!�,��O_�{�k�u��=�:��0��`�#0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
LnƼ��8�/����#V���0��$��0��������p8l��i=��j�\N�O>U˲�L&��f��唀���w�a���ٚZ*�[�U8��۶M�F3MS�/�`��iZ�_���J�H��u݂u%�,�0�R]]�����TSSS��ظ�ڵkm F��`0^50�a0�z�)���=2::*
���� ��,�l1��{>֚Jf���ԛf!�8vԶ�0���������R)X�K��S2���zER�!�qJ�RR`+WS��F�4E���pT�<��&e�� *��	�"a�5C/���em���9�P?��@h���_��Gft=�jk�gkkk�`Cܪk�+vǻ�p��u�
��x����`���LC�)���Q}||<8�L6�L��f��xb&�M&�=�XK&�[��fہ���h�L�ֲ�0#�� *�8����n�w�������Ă䅾�P��Ђ��'��jb��E�c����a))%�B-���?UU���S8|����)���>��\$����>2��I���d�&�hji��m�o4�P#�x�b�;���_Ln��
$gΜ	MOO����Լ|�k_k����J$ҭ�T�9�ɴ���i�Jg��k(����D���l+ �@��GW$$H6���B����i��T��|� <Hp�x2����
�߸�C��q�@ ���������M+�E=�����C��X8�
��Ñ�T}c�XC�v�����M/_�Mc�+V�����`�J�1�;4�0j��D�������['��V�%fWX�B�i���B�eY�}-,1`&! z�h�����@xv ������O���b=�KǑ56���
rC��@�>Q�Cǣ�H#��l;tL�d� 7�YBҦ a�?��9p�j|<��|O�@2
��6
��jjkG�u��O~��4/�iYؒm�mM����6m�:��a0�`r�`0~!Ȭ4::	 �Y��o|u����T&ٚL�W�2�E�|��y���5��f� |�iU���x���kT���ք kOp1M�}��ɑA���k>q��˟��Whm���_.%�WP\�Z�Y
8���1��H�����#p��b.�䵌�B#d铓E��q�z��Hx,������o{j�XGg�ضmۆ���&���]]]h�2�u
&7� !�?~<:11����n����R��2�Juer�e�lv)H��|>WcY6��,��A�k�9�B�B������Gh�m\�_���}�����Y�"���j�K��2���b��������&0E+k����cym�~��K��ר��i���� ��dR_g�5���944�9p��X(<[[[s���q�����~��cK�.M����,Y�W����0��AwϩS��'�����[<6:��\.��P0�l�j����,�2�n;�_G^�|kYT���TiDׁFS5A� �$(нm�*8�w�#��1!2��`���Dl�5E����ǭ���ۈk���!SZ�1�GnȜ���x��)����#H95�bC5�d�m-�1r;�W��{0a�*@r�,o���1SG���E��Hh���������t/�w�碥����Ln��!<3S�������Ư~���FF���&W�3���|aY�X\ �6V(�1�Z�PȒ�MB�'�]-_�2�K�3� 7��n�6�Y#��"2"G@ѧ�W#������վ5�KU_TDJ�o�v>b��ST��D��$b��-�)G���]���»�$�
��O�>�����un4���q	��.
�h3��5ΜcNONΞ=3�?��!?�����{�w�����رc�V�B?Mg�+0�a0^'@B3::����MgΜY761�6�N��e�+M�� BS�2�cȵ���cq�f=��p�D!L!�A�5;�.��"�����D�@G���e?ܖ�Ѐ聊���Fv��v���.k^\�u�4�XAl�^I-	�&ks|m�w*�>��JS+�]$`T� ����D��KrBA�zH;&�|�w�Az���}�����`:�������_v�ԩ�b��d49���o�h;���|����˧`���͛�W���c��35�}}}�ӧO�~�K_�z���Ԧd2�
���N�	$����
Uv�E�E�UJh2BJ�"D�K(���D��IJm���vY#��B�G��Ed
�F����i[��G&
2��&7����
.o#�����<°���w<>��p��Ne{}'�{9u�IX�V���lan�����hʲ�B�*���9�D���8��}]Ŝ���Y�=�ۤ�f��n��p6�o�{�RU'���>u��?��Η��k_;���Kǻf��^�5&7�<jg�������x�������GG����ήO���AN6y���
d2��/���
W����\����@PW¡��Q��]�Q��OnP#AA��� ��(���`6)=H�`Wi��=���7cY^�a�#N���H�:�A�JU��U�GF���¿�	�`H��7G��%d=�k^BB��*����>�G+y���Dֆ������������I&�@�5]�vQhy�~ὀU��C�3dR�bmA����Y�U�js�B휑Z
����9y���C�ښ;�;^zꩧN�Ituu��G��Z�c�q�zz��|��ԩ�����^��RXV�p���!���y_K�ڗjGY�����X��Ǖp8���ħ@\�l6fN|��Y�i�%����- ;�h��-M|ZV�#em�A6�TGGU��P�#��m�o�o5����gu�����"�h=�!$Be�d�:Y�����v��*�� V���l�BrD�զmzd�#tZ����<����7��u��}����u#�/���K8�H�O�̬���������=�_ll��Y�l宭��M�uӦks;��0�A��ԩS���x��ӧ�>��_299y-�� P�r��4u�dB�W�`	a�rGV���D�-=�P(䓘��6%�)�hT��4)�����Rff�yA2�N'��؂�
�e@�M�$3�7��(��v��Fv��>�l9ނ�*�ЃX���l�l�n�/�b�ۮHE߁t`y��4�6�M�.u��8�|�qS�Mu�H+�̃�-l�c6e�磸�ڢ�A�K$B-�H�&&Ҽ���i�|-il*������7�������l�#�JDG���{�z9�1"�	���ద+-F��855qۙ���b{�{qk[���q��GV,Z4z�UWa"A�5:��Ln��N�<�f����_��߿nppp��@d�8���X4Б����!���	hJA"�������Yhi��E��dfllL��z!����J��б�3�0 C�E��z�%jxPH�"�;�aCl��-4]�`�H���
�`%���T�X����C�º\0��߹��䢑h:�e"�0��#�H���.ה��i���#��2���p.[d�J:PŒcß�A_%\��1�miE��M3�g2�@6���� �u�6�h2���M$��|-\;���7�ŘU*ƊE3
�@fBS F�!9���LM��x"�H$Eז�a��&9H�6KQh2�I�Y����!�dZ'k�<_'�Ta�aؾ��
��x*�z�ٳg=[����~�o�ҥ����7�y���`\$`r�`�p��S��6|���088p]&�� �h9p��B���3�L`�8�YIja�����6�455	B��zP�7;;�LO�ňennNI�R�(��dj�E��+�,��1W#��
��p�Q�������f,��ж".@ZR@Z����D,����@�&�3d+Q__7W__���i(��@bb���ڂa�3��!���)���	��+d�B���|��V��!EƵT*�[�&0�B�Ā ����&#��H��@���%��@?6��Kc6W�C?�a_Ch��f�ղ�r��+]�����K�����QR���aE?�P�9�Ldg肄��/���}Wӄۡ�'�Ϣ-���4��WfR����>�6/<����g�-[;~뭷f�l�x��������1^|��رcǖ���Z���}�Tr#�n8M@2�����t���7�#�immU�$(uuu��(�EM̙3g�ٙ��Ҡ�$2Hj�!�B��h#���(�C�H
��^RIhJ%����t8��s��DWw�@<^;��l<�<��T�b��6"����fW����⽈M ��Ż���C�ƒ�dpjj* �����kNL�-휘�lK�&Zs�|<��5X��P��˴1��f��҅:��q�R??_�����O�)�_�C�+��
�wn�AS�p��0�.8==��#�@pU2�x�����Ç��>p`�3��ַ^Z�j�ئM�0�Ne�#����q� M!G��>����?����#��o)�+�M�~G!�R$�Kd���dn ��d}f�̴��	a�
51��R2����BMr�����I�\��#1&|G�I>
���3����4�6�6Nw.��X�1���<Y[۔hh0�L��x1�wQ-e����	� X檷�{>�(��33�����tn:4�7阚�i�ߖ!Z
���I-.�/�"$~�*�k��T��[ł��x��_ْ銶w}�<�fȱ}�U�(��1�
K#��u@�~�����v�z���۷�衇z���3�?�q!���x��B��k���<q���cc��d��K���s��jz��rF���(dnB�����Nq�300��fc$45Q�>������A?<$3ؾ��p(:��h�o�kni���^8���1���9�����W���<���f�r�����.fV>?p��2�Q�j=���p_��=���0ٙX&;h���|Y3�g86�9+tu��& ���O�݃�Su�� �������;vd[WWǮx�(��+V���U �S�NE��,����K��O�����m���QC�%~��2�G�������O���}������I
"�I��B ��Ba���k#��J�����z ��b�	X=�&���ӝ�m������|�PWWK�ЁĴ�)�� }jzzz4 �j4:����T�O���d0m۱b>�2��>��0ܧH"���=k��]����~,D'e�O��75Q%��_�tQ&3�Y�S���KH�*j�0�@�֑������=��c�/����O��6l�p���kr���E�#�� ��0���������|�3��<y��SS"�	A�cEmz3F��Z":�A�/�@P��Ҡ���2p?�	J&Go�x,
�ƿQ��q�ӆ�PB"II��O����x}���Ovww�.\�d��k�Lss��d�\�6�kph�@`rR������L��o��o�3�L�i��i��V]�*�[�b�e���������,ۊ ���߸.���nra_��Z^�yx����At��ב}x(2O5�5z���G�%�+)�V3`�Ս##�g2���������=���#H��e��
�;v�����M�c�7 �xS&�^Y��(:�b.Ҧ�~3�ƲJ^�Y]D�Æ  ���hjjQrق 4�䘛fjJ�Ԡ����ͣ�Q2FH	xO>�5{9m0�:j)8���MM/uvv�X�lYߊ+&0bi�ڵhR ��������{zz�Ã�c��|p<9����}����V(�ڋ����2�(����a�ڒ�D`�0"�^aR�ql���˓��AU�d����~���Y9��AA�������l��sFv��&=�G�yud�i}<£�8aAOX���]�Je�ݻt���v�ٹ���cz���i���3^0�a0^!xZ��}��wɡ���''Ʈ��o��D&$r�(����!�B�uQ3Co�HD0��A���Q�������43�t��ojg��e,�n�t(	��Cu�����]=+W.;�t��i 5�ŋ^ς�#0����ԁ8���6�e�b�����!ݘ�����2�2���
}�;�5]Y����`���ߦ��9f�D��9��mS|�!kb0d����y����*�#�dd��'�+YTm�\��q3H�IFZ�b �5���C�7�����������466?��Sc����U!s����>Z��.��0/3����l����������T��i��${@@0	�of��͊�]7����DB�����53�T�X��pm"7��@�iKQ׵��j35�5�����6[�|�u�֝]�h��9�y�z��@ڱcGȌ�H$B�јϧd2��l�����.�.uA���=�����m7�~� .����c6c��e?���3������O��*k`�F�d���]a=������ي���s=�-�z�l�rm�3O��!_ʕC�;"ŏW�L��㖏����Yeb437�!�m06�'�'��}6��b���H�x$�oZ�r��<�;�iӦ���V�����x@a���ٳ��_���cc#�67;�F�� ��E�L���	�Hm��Bk�d�j7�@��M�#��Ar��X�A���f�@45�I�su����Ύ@b�\����'��k�@h�דό��Q����`����5###ᱱ��]w��+_,t��� �%��"�Tj�T�$r-܃���|-��R��$W#S��[�䓛��!�
Ѐ���F��3�H]�V�_��6���)������K�,��s#�P���V��M=/���ȹy��ѱ��
5[�<��O50�;�_6)"/88}zp���H$���������ε��d���Z.��8/��0�`��3�<���/|a����W��Oޒ�fV��k��o��z�R��~�lo�F�d�i[�dB_���O\��QK�@�TRK~)�7��M 
 ���L4=�����ʕ+�Y��DWצ��Ж�/9|h===��ՠT]WGF�m`=jQT �f�����l�؜�$�䲅%�B�ö�v8b��
zK@��E�1Jt�J������p��I@u�'q,�
_��e-�8�B���a����L�Bsb�E�=�P����)9wQ9ܻ2N�FY�69�YLs�zaJ���MI�%jz	������1\`U d�V����Rnb|l��@���z��p�}�����ߏ5�\9�e��¦M�,&;��W 
�]�v�?��O]�w���ѱ+a�:tb !5<����O�I�5q%�ݲ^N�ACf&r��p��)V����&�O�`ssþ�΅/�X��Ě5O�]�0���^|�%�{��ux;Ggk�K�������W:��`���>�\*��Q	C7�A�E��AF�����`�d�@ah5��Z,X����l��:�RC�^��s�uT��>&mB�����AY�H^H�c�-��
X����)b�GV���}��u�Y�H�-�e����w,H��T�[Ǐ��f,""�7i�ߤe�}��&3����F��ѳ@���:��������$�ϧ�v����������M��g���P襗z������?���}n��K/�^w�u����xy����%!���z�B˽ﺾS�nN�2���
�-��A��HL��+ݠ�Eē�eqk=Ţ1�4-� 2C5�p�U�("������jjj�B!?�P_?\�X�\wG�sk.YybŊ7��nJl�$�5_4��d�eǎ*\/���������&#�N�=bۅ�#���9�˷��5ؿ�4����P�¡j4M���VQ� :�a���R@	�b���Y��h�d}b0|�2�i�!դQ��1�M[Q$ӌ��Z�y!_`+��ZWx�.��߉�`�-�N��91�q���) 
����ȭLn\Qr57%S�aA���e�����H��|����髤��,�t�	?�I	���+� ���͑�MH�, \�Ui�+�Di˒Q,�͎W����!�3�P�*�a,�	WX��ŘP�(&ә���������{�߿�����u�{���E�%��yg�oUvJ~=����K �q�{��ؿ�����r��� \�s�|�¸剜rҠ�@� [���GorrR�����|p���&��"L�	X:Y�lٮ�kV��]q�ɋI;�o�>|u�5�O��O��d�)�KקS� 7mɹ&�k�� B�FU�Z�,���� ���h�,,�&&�l����Od�Xt�`����W�eAh�����V��#e�%�} �(<g4V�h�����M���x�L6D���W�,f�N�nn"��9���|�^ ��?�[\���T2=R�) �X�	� Q�"��أ~�%-I�ϏlB�6i,OKC���HZ�okYd�� �Z�s�1�H�p�v4L�㕠h��͊ZZ��B>�΄���#=�'����~���?��S.�Y�vm��:�Ln��(���=����~�ʱ����
��
�|7L�Q� ���槑'g�P}a�:w������Go�$�h�v���a�|fB��T,;����Ժu�nXyɉ�V�tuu.���#D&466V���u]"��6�fK�`u8�� YZ���Nu���4=!ID� 0�����b����WZ"�X͇��,9�"H�cΟr"<UhCQ���|2��?W#�τ��s��$�V��$ryh�)��"���)o���}D.,�2��r"H^�RQK���`��K�W���z�i�̛�I�S�\�PNHU���i(��uD�d��kFd���N*Qa���TDrQ�eG�K%/���72̢]�V��Z�>]� �J%���O��?��g��|�G5/J~�����Ln�� 55�v�j��w��ebl�3�s�aN��\%�lV���G�<krN���0C� ��
~ē(Ri9�n�9[:�jaZ�}�`=f޾|��g7o�p��.]������ړ�����/4��l��km~��e3��]Z�k�"��v����}"���#��4%"f��JԤa��D��Y��w"ԗ����fs.󾟊 3�+�K�S���h&�'<r�~�y0�����ܖL�T�"�J�O����m����(��`>���QL���J�A�
�E�8x&#G�v��������H���(�סu�<��Fqo�9�&,oeET�LN����!�S�U6~>�S�jse�8Ƽ�h_�v8֦|���������̡��ٽ��]�;�:��.]:���P��;^7Q��Ln	Hj�������~�ꩉ��fg���l{A�XQB58���8��3�j^n����GA�� Պ����_C�'+k'C��@$�Y�pў.}���/?�iӦ�����2gΜ	=�;x��x�/���MO':�z�����`"�n�aB�Le�U��/�BN<H���ZY�_�tc�D���{2��S[v����5/�pLh0P3��%�#kB����s�f<3�C#�hWw7h��Z���!D���_�<v���$�l��yI�~w���P���H�B��\�����~��6�>��N�ܔ�Jɏ��cT��跲vG=g}u��M���=�9�&��7(�8(��|��˛a��\*�d<W���.>�w����g����/��'?yj�%���~�E�e��`r�`(�6����o��׾����o�7�ATv�y,����I�.�X-G"4_0�
ArFm9�`%m@,Ca��`��l_�~���KW�^q��ɮ����oEB�{��5�=w"��H�����t:��T��k��e�v+\O����b�`8N	�Y5�="H>+�`"����:%A*�~��.�HX��	9�ʚ ۩$�Q}�Ё�Վ�>1x�^����hƏZ��G�%�M�Y\��&���dF6�&ڶ�0��Ne�F$ζ��`��j�
f��$D$��F�`��N�{�*~�a�G�*yZGZ/V����9��v���Wk���KW�
�F�B������؆~�ȹH6����[o��}cS/;x`߳��}�s�333��ۿe�����0�}�і�~�������{��w@�V��~Mf�p(�	�3i��7IM�b� ���M����������m�F&�3�g�.]������nذa�Bfb�������@___s_߉�?��?^�J%.�_�C?,/�X2"�&�¬$¤�p�&�%B�QP	ł����}?�5��C�I�20S�	�KK �AȡѲpv�yn���6B�m�5v-�;��N.�z���^�%e61�-<���U<�Ԣ2���"�� `�$T��-Ƃ�*�#H��*k�L�{��p��'9!e6&b��"0��\/�H�����5T;6S�i��#rC&$�&�9�
�;GD+��Fu���}A���fٖ��T+˿'x��OI�4qm�N%h�_�b�`��b�c<��9���as�$��"5������?�W�Z5
;��l�����0�����}�cW���ߐJ���	q	�0���4Y�B��ތ�W�}�W�7d������OZ	0p,,Ti��ihš�֖=k׮}��+�ܻbŊ$,��Hhb��˱c/�^Q(���viM��t�ﵘ�C$�S�0_��C9P�ܜ�g��N��D��Z(�%u�����9�k��Ie&��Op=���<A�&"OH���n�g���52�wڇڃ(kl����!--¬e�D�.�+���}nd_�ܠj���ԇt\ٹ���dd�ze�s���q�����N6��~U�1xn�4>ϩ�%k��<�ߚ�kE䍶!BG�#j�J�3�w_05&��m�4���Fkjn����{����Z��}�_<r�嗧7o��_�b��`r�x������������o���	&�Ű`Z}M�O ��B�$	9zKF���Ȫs�HQx����9��iX�-Y�dۺuo�~��o:�iӦl�&Kׯ��{���egΜ��`����Z�X�9b��I��@�.r %SE��Q2�YH8�B?�v���J<��wE!�	,��=�5D�߲ sM}r�.[��]��B����
X:Vɓ�r��,��Wx�|���rz&-�]cu�^�o~��|�6��7����>Bd��L�7"�31F"��Q��Z��~V�5)X@�2Q_u�`;�3�$E2�A�E*�
/���s��3.[�[�
�F�{N�`��S�VҞ
�g�o@tt�[�{�C⣔��ggk���U(������w�����җ�tx���3R~���u��9|�p|Ϟ=�>�������č�h55��P��!kZ(�*��B���5���G!Ǵ�Ԡ�i0��Z��7��M=W^y�8���v���'44Է�ȑ�K?�ɏ�!�N�M[��	������t�$0�`TkdH�� ���kƿݨ�rBB�д���j�(X�Fi.��H�����vr�<2/��1X���]�bTHҰ�vG�,�Ʉ#�tP���Pi"4�;��������o�?��O9��r��6ˤۂi+�� d�C�5�W�/i�W���o�2ñL�p���}�d�,�\H�G�@ji���t��}�Ҽ��W�2B٧1��L����:Mՠ�"��a�h��^��f�=�J�{��ч?�O��q�ƾ�n�	�q�͹���1�188y�ǖ=��[N�<�k��]��ZlbjRs�REvZ���5u�*�`�̠�FM���ր&̺�:���k�x��,L���/_��k�ٻf͚�ezB�ӳ�>����|a�K�^�ljr�j˶���6� ���F�6+5.�r�D�ܸ�F8���[�	���"2�a?,]���|ۡ�#�O>%��7�~���Bθ�N���g}��q�\�+2��*�`��lK�(2EV��-�'��j�0	#�k���r�*͇ⷁ41�x>�q*�W�1UaS�ٮ�&QUE��e�9��xE���B�kj��oa?;��E�ʄ_W�:�T�}�k�C�i|��>��)o�)����'�f����.Y.�sl9%����R�m�	j���Ɛ�+�������Y-��l��"<��<���Zg��7�LO83xf��޵k��UW]�R��0�-Pc��O�~��_�������06���s�x��s �r	�	@�I	g�0I;^�(Λ�	�Lss��u��>u�U7�x��WL�i��$�����󞿻�cG��Z4���eж:��kW��!A����k4�_ԗ�}Ad!N�FD�P0���	��2{P���d� 	P�>Pn���	�-��Y&L�p.��MV�2C��+�]QQ��w�r���,��J�Za�����y�T�[6���"��i&��@�"u�tPyV��q���!͆N�R��1z�5�����}��L�t<'rU!�oHCc�4\h�����(�M6A�f͊(6����9�8j�Kv�h4�还P$���y�N��Z1�T/QXMO�td2��ӓ3��w������-[�l�mo{��c�Ln��������|�3o:x��o�%o��]�w�		
7�|e���{��A�=�8^���`%n������H$�RWW�s[�lٶq���L_u5^��^����]����7ݚLέ�D�-�C#Z�f�je<ӛJ�7�D����F\sR���d=g֘0;!�A���mgf�|�*�m�#��^��D�0�T��S����������<�8e�^�|B�z2I�{-Wr�6�!!2�P���	^)?�r���z�ㇴ{�J�L'��U��5�فX%��>,G�Y�H+�L����G�l�}@f��k)�C��TF���9� �wl��rV��~DD��˖]q}46(�̲˵�d��k��s*�M��`�=>.zf���N��*m��`8�����bG�)]���=7�8u�_�򗟻�.d� �Ln�(�������wߚ�/�x}2���l.��
�R	��*ke19RVZ�pI��i��A�ŁŁ���Px
V��[����k�9|�W��]�6s!�4333�G������ґ�+��f6��u�S�����I�����"14ø׏f)W3�:Gn��r)�rx�{��,X�@hk�^2��Hʂ^��p�e�S�+i̪5'�&Ā�������o��f���o�|��d�V�?F֔HcMlSD�T/[���Dv��wƅ���Ǣ�6�y�3������p4��)9��=��.�"͙�~̘-�C�>/k������5��zY�V&�����G�$�I�M�WBP�#"j8��I�$��Z$D�C��ʩ�<<�NYK%��v��֌���pr�jl�4�OOO7ټ1�ͭ���������{��Lwwws��&7��<�Yxtt���޸����g�H��+� #V���e��(q��m��'ri'��P:}
�ERK1��Fc�u]����K�o޼yx����k���~�I�����& r�|�������U#��+��L��E�����u���OD *�Y\W<g�r������证��ѱ�?��쬟�Ld�"Ti��!"�����[x������%P���P���O���B��4��t:#��=����RvJEIU�K�%���2�X�-�I�Uը>�q�n}'Oc��'72��I�!����&/
w�dO�:$������`�f���F�ı�<8�+��#k�^��!Ⱦ6��F�M�#�X�$E�'F�Oږ�̤?ְ��%% d$�3C������&:[rR�JRb@�vm�b����`!�!��:W�W������Y�N��jk�.�yi��'���O~��-��2�^����;��0^�p��s�CG�\�c���������dr	����ry��꿍�[N�F�M�T6���r��BB ��7�aat,�I�����mm�Ͻ�Mo���/Ȅ�������3;vܴ����:��!�L�����^/�V��l>�Jg3yO觡�/N�2)�I��!.LP�=����C���H������˕���K&6�������ǡ�sM��,�-�|¼6�T�U�/GȔM_�&ZHK��ρO>m8v	�Y)
��RQs��唊�(-�.�-b?�J�;���PIS� R@t�[�Ȅc�H�˙�m�8��&�.��y�R��-ԼP�:�>�V��x�T�js��\L��Ll�Y&��T�#�LĂ���v�8�OJ �4���zc򺹹9?��ȧ���'m�_r�q�D�uXW�*k��
S�L��H��D��H��/4C�4`9?�K�`��ݚ�X��'O^/"�9r�={�`)�Y��z����:��׵}�ַ�ڵ�7O�>�&�z۴utN�7d1j�<� �Ŗ��e�E�M�x�w���f]�	8�N�\�uww?�ۿ��C�4�����\/��q߁}o|z�[9rs:�\�7�1���iU�ъ�0�b`z�t�[��QK��9q���C�鴬�A3i�܁��&'�}!V�UĹI���J�6%��Μ�G*�Gv6v�g�B��!	O�>�_.A���7��O2���h��D�"��/��*�� OAq�m[-������,�3�%A�Mi�>ci&	�t=���C��c=�3W��!�,F��Zu�i��p���qM��\M���1i�j�N�d �Q5i��UL��|K��N�ܗ�1��bA yA�*�q�hՈ��̎��[j½�HJϙ6��U���^�7&GT�r�#j��%�>��n�Qk�փ�Q�G-G�a���;��:�N�:cMMMp!�Tf�L���r�d�T�����i�V.u50#��α�q/;Nc�?�̈}��]�m���!/Ɯp���/G�厽��-��>?��إ �����ٷ�K����Qoo��u���+&7��P[3����К'�m���C/�&�Nt����Ɓ2㛜�;�
F]����s.�:�#�|bE�P8�o�(�Ƣ��X���z�����;����7/ȵ�G��ÇW|�;�z׋�^7>>�&�(�M��gA
�rR8�1�fX� 'bR���obbB����$	���x�컀Z����=�����$�dg��dx��N�'�i�|�섐���9�0f7l����e�X�~:6it`��A�·��/�si�>g��?����`�o�\ccc���ٌF�r��F���\��+W�NNN�����E\Љ'0�F����X29��SB��\�6��0+4��6ht��8@��٥0L�&2t &���A%-�0�o.�@�}d6!��T��g�R�����l.�f����tdv�[%-��k���q�#����D5U]�'����E�-87��ـ��iu���'�M����vQ��>(7?S���L�)"��:dbû��1#����gCvȖ���0��G(��N�Ŝ�mI�
F�A{��%�o8{��w�m۶��n�Q/pݸ���0^3��&8::�t���on������\��X��}�/y,(�\В���$�o��l���H�(�[�,L����\�|��ի�������/_�kML���O�����ȭ0��mx�4P���lo�w|M����W�Pl�\�Q�����W@9�V�����OC&%ޓ��ɂ��^�$mW3��&'����!D�Ȝ���8?��(
�+FFF|BC�:.k��7z�	q���p�I۶�A��6g�\�����pMM�p,�[�~y�A�^���1q㴼�������l����@<����3�tP����p� [��:�X ��~�E]��e�2��B/2?"i%_�p8���B�X#���h��.E�*HtI�� ���E�ښ��H4��|�>��$�gg���Ba	P��~Mɶ;4Mo��Zm���θ�]%?8�C"�b"eD(��c������h|�x�>@-%^?i���5b?ʭC�פA��Ȅ�ֻ�����c`���YN��q��I
�`0���v�С�ccc߂g�{p\��z���qу4/�߿�gO>����X(�g�� �Mp�����͋rf HAoq��F�=B�r��`�J�dx$����i��7_�=�yOZ��E,SJ�i�S����O�H�X����y���'N�K6���5,��(.����}Np7�%�ބ+�߈��Z��%iGH�TV�V}^W;�Y)���/�:Ⱦ#D�H�"��He��{w��!���r4�O�`�p]Շ�M�a���t�8�EN���L�`�hmm�hjZ[\��ق1`SZ�x��G�������8|���߀��g["�i�Dԕp-�,�2�/�����=ŐdM�F��A��P�4�#��_rG]_R�Ju���{"B��4u�&���Z*;��KDl�~��[�\z������8x���M2N�8�Z063��셪�/�gx��V�}������,�!;��}%jq,/hm��|��@��"�Ns epN$g}��(wT��њ�n�@Y>	�����	��s��D��~^���o����c�������=v����	 _F0�a\�@'ڡ�����{�7�~z�oNOO�Eu>N8���9�e�&u�(��,C�5"5~�Йl���(��J0��a����lmm���W_}�O��O��������:Q��O�:�~�֭���{�O$���]4C�DK&"���o�8�����^SAjI�А�pZ� �v�I���A$��¹�����B>���*"Urh5E"I�o��2Aq}������4^jj�C�'\�<I�*�0��֡��t02�(lw����$���dV�X� �g�~��¹�b2xm1���k��7~<����~Y���a\�j lmp)���a��Z]�\��fY|~PЧ��三��Z`����m��VCq������~�a̬��~����3+U5�������9B��,�������'''k�5$��u�b��X��, M�M#,1��y�@#"M�/�:�~�;E�ɡ��+�~�ւ{=���zr�mQ#'=$�ee8�^�� �q?q�0���5gJ4��u�}'�&'�ϭ��O���C7_}�8;�<`rø(!4�T����/۾m��/��^��N�/:̊� ���E�d�3�酟I"�clׇϋ�pB�H���@|�.��UW]��G?��	0��z��UA����\�uۓw��L7�1�O�I�
N�T������"���F�677)��E����9\��\�Κx<�!�ąDd�6� ���}�mii���ތ��R�o9D[&6�.*�H~2�v\P�@�Y2
���� 	Ǟ�>Mӏ��Ԟ���=�u��K.�����}�k���Gxp�{�$�>��=22���>;�\Z,6¶k�?��o��D�� ��Q헂j<MN��Ǳ��	�2
�S��>�(���̜ 2eE�B^�($RA�{qϾ�������~���᭷��}h� :f{Z*\��2���~�T&������Q8vw�`.�VX���)9a|,�t�A�4��h�RI#�:�of�*�8�(rI�AI�K&N\򅐸fܖ40��x&H�Hٛe"�>�L<�ܜ�� ����f�=ONN��N��f#,�?���:f�f����wv6����jk���;��<y�c�>���� ��X6 '��@X�w2"��9J%��]��T�|&c5�}��>�v��W^y�it�����y��C���xb��;r�˶��`
%�s��\+F����$8a��o@�O��@RC4�aDN��/�m=����XGG�0Ea���"'JZ8�ӛ/i���(@�ٗ"W(���iHۃ}��	2��s��1�7l7��������普�,c��h%�ga��"�������E��nذ	�5��6K�,|����p�v��N���Ʌ�L~C ��7-�R�.u;�Fn	M��ؔk��=�D�F����d2�;�"���b��CrRA|���6��T����w��ܷϲ�o���m=���V_�}��MZ�$\�|<}�t 怶d2�iY��B�
�hn2���` 5t=Df8�Y)�5�;��P8 ��5Q�����3B����cҍ+ki�{�6�<�O��r����Vb�`��x��>o�w���~G�,�;��D����W���^�º�Ln<�L����7>�s�=���`m��G�.hb!GA����%�Y�yM\�W�X�)#WNE���@T:����M-߾��������g>�y�Xm����|���Ͼk`p`3L�5 PTl���*�t�QyR���0.4A�B�)�	�F�38awww*�/�+Zˤ�LH�e��t�����K�	��߬�C�Dl��"VHK���dz�4< �l�4�a��qh�0�?d� �CHd��V&���5��@�b�Gt��2�o��п��'�6��ˠ�6h�ѴE�BZ���g�>�8��h׏�Q�׀���s�����Y԰���|��;�ڝ@T~ﳟ��/�x���?�l�r��%����>���{�������a�4�ؽ�U�䬆ߺ���0�j0_�xT$e�V$b�6ҲT�T��׀�>g��$��lrn�M����ʐИG���\��!���'>�ccc��ƾ}������C/�_�M'�c���?ٸq���T���0.
��@�����߱c��w;~�����(4��{d�>��o_��'�L\FB�H Lx&�1x�{����u�W��t����}����S�y�'�ڿo�;����j���ׁ93�e��	�!^/�AD�����V<.�>08ac�5�4a�t`E�߅�@[[��r�Jo�� �r�Ey!�
��)��}(q�����"P(c.��������4�[�u�qP��`��@lN�B��X��Pcc�DWW�(�?s�wx�??�~���9��~����Y�J9m�z#P�7��Zc#���dَ�"-��\R��D���r�G�PW爿q<"�6}a�w}}}�����I�ɓ'����w= m��>�K^��)\��wMN�����lf#�f-��50~:��Qx�BDذmx8')��J/�$Ҏ� nKZR2��vd&��U�<��Y�9���>4�񜭭�J{{��	��̴?����@4G_~�̙�o?�`+<#��oh&��Ln�:����������zf׮���V~�S�MCQ9�m=�h��7��NJ�d�-p�J9(�`�9�j��V�X����7�j�`����~z���<��]gΞ�5MU�u9�������&89"!M�-�k��"�=OMM�A����j�@�,�������10O��ʹfH3�����q2�{B�0�ᖈ���f�n<.E�Ph:j �M^�%S�W��������L��@ ����m7��̲e��:;;���~�_Y����R�^���9@��с�����\�I/�B�50�.�~oT�RXUb���*�\��N!����^�U� 8D�lL��y�a���g~�{�n�����Goo�ck׮���8�B��V�=w�}������<z��'�V$�����%]������XՑP�?�[�8��]�ь .��8E҆��2ˢ�2�]���J���<>�i�%#�'�O>ADpP���$]���\�A;CE˺�,�~|�%�~8�Lp�{`r�x� ,FW�����o<���;a�[�M�4�B��nS�������&_N��b��I')%Mq`"A��S��>�����_���{ѯFQ>}��U�����G���G}�=�&���o�Dl��H�o��/���L�%�E61�:t�K�bu,l,�/����j粹D�2{���S���Ovtt����0����677#&SQ~�+*H���	$~�j|K�1��&�+x���%����|s��w���1��$�;�2P1�k	��Jc@���o���w,^���K/�tͅ
�e�g�A5�ޑ����{fg��Ύnr�F#���j_�p?tx����;��	��.h�%�/,���%
yJ�G>)^I��:���ݻw-=q������#t6~ɋ���!E���6�8q��n߽{w}��%���a��]Z���i��3��%�w=i��Y8OQk���a�gϞ��U�	j||Td!v�L�8h������Nh^D�[�]��𒊢6�LVH����٘�E_rj�4Q�"�Ҵ��e��<��"KU�׸�i�����`r�xU����6���;o۹��w���B�l4����+ȱ�B�q�D!?=Y�	��R��`��bw�dm����������{f^�0K$q}}��>����x~��w�.h@��]Q�rF,�t�@8�۰H@�Hz>5�dw�&X,�-xO�9��嶯^���+���Ѝ7�=|��[<���ct���S��Co��w
�Ɖ����)���W�����`�ľT��N�[�����a��p_�ֳjժ����:�y�f.0xp�}�a?���
�������L&uܫ��>��{]�&c*<���1����l���=.��k�D��&��ycDmii1`]w__�|��X�gϞ�Ë��k׮���fFo?�\�o߾�m۶�ٹsg��������ˀ8l��dECUsa�ha�%�d*Âd�J=�8F-jn(	:��k�m�����{���+�tR��!冓�Ĉ�wgg���`ppP�K&|�<;��8��'<>55��^���:��6�2`rø�����Ǐoٺu�=�����Ǽ�&M4��S�u�8��#-
X�p�<.i�ԨJ�Z�������`(�������{���:P0���j9r��o?�~��MЦV�d��L�+O�*��9J8��dB?����H{!�%u���@0r�Ȕl�D6�����]w��{�q�s��,��|��#Gn���B���'T�*"GЁ�5)ilh�|,,AHp�wO�<ݯ�MQ"r}'?,=��mvn����|�	�&a�c��3�h�Z�[����k����9>^x�	����<�H=
������[�/�����!�~�S#8^�P2*�@��(�q;|~�7u��E����7?��S�gϞm|��޷�=�?���1js��?���[w?y���+GG'�m���Լ�̦T*�1�R�E)�� �Q�y�po9�PDc��.T���7+۷�p�BzP����&f��5Y�N�D�0��59c��h��K���j����ͻw=��/ y{���/��j0`�ܽ{���v��SxH�[%3�E$��@�981��ON��T����y.Dx�p`�����[��|{Ӧ�{?��e���Sܲ����n{l�O�ɇ����=R4~.��x��LdĶ�;D$�uZ4�$G��������|>�:�Fv��6疷��%x����g�}杏<��]0�n��0V<N��h�w��7��H�|s~�zz�t�5��Ihb�qAj���L� �c%��X�Ϭa����@@}r��U�.���q4;=��C�?��?(�W@n���!����;���$�H�d���B��f��M���^=)��☡0gGh�A������1�������`�Ԃ ��������G��v�m�<y���+V���x$	�3�˃>���Ƕ���\c��H$�yzzr	l�"5���O�`�V�D�<.���]^?�Y��曕G}T<7nj
��CGmW3k��t�/���X:���퇆���1iH������p�[�ٱ�����+̝ۙ���`rø @����g�}��w���[K���s�������>�����N�(8]����J�.)�j �ɀ =
��_�x�#�ׯ>��U{�aҪ߹s�͏��?J&W �	������QU��h�l��q�E�/�m�h)���`��(�2�8�xc����^}��믟���ە��sO����zv׮�f��V�a�2-��c��=�̇�(���Y1�S~ ��\.<���ȑ:?�dxxX�ǭ��@[�p� 5G�[��P�����^w�u���rK�#�.n|����9��FN�1�J�P�����K��\�p�w%ό�����MA3U��q�`A��|�ϱ;FlQ���~�Ǥ����������׭[7�r^�w�!�4��/>�[�Ϳ��50�k`�j8��a�|.����sB��\Qz|N0���E�����g;���ry�]��O &�NZ/��y�O�F�h]��@�	��{g�:N��s����P�6����������\��h"�)�O��(8qR!�7Aݜ�(�ə&�����1Y�������K/}�3��{������;�u�Ooz������1���Z&�%�+��PP45�'�����oK$%����Ng禦'�k�ozh��O�ٟ�Y?&��җ�d8p`Ï��?8�{�6�p�=M�hB��4݄���"
$5^}�FU��D�:��p���z�F�ێ+�S����	G"bVu�۞�hݶ����k֬9�e˖�������k�r
>���GOmO��n�M��@g���Z 2m�qL��EV�8��1�G���ċ>��`��M ����OvQ�����n���ї�Y���+s}{�?��?����Bu-�Ԇ/\T����[o-�W��PpzV��u�;�-�^�l}�g��/m�`E�z|��޼�b�&��*��,�,�C��ل�<���
T2�D�r�������~������z��+O������޶m��w�:u���G��rCJ5ŝ�,�C��oBɀx�s^��p�C�A,R{hN4�D"��b�xɲ�߂7����w�j�oa���s��'��\�p�=YFSt�*�i�- 2�����Sq'KG-	��@��~p`�M��T*�ӕ������F���1�|ǎ�>��C:4t��0�FM�Rɇ����A�����N��j.��׸������n����Fu�7VLL
,���p�Ӗe>W[[�tGG����nt���`^����~���o��9����`��1t;Z �C��8��u��+)���*3�s��dI$�D�/S$,����������%�Q���w�%{H¾� �,*("h��n]�U����竾O[��Ӿ�V}Z7�pG��$l�@ �,���e2���|���&F[5H�{��3��n�s~߳}ϴ������}kj�>T�tk��ܴ����޽�����{�|FbT�4�s1Rm87� ��!%sh�07����}Ŝ˥�7J���pQ����<nI��^.I*�,#����z�x��F'�:"C�{"�`���>�𭷞�e�M�i)�΢�MN� j@^Z�����9�y�P��mf@�����ydco��`!e>���:a$��b��Cf���h4o���Z6{�읏>�h�[o�uFϹ�Q�|�'���I{��aTCC�	�N�P��؋�[#����J\pg�E�Ճsеh!�p#]ӕ��rS��o�]�o�>�O��,]��[��'y˗�v���,�r��wwp�D����9<���:(\��7���#D�牓��	).t��'�J�O�8��N6l��c�� s���;�&疼��Ε+WJOO/��/� `~�.��d2����h���5��8!N�]�E�������В�G��w���bSee�"�t{�9�I����u��5���?H:3H/�P��a�X7�^]]� 6��%��NB�'����G{�L8M%�����PDk����p퐶B͒��\�N2��B��n4�f9|�������X��t�h�������1�7'ߙy��ݤ���I�W!��#d{�@F��hXM�e��|d@+ɸl���~��(�3g����TԲ�K��8p�7~�o���l��!�&����
�0L<�݊�y�Cd��d,���Ř1c�<���'xV�b������ɹ���xz������\�J`�E��"c5�2xd ����u`3F�GE�)���\�i{)t�_�)���~�0u�T�VOsn���\�hѢ�G��).>6����I��t�b�f#�Wt�h3/D����1�q�!����U��_��w_�?p�������_(((8��Ɲ�2��z�����ޫ)..�t����3�1�����Y�y��
	�p�رc�7���3��ù3�AdVf7��h���:�����L���5�V�������/~]8џ"�Ѥ[�2�3g���������$�)�<��M�}ra�QN;E)�,�Pj�>�������3l�~�:�x�ȑ�?饗ʖ,�qG't%Gi�b6;Sw>n6F�1�`�0��T���#<3|穄�.�����^�,X�`;��fx����jժ��=zy�	��q�
wz�0	 $��``a���������6��FEf� ������1^���@���z�acRR��C�)&��
@��Ӝ_��x�ת�:��X�s��r���K���n�a�G�'G/h���_/9�-BؑQ���ȈD9>l��_��~nnn����ۺ�<0�L j�|P���I*�E�;�z��P8~�RU<��I0��� gaҤI�9�B:)�=�2f����[�.ꕘ�'M
�����z��=�|V����X�5:Y4p�I�	
�w��q�ƍ�-+?9�:J
�t��-��/bj/:%z��9�W�Px 08 (F	���r�����~�Us�~��8ܜ�S��G���.�ؗ~��l�	���S�x�t�96r=:KRMU���q��MMud趑a{������裏��UDl� �~�w...�M/Dq63�22m�~\#í�����U�N��7'22:<�R0+s��ԓ<G*����-��	;i��:th;��3�!�I�ܣ+W�<J ����������t]F 9���ݠf4�Â��;�D�t�5<n���ʠK8FQ�#ה��Y�x�	sZZZ*��O�y 2D � ��K���o!}��t.�g��  4�� ϋ��9�#���7��\ ]t�E�iCG!"���.Q�>��@w9���b��E��S�_�j���E��A��������uWй ���\R���k�^���/������t��$U�aÑ<��4�H{T����g�� (�"f�\�U^y�]�� 5������3�>Y�Ɍ�{����42P.��9K<�����|[�;&��1��}m��$_z饟�v�m%J���gس'e���[������kL}m���M��+�p�p����k�a���	�P�Px�Ũ��*Dǈ)�M ݣ�n���L�8���c��!j��^�$���������I�o��g�[&0�rWrRw���kԙ ���&ɣ{Žq����=��׿����_l�馛��<�{	��Cv8p���ҝ�UEz�gfaA�L
�3����2C� ;B:#͚5KZ�~��tR'��O�Ց�Ck�!��6��������l���z}��}ߖ���	0.���H�h�F�$H��9�I�[�������F��f�GΝ����F@o�4PN��ؘ��P9D�Ŕ�}��m���I��!����{MOYP�zژ���͛7��t���*w%��9q�7�[έ[���������w[YYy.m��;��W^yűj�*��̻w���k%�=���,��gc�]N���́}4L�PC��IH����fcӊ�����ѿU1=o"P�qҤIG���?5-[�L"Z�D�� ��׼�{�2+++����^���jO��7ʐH����!��O(�6@OP��� t8���+/�/^�x�/~��q 8Gi�/�۷�V[[v��=s�@��D$
�
��P�����#p4�&]r�%�p(�z��"�{�E�G���
u��ɺ
�=A�9p  �3��I��=� ׏��>���5A�tڴi��\6�h�wȺ�n=t��=͎������U*�Ɉ���1�KD��ୁ���q�F�q�Jk-���Y�H�?�����Ν;ǬZ����?}0��<̑O �����A�Έ����g:�wx��/}����@����<m�򥏻=��hv���	��lq�q0�̝���X�gcm�0�8|�n����6Q���������o��^cD���%-ҴiӦ/�ޭ+**��l6�9��_�\��ȄA f�ffc�� �ʌ�� Vf��$�?�hћ��_~y�c�=vZ"8��SRRJH��LOO�q�D
HU��W�Vؗ�Og]Gz
� �����R3{8t��i� q-����N�tcx
9"���Q5Օ�Hޞ|T�O:oi4p���Dl�{�zͺ�e8p-�}��Wͅ��	R8�7&6^���v*E����^o���˩&�^C���9s�EK��C)����o���7�{���A���.��&�#�C����#�cH�,H�����6�Z���Of����?�ڵ�M���W�hni���a�i��S�!\��'�bJ��Y���o�y��4ܭ�]+Hп�_�����6[Ē!C���E�=	Xjr�f��K��'�=~���Cn���t�]H�ot(�����4�eܛL=��IɎ��o8��`��իW�/^���{�<u&H�gdd�c|)--��;�xIm�2{�.<_�f�<<|}cB���Li����ԩS�)((�����J�'�9�>�A���\b�m�<��H���� SJ�J�o�>�f��-����;<�����+V�x����g��q ;^a���#F�V�����E�.��~+�,�V(�R�ቈ���x5y8]r�%�ꚓ� ���ѫV����|=(�1]�2�H��
�1���"^x^����F�m�^������u�-]�����Y��������'3+F���}!� �}����d�>G'�������$�䎎��1��cc��ϛ7�xg���&�G�Tr�ʕ+�o��%��U������8��C�y0��)�h"�0H� 	
���ut?u�<�~뭷,��>�O��#�C �8���w}_G��.P��S��x��27�ǎH5 � �	�/L��Թ@Nm�c���F�S��pm��0��ZWW77==����B��t�n4�Β��5�<�_�B{skK<�����F�����B�9\�E�̤�M��[&�S��������=eʬ����=��u6o����ܜ��uF}�vO�!���
fVw`��>l2���C]��H �������%y������0�@�}!ua򶭿kin��p<���]�r�����D�v*�T7J�0>
�U��K�~���-.*�]����wY,�h�袋z�����e8�v��Y[RRZA���� Z��X������9�8t
i*�b���)B�,�z�������|��g?AM��8v�%]z7'''���U�����Gz�"������v�����&��"B
Gd���Ҙ1c��k~�FGtM*΋L\�G�8�-R���n�<��O6%�H�v�=9T:�9����iiiU�^���Z��L4p�ɿ-���ݻ�/��?~�.R�p䂽���=RPD	��\8��������� )3y�_��D�1eʔ#�>���xD�I G�=u��m��Gا;�.�H���6P��0��f^
6XHE9����6]<��Y�n]i�"i��6o�|��W�����t=M�T�gCn���%<=�t��n�)��J�����uDD�����O����O�t:��qq�����+�@�&�S�Q��<�̫������t��]J6"���q��yee�Xԑ�B۴��a���l5�����1�%�����~��SO��� '77w�믿BA����h���[.6��B'1v�9�d�.�8/H��ѣ�$qڦ����\�&�w�b�J��+�Q��-D�aW������@O�PWW�����K�����:� �n4���f߾}�h������VR�8r���B@xF=f�xã���K�mR}#fD���Dl��勎�,�Xl����{�M7ݔ��=M����mܼ�gn��R��h�`�APF.�V���>����DE�GSSS][[����|}͚5':a����'OY�l��t-��6��P*��?�S"60|xpk)�OU��ǿ�(86ۤ�I}�w�;��ғuV�egTd�'�F����O;u7�&?��i|����geeU���0�{W�#�M\��a���a!�=��N�m�b$����`��o���FZ�?@4�t��(�MKK�x����*��m���`�đk�(�_&�3�(Nd�Y��=�mx瀨�R� ,���P��Qf���a�?\�l������U�۷���+A��u���Տ��]䔖*C6{�}=��M�-IMM�jժ��븇��wMM�ކ/�g�-!0LPZ���2'����U����썉�9j���;|��5���OU�z(o
���~��9L��X-����sF
�;�8�#��`xV��_"���X߰���S�}��G�2�){RF|���� `s�i�6�#F? ���:�(��� ���O�~�XN�<���f�-�ק�'s���G�@#����t@.Z�h��\t_z	\�cP��{�UN��^G���ڐ2�I�̈́i��<�t�͛7���><-m� ��/�.]�������(F���&tQ��z"�#�ؙ��ћ��.�ƍ'edd��8�a� 9��ʀH'��T��ItP�z�Qr���}ˤ�nL[����������t��n4�VA$!%%eyD�����Io���q���H3��4�&%&��b�ee�2.$Z�#""�v{D�Ao��x��)�������Yꉂ:���_4�����DEEklv�Y���GtEq:J<zQL�a�`�LFScEE�q/xzÆe]Dl�������r߀����S�+ߓkl����2��\@�8���&�I�Y���"�{̠�<b��%/��t����L
:�X�'{�?Ũá�}` �3p�Gr�_��#p����v�o�^���>��s�o���G9-E� |饗��۳?TUS�_tl������b���A$�i�g 6 �E|��I����Cq>�5�⼡�4f���r��R���`��>c��/h1M�7oO�^[TT����Û��@4p��7
\2c��
��w���xRZ����,)��e��D��f5O���FD��n�@�""�k�S���^w�չh�z�����Kٱ�&��4��]��y���#�8�"�Z����0:m��iN�pѦM�ʺd����{�759�q��q��1�h�p~���6h<�^"<HDl�E���xv�m��/�`\�O>Y��>#i�ə7��+W<x�]Z��j��1b4�8H�`a���(�x}��\l� �#`�U}H||�}K�.<��s=���e1��_[������t��<9:���6f�L)�u]�q)���`zРA~�SWccS�P�6��� I�~[[K8������.�V��"���$�;�vpFu}LAaт�;w��o�}�h����M�Ю۲n�͛nw����{���B���C�S�h����f����B�k���:��X�,6Db���Q'H���?pŬY#`ӣ�WKJJ����A`���=��]g1Y	��$tI��^�^��t��>�U3�8Qtp�Ё������6eee�.|�Ϊ�����xxiF�^�!�*-�v�Ԭt~��2���y���a��.�F�I�~%GSS������uWlt��]vI�/���P��/
�qٟ����;���M������x|9�"�Dd�����D��J:]� 
��[���o��b�59g�\�ᡇ�v��4:s�#�<��%�u��j��H�	@�l	���!"2�� =�U8$�NvN���#F;~��!{��m�R1t���-��~d�*�h�t��(�76���
�%E��O�)3��N��~7";7��/S�D��Q�9>>E7�|M��Z�v��5�V���q�DJ�!B�A8���Lt���m����a!�
傗b2YB�U�,f�q�G���?�����A�꣏>SXXt�d�ȧ��&���t�|�c��U�WW�$&�y���������)�>���kJJ
�}@d�`B@�X@p(�x�k�r�x�BCxo<
^y�YdL?����Ob>�sڠir��bʞ��Eii�'{?QWW7��79�:,����C�yK�̥Czz�?&ze�X~�|�r0�9L� +W��&�����Q��Ek���A����n�3��; e�������'7nLJQQ���֖+�V�4��߃@�9J�r��TVg l�x��e����\_�p��#�����4�$����&�O��t�5��x�?%O!Z~_	s�Q����rG [p4`�G�pCC������}�pYz����ç|��O4?��RO������۷_���`0�-j�P6X�I�m�0&0��.d��>\I�n�����UW,�����O&��K�?������Ձ��y>w` 0��qN��+�u���3ν��Ȫ$C��o��K�O�^L�J6��xA��K/��qǎ]Q��1�q:�&���f,�p�����J1b� �Xđ��d��=����# Ҍ��J+z�
�N�6m:��~J�:�l�`:N=�� �_#���>B������L�e襗�X6mڴ�nM�,((����T������]\�V�	{��)Do��.,|<H�ͻ)==� ��幜����&aA�bɧKF�n����Ʀd@0GE����u�QoO�56���9�R�FFF$���i��~����l ����Et>���Xn�T���Y:<g��w��!��A��n�aI�YQ�>t�vm�n͚G�:i��6�&���v���yz�-��ǝX�
�0�0�d�t,�X1y�ď�z�J�V8��Y$�?���t��{}>�c���B���="R�@�<<ӎ�hZ�{S�����H g��`ޞ?~kNNΖݻ�ƶ��>@o�"P�c�M�0��pD�q�v����kjj.8v���I�.����_�z��̝;w�)͢�Ɠ2pd�Et��a�
��l�>c0D�1��#���٩ʒ����C����6�)��DRQ�~�d��/�z����V2$Q�8딉��'�%<�^�<�9l������8d�[��;w���4�_Ijjj�������r�zt?q1#��V)���;��k�%��w�ԩ��z�o����������t�_�Wz���eZ���X�e��'%��ʧ��X2Z4Q�D���� ���/��!�u�s��D�D�o8K�.]�q��Hҋ��H0���)\ၒ��a����Zѭ���!Za���"��}��ǯ����3gN��#�y���������	L��@N�2.�	<� G��xF=]YYY,���źsܸ!�-Z����Z��ӟ���-�SEzo���`'İa���l) %�>��W
�ʹ�+�g�b�w򻕕���A:�&�k�FEX�dɨ�۶<�hi�)��>(	3�rĆ������;>��g')�26�M�2%�l6h���_�
Cx�w�#�g�Q&�bb���'\:� �����K���̮H	Q�L�{NUU2K�K�|8�&_w�/����P��y�!2l���,Z^�=��-��w_3-�&���B:��t:�<�9������ɶx�� 8� tP���ۦ�Z+��euuuͯ��z�2P��Ӵ7�0�������Ҳ�t|*����`���K tFṢ��oll�u�w�>JǘO?9>r�7�/��Xvv���|�����j��5>�.�&L��58���5�m��~b2�"�


v�9�JQi��<���;�u���555�HJ� �H�[a��O�M(�<�V�<.9��VD6�2A��d����~��e�C=tVy6lH��Ͽ	Ž~�F6DzQw�-�\��M��
��F�N,X����>�ӊK�gd�����Vg���t��n �l�h���9���|6---^��ބ���f͚�� e+=$M49�:ER�z��w>��� 9��hlt�"#�t�\���������j��߱�����b����?O�-��t-�/^��ܼe�P������)\DlBz�Q��%��6SQQ�����\r�����Z�Y%���~��rӦ�w�h��0�V�t��'��]b`o{�S�������G��w���%��,V]s�#�����������RG7� �|���#�����֖[規�"���7 ��q8�.�V&�#� D�����ܹs��t�΂�ʢE�.#�q	#;s���m�~�;2��J�������7bĈ�O?�tCW����X��.��T�g� I�|���`L:ޯh��yZ0>�T`���SOCC�~E�^q��۵VoM�%Q N����m����rذaqz�0@�-$��%��a�ŷ2OL���!݊����R���Ͽ��v7�!@�D`�3�����.,�]����9^s�Ϡ����w�ر��"�RRR��ET�~�:v�ȼ�>�"3?�诓��FTWWZ1w�Ng�N M�k��}`��)��]�!C�ܴi����dw�+58�9����!�S��kw:o�x�����e%�S��x�EĀA�У3JQ�QRdDd��lNILLx��;��O�Yl G��_XXx5�~����ɢ|�}Gk*�&w3�w+�Ȭ��o�ו�xz���	�� �,�
N�l�"�%w_E8Y�r�ڝ�pQQ��V��P��t�E�&MЀ�&�(�2e��a��$z^@ ?��L�$ױ��S��Y�9�`����"1..涵k�@�u	����ǚ��[Z^^����'�9����=���ı�p�^�q�JQ�����rX~z���C��je����ڷo�ҷ�Z��������UUU�8g�R��b�3���̬n	���5x����I�+�oߎ���2΅�n�CA�iÆ�6lX��vg�]�}1���+*(����P�%5�tll�n�;,6�椤���ϟ�l6(�{�?�"�6��
C�6��-��(x�4B��������o�}�5�\��b��W^y�'O��f�"��G����6y
�&���\���8���C#��#ÞI����ٳAT�M�Y��NzP������ԭm��N�?B��&A_��XD-`����͒���v��''⁵k�֮\�rMwwPa����˷/[�b*���	�D3+1�������������ݮh����=)))k�̙��۾�KZ<-���OJw���9<���Fd����6���*�\*��l�;���#���]�vY�wo�-K%�M:�E7� �$'''nݺ���ʊ��!oZ<�����F�҅��4jk�ĭ�PDzEEG��c�һw����sO��i�|�Y(�!���˻�N�������VJR���[��p�~2C�]��/Խ����k�����֭�w�Q�p8JgS�Р@[�#rc��p�{�\.�X9L҇龴��yg���O�&��4Q"8��z��m�R�I�n��#8��E�
�fx��h!�i�pf������{?���]����;*����gg�^H�y	"�<2�TjJs�3c�!�b0ѝ<Y�7::�#G����S@i+))��ݶm��l�U�vF-�����Bz���85�d0�&�����VK�~��ÙV�o��o8�ST�9�����1�7o��ĉ�X,�>mm-z9b�S�-/2a\0�z�^��@��ѭ�yl:t؛W_=7�l6������I��5��0����5��C�T�c��PL�~y������Q�IZ?�x�\��8��K�u�`�+Q1c����tp���Q~�� ����+&���O�S�O>)i��� J'���Ez�~\cs1�h"�=��."�nx`%�q"B���t195w�Z����Yԝ�7(�ݹs�����m����q|�#�}�PnNP:��c��������Ǐ��w��"	y7� xTVV��o�k֬�����Ц�وmpg%l93�C8O�F\3t�6��������<��lk!���l8�9�7����o����/R�1(h�vP~p��O��	�<b�\\+�����6�M#F�6���������?������5�K�@/�p��9\T��\���!�Ȑ5jԦ��s��6���D2PwGG���_�.�A_D��)G�07��@f��&�r85�--�:}U��4��|D.SRR��.�_NNN�tdnDD��G��S�)\��V��r�W�"�sӾ}��}�YR�u�q^~��u.�d����f�Sc���^����˺���� ��loק��紐w�>�����v��f�ƍ�C � �������evԸDy@+A�)>��������7��9�"��9O$--ͶnݺY����n�Q�h�y%���͞�!j��Q����נ�64`��^{Vt��A
<%
ڸ+�I�`s�SLg����Nץ�~���?�yNW�d���l�tmLL�4F�����5G�7�'"6^���0�����B�f}CÆ>I	K�L�R&i��y*�;YYY�P�)..N�E|�	�%����z���xQ��z�]���͛7�lڴi}wwy^��'��r4:��~����3��Y2�!��ب�7JM����v*�笕+W�uE/1p�@���
�������Z��;�pd`����5��9���ѣa��>3�홒�y�w�g@��~��H4ps�./��´������@��k��ߡE�yV���� L�X`{��o<x�����/sǏ�y<��̃�ɦ��z.���3ө��X6����h:6u�����sO�����a۸����ON�k���{4�6`l<��>�D�N�H��\����j��nOccCfLT�b��a����&�L�4���);����N�8��V����1C=� 6 j�c2��#��(��{^}��└�#��!���'����YSS��h���n��#:���0�a;̅���f$���������6W��>Pd�x��G��K�|&���-N�q������v�����
�e����l���g�#�qq�%��=CugO�J7�@�Iag�M�)���Z�c�T�e��ψ^f$��0)}�K��K���;�#���YYc�|�kkk��s�Ŭ���燴Vs�R|��B���g�>�U�~�Ν}���C�t,S�-1��=!u��_\��F��I�A������s����hr6�M7�q,[�l��؆���Io���ŉq�>îa��ar?�Y�{$�s�566�bݺu�����y��G�rb��#�����INg�P�@ E��:2Y8҂c���ȅ��ʮLKK[	����A��)S��JOO;]Wx��3p�SR��+Yl��:p�Z0@:t�������Ԕm4�t�TVV��-D�9������z8���Ζ��0[�b)
Wi-���2Yō�!]|�硐��������7�|󑳵xX-��y�WF���q��Fׁ����]8O�r�L��v�����1bϣ�>��b��|��2�q16s�0�"8C����Au>`�\1��IQ�vp�T�#���Ƥ=��l4�D-w�ygCmm�jZ���^�K�ͣ�455�g<0�]�p.�F�Yqhb	L\�����r�ʪ�l�6M�ۺu�c�������1�6�����"��e���h�kp�-�z�񺱱�W]]�,r�R�'��ǐ!C<��r�Nr�����01��,��-�Qo��=]����������a�!���lCKkی�_%��Kٰ�y�z�h��,ܫW�N��ʼ���a�Q/E�d�0#��tx ��[�3Q�J�-&���7ܰ�<��Mjjj�Ņ������5�n&�=]jH��>o�u��(���/�������)..�G�d0��i@��Ɖk{Х��������p��S�ֈ����pLM�QX������}P\\<���̎��4�� Z���7�) � Z�T1�>���?>@�����SW^ye]jj�g洷���PDnB!}��t�\��E��Ld��VT�����R�U�נ���h͚5[233/�s�m0�tu��%��CR�S�gpq���-�'G�u��F���ڳ�m�՜���-�9GeÆ�Rw��_]Y�@��K2��:L�Fk7/�b!Wڏ97��2p�}\\\�^�GEE�=o޼�H�Ι�5�XV�ɲ���<#�혊�rNZ�,,�U��7�q1�2���%a߯��E:��
2 6NgA8�1����.,N�� +�}dp�����W^9�P���D��E��&0�2��8��<��̈́h����4@��@�9mC�[I�..))��?��?_��� JiiiG�����qj���ҩIR�]S�GT]���u�KJJg�����]�E����W���lI��h�0��\&�1��#;X����jmn���m؎TXX(�黸n��!�)/��i��]t��t����sP���ڵזWT�M�G�N���X��x����G��n_q뭷~:w��&���^~��.�k��n31�2��031禙��p�]�+����
l�Z�*�ر�kl6K�@@&�b~	��䨍����ڀ$��f-}��/�����h�ɷ"�v�J_�bŲ���D�c�A�����s
0�YRs�D����j�N�W�W[���f̘�X�~}
��+h���8�Q�@���,���������C�o 7�ٳgW���JKK��y'�q���0X���r�J��"k�����sd�k0c��b���nZ���666�=��[�S4ps�	�}�ᇗ�?F�MiT/�L'��A)�U�z��+��!R�z����+?$`S���a��"555֢��)�!�������?�B�p����)�F�Q�{֬Yd�:l�6�=��ј�r��lH؀����a#�)*tF%$$�WI�l���w��]�c�=&i��&�.�]v���ɓ_lܸq ٯ���"����dn,�X�9�p9r��5��`�׷�]��8�����l۶-���h/�w��h����C�>�;3�+�B�l0���v�0�]�222��4s��y晔E�]K6Ð�؇�i������x�}�9T��)���8�J�E�r��'�99����lcOm���9$H��b;�x��_����tC�pCC�ƃ#\,�sH�ȭ��P�)�蛮��wo�����=�),,����O�i��\7�cB`NM�g��,V_��/'�nWW�������yא�	�<��k����� S&�������I�&�K�RMN�(�7���Ջ:4� �,r�,H���Z�H�"�T���$�&��8}T�]�G�b�f����9d'�q͋z��zj8w�"Ov:���~Nrr�:�[�&�g�>�|��}n�w,ِ(�>���^_����4�4h� )77W|��T)�|]#�s�IL�G�M:���E�5psɇ��7=}�/�~�,�Ym�@��
�M���I��c� )��P��ɓ'�����,_�F{���>����mζ��NĨ��Ϩ��1<n�kf�{>�?p|���M�}m��ӟ�47;."�bUS�s�����kl��@'}�uܸq��w��3�&�h���E󉆆�%EEE�i�T4����K�����>�<�U�ݑ��W�ٳg�M��t����~��ɓ�>�w���`�;Bl7�قp�����2���d��P���o��C�qL�2%o���utQlÔ�Kxہ �^D��Bc�ְ��YpޘMV)�IA�B�Q
Z$�}e0��t:���;v�2!6�AǛ��0ܜ#�Ψ-[����o"��u�yQ�5��@4��5��Q��BO3f�K���-�CL���#�@�^�G��]2��aO�'�*�8!�v�@ x�������>t(�J2�c1��W��R�9��t��	����|�*7����iQM4�΂��d�jllAz�+z�3���
�ar?ϥBD��7�^"]�s�ʕ����nq�Ⱦ6�����K��C�FǠ��³�����T][;'r�����xg̘�?%eG��P�"3��}��_%�[��a  Q���>�hB�Z�S�4����U=ٮ�f��$�9d׮q_|��������M�$��1��p0$�ył-��y=�����fV
Y}�y��ѣ߼��v8�ǅ�C�c��?J Ĕ��ʼ6P\\N�A87�t�t����z��A�]�������ݻw�H!�ǠRM���ۗST:)>>A��։@Q=�u���UM�7��kj���?%�F6���x3k�z����ő�S��M			��ݻ�ڿ�����n��B�yIQQ.ٕ^��`�
�a0��L ��-�-��͎���߿��/�+�v###�8))1���\[�VTD���ͼ[��#�(�#{ń~�����h4q�9%=���յ��toINN������@[��CD7g����80����.�Y���s�;����.Q@�v���'�҂짿O�;$})ϲ9"�E***z�ݞ�t],jo��0�p����?pr䘑��ے;|������3�=��(�z0D��Ww>t�@H$^��"	�W���������4�D��'X�sssJKK?~|*��HL�{1@",(ԭ��O��y���{�k���؆V����5��G�ԩ�5%E�:���lҷ��G�������ң�h��fs]p�Ĭ�;w:n�)vu�m�z:9�C�k����H����X�'Jf}kKˀ�����m�VA�:�M�����XP����Ϗ�9�����y-�&�M��oU�}�"�@Hr���L)�^u&&&�ehϟ?�СC�9,Ǌ�%�=�����Ev::�z��/� ���=�ZJKK���ƣ;At_q��ۄ;�������:�/���&�t�`��ꫯ����-�?����I,М.�9K<z"w1	�i"�\]]��_��W���N}wץ�^�ܺukZccõ���Z[[��4���h
K�I� ���'@Է��lҺu뾢O�����x㍌]�v�ѹ���3p�;l�`�Fn����f�s���O�2��Ki)�.�_��769������6�Rmg_O�]�9K̛�V/���� �x���v�����H�_CQ�^_�X�*�<HY�bcc�_s�5�v�p�kRZR�DJܛ�X߹�)$�:x5b��Ń4d
�ht �C�������h�L���p�K�N���R�����;�t��'%��y�7���&�������@ɚ={��![w3�E;��0q&wEvvp~|����皌��+W�L��) ��������$`3ɀne��^��<�O}��)<�vg�EG��#}��L�<��lK���F��ƶ���;wq�z�nq�.$�_�F��t����(���v�ڟ�q2��`��:��n�RټysTڮ��8��見@j���!"B��Q����f��J�V%@����{�����ѣ'�K�j��H:)V�Q܊0���SG������ut�:�����,��9S�fS?@z;t<�[��߂;�`H���9��@�ԩKε5M49�2�������eee���ӯ�=������J� g =~�v��\���;l�ԩS����Uf]C���/����hV�Ų	u�M^.��K^����/:^pS�M۟9sf���C�dee_J�aS��������V�0�VEEEx<�

Vg�����t�O߱=�@��iӦ����9u6�;�]]UU���b4�uPJ�t]�t�����*�B��3�E�K#xi����ÂJ���ēO��+fA�K�YW��g����7��ݻ�R��TRrl`mm��^�"a�������:�S����^"�K����8������o�F�QM4���	����v|��G�l6[����3�L���!����b4�UYYY����r��^�����:t���
�Go�0턪���oG]S	U�USh=80g�wW�'��{���>���UKۍ���9����Q���6�����D���.1�YOσ
�>пO����g��V7g���o�1��X�Ct����?&z�{��F%�������-��x����DF�9|��^��;O"���g{[\��dz����";C��k��rR�O�1��_�I_M���n�ε<�fN#�KF�MX���	S�%M4���ddd���ΞM�z)�xc$f/��h 0h�� ���nݺ�>����[�u�ֲ��9t�i�65�9�N�@����:1�(%	�o��̙�~��G����~�_��I�.W�(�VApm�6�����"�h�8��.����9ٷ�5*��a���!�9�$�L��<x���}z0�B�-�b��L){ ȏڬ���l�`�Ȩ������͛�%11��p8F��K
hPw	�9:�1��F�F���oC���Zyy��ȑ���#�E�k͆Hކ�k�6�9D��	UWW7�L��a�.Ң6�hr�D^�_RR������0�:�Ŵ��_8���SY���/��ͽ��?,���������Eo��0��G]G���UM&����c��s �^�]�(}K��ȑ���VK��뛁�@��S���M �_�F�d~�'�}A� 6�#xp���#��}�������

Vb�tD7g������ص�ζ��{B_�_A�V�M�M ʗ����Qm�N��!C)2�.%&��Vk��d�|��׾9~��;��tHEE��h0ĹB!�h@�G�s��ੈ
��~��>�\@��?~<������b/�=-5q"҂�u���G��-����`[[K�)S̘1��M49_d�̙��k�nY�fͅv{��6��I0��E��EJ:��Q�C=-򽣢�w�\�r7}v���`�����U�,渶�&l��;b�c��6��Kz�]���׭7���a���V�7�`�Ęcƌ>�o߾�?6��(��a�tAeLN0�".f���b��%>KJJ?�d4�E6@��iv{$�� �6;$��&h-�=!��]7����ov�ޝM�(�Ld4ps��l:4���|-���D��#ء�'�B�7Uܬ�h�ǎ+��r1?J�455E��\v��`�t�S�tSR��:9<,R~4�C�#y&1�g���Ԡ�sڋ��
M�����1bD�Nk��D��.'N,����XZZvill�h&��p��\g�7�*��G74�^�dɒR��S��2v��ʴ��c�om����ڜzt�5O6mxyy9��.�8̆^I�G3mC�4GG���0e�]��ۨ<DM��~|���b�p�]t����n�L�F��T�A��2���M�+<~ۦ�TtN���S�9���{�Oޱ�;�����esب5��F�N }%&&��	&|2u��#��B
@�瞋B�Zo4ʍ�B:}'p#�g���A�:����?:��{aZ.�ɹ�X]�ǹm5S4�6 �d��cbb�Ǎwޤ5��L�СC�k׮�W_߰�t{�G�*J�w�����C��t=��p\�y��Tz���ތ=��l@���r�	����br͋.̬�twEXR\\!}3��9��Χ�#A�.VVwMu��X�5A�"7>oG^0D��I6z�!�&���#�kj�g������?vzJ7g�l۶-)3����--�覉ө�(���\6�!���
.�/�BZ2x���7�pC��@�-bp�Zc�7�'}��^2Y�����~�����ϟNK�����󻀔���_j��D~jpP������!C�d0���5�D�O,XP��_�i~~��������zt;��p^�9"΅� ?��&���+>��ҷ��;B��ݯ_�|�'մ�X5�D� qM�Rd$�3���Mu�0�!@@��lN)mw*m��vH��uF�3��!��ac�I&(H|aGݺ��LZ�>�؊ʊ���ec�z��#�nz����W�Z>�����������!|��2�sf�D8�W�^��]O���x�[�S`#�۝��^g�ώ!_�׼Uۤ?22�V�"o�R[[3�b�Z�À;
�3�n�{0 8��<'	t����h�	�ݻw-**�I`e�7� J�[��p��/����7����򌌌��w�<� 98����דy���:|�Sڛ �<��h�~��{���u�����G����:�Z#9z�up�k!G��J�Z��K�-�k�58�z�\��˵;N��B�pqvV�씒��9C��h�nz��ڵmĉ'�p{ܣAo��S̨�=��yp3"�A��tCo�ꪫ��7�I:ODSd"I��J�����f B�z���WUU���2`� #���I�xm:w;p.����HF�E��1bD��}5�D��'�^zi]rr����ȶ�G�0;�������VYZ�Lp���1)))s���!�.�~��5���#�p��Vȩ�S��
::����K]:H�M\\\�ɓ�>L�gL���q2��kMLL��D��1����'<U|��5Z���[QQyˉ���y���i��_|�e˦��|U����:(GDT!x�>a`�ya���G gߔ)S޺�kr��� ��������:Y�ôr�W�.
�Rd��9c�A���k}�`�Eg�ɤ`�:(�q����ZZ��ccc3Ə�8i��&�_@r�iӦ�������������=�7�"��ߒ�cbb�477_�cǎ�����9����QGNOe{�ˇ9P�O��(p����<���j�*�7m�l��\pθa���4zGч�)$���[�v2�|~�=����' �!���*��/Y�)��\N�����z����i��ҏ �顂t���˧544\K7o�$�A%��&��;�/� 7|#*|6z.:t�26�g�-�'HMM
��Շ�T����6F�>�A�����N�,�C�>J��n���1��L��{-�r�j�$M4�������8�%��|��a��H���BO9��if5��W��霺k׮��~�iy����Z,�&ڟ��!��mɩF�+�7hd��ۛ����CF#]ȸq�|���մ�6r�v[$�,w�Ju��A�Gͦ�악�M�s��n_��`M��Sו���ښ�9�D����E7=P �_~��ѕ�e�3����(�d0J~�|C��+党s�HE����fl����p�Wn�ӧ�nW<�^��P�'�~��\/�.��{�7G�>5��WVV�X,f;�6 ����hJ�V���c�D���O�,1bD�L�DM����{6n�x����>��}I�m'�cԴ�h0А�qD�����ʙK�,c����			ި��F���$��̯�H2wK�}�(��H@�?�0wAd�g�i�Z-(K���U�2�#B��ڂ��/Dv�:!!1�~7�l�DF�:����}��3y%�N/�
8v���@������+��كYX��3T7=P0������ֶ�馵�[��(����H�(�MJ��Q)s���h�ԩg|BkO��@A^�#�(�"K-+�)/F����ao���P�p8b轈S���Rs4��ŕ�<d�������D��$�{�n�ׯߺ��������3����T[8Gr����i�@_+���@�!���RQQ��h0O���j0QHA�mmm	�o�>����C��T4�M¶��^�������=��<A6q���4 ���7���q��ksp�=]kkk��b����#��{駻DB7=L�����P]]}yIts���=u{��t�pwP2n�>}���袋>�0aB�N��	��v.$��k�>��	RP���!���lht4ƙ�V��n#����ſr�z�ۃ'$%��f��kwTTT��!C�pM49�2m�4ߊ+����e�N�%�`AJ�if.�U`��DM�0�]���=��S�}S.dǃ���.`v���2:�}����59����-B@�C�i���5�ыsUt��ĸ�Y�f76�]�rY�{�nr��¦!��8$jo���� }��K����v���e�#z�+���nz���O��[\r��x���Ʈ
�:�`�0bNQDDD��n_5gΜ��k��7	����N�ЬZ�p�.�؅���&���yR�-ʨ����kmxМ��))�D��h%�������"S�D��(�:A64������Ⱦ��:�a��ε)Dy��jii�d�i����|$'�o�G5����NMȩ���Tʃ���jnn6I�"�T�9+�"7�ו��S>׹�.Ck��|�ݷ�=zt�kٮ9���ݹu7��q���H�p����k?=|��f�M��4�e��M̎�9p��&G㵾�?���;/�r�/L,�����u{�ϟ�����q���(d�B��|�ý]	+�𢤐��LX_PX����QЧ�m��{�:-��� �Ж���7n�n4��ˌ3<��طo_>��>��cD���H���� �|��G��s���{��@DD��h4���Cݐ��=D��2
�lhh�ִ7ĕQ��wRR�ȶ�y<^��	dee<y�d5�A�Q��i)��`HDjP{�7�$#�G]���q��#08�XQѼݻw��.N5�nz� :��/�w��,�z}}� U��U��L��~��lF
Fo&L����ѣK$M:Hbb"�}t�Bjr���S�O����t��ƃ������;�� (��ٓa��<��)66����D�3,���ٳ�����Y����I�uͣ�pM�Rw��r#�?>2%%���r�(4��䢧ց������^Z3�܀z��۱L��M���b�B#$���O�2}{yy���T'���3�Bʺ�v�d���"�fyp���.��h�<�X�V�^�����M�իW�)(,����^���d�jܸ��d~O�pX(z�SD��>}�|2o޼�Z:��BJ"��NM}CHV|��V�3aKs[[�NU��hz��:��أS�����;�ѿ]S\\�kZM�&�� �9sf�W_}�\^^~��n��֮Ss�ԩԳ���:�M ������=���r��Ln2)��
�>;(.h��TB�}��A/}��6"����;�Bd�p�!����%F����yyy������\.s�1/�Lb}Rϲ��&Ӵ���+7oޜ/}�H׷�nz����X�z�-��W�A�n
����;�5�`2�d�G��ftC�85}֬Y����v!HKYL�����	�A�����Hz�g����7[MF#8s��*n����R�<;nz��Ii��&gJ@�t�Ҝ���c6��/"2j���<VV��@-�V��3!'''�>o��z��oذ��0��ly�\d[l���i�\`���2�+pC�Dͯ D:���!�NuH|G�nowzM&s�?޻lٲ����-~_�^��C�CJ*��ވzC�AdP6��0F��T_s�ĉ���#�iܜa�d�[o�5������3m}<?D,�z��Zo�+�ZO��-9]nɠ3�"bR� =Jƌ��UW]U�;Ϧ}��B�/۫WS0��.FQ�P�m[���dn��O�ZLR[�G���cǍ����t[���bC0{��� (��059ψ�	ɣ���E�L�DMz�L�0��СCi.�k:�����Z18���vHIbh�!����� �����ѩ��'��95E��i6��M&2�2P���� k0��g�ұ�f%e�B�-d4B��OL;J��1U l"�!�����^oK�u�o߾I	�ۚ�/�����$04�_m�Vʀ��"'<�
neq������~�nliY錴����3gv{�A7gX�m�w�d�퍍��3�,�2�~��C����)]7 �0`���/�|X�%M�I���h0��F���9�QykF����������pG�z"�G���i��DM��L�4���/����V�������u7�3;/�5�u%`
{����{�%u����ا ����\������cq�:
���g>Gu�'�9^p��������]YY����u��f���2-��G��v��5Rn�y�nAQy�6:���`k��
�����+�*�A�\��A�Ry���4k�����c�i�6�5J��A:���n1�LW���'ֹ�^��􀅉/))A���	����յ<j~"ޞ�O7Q�'i��&=J�v���(������C&�#����[����2���*����}����]�	��)��!������2�w|�n����֛�E��M���`��B���Q�h���3~�p#�2vH�+�S��t�-�)����崹n�������7�V��_�jo�(�|Cˎ<����g����<x�ƩS���Q�Z�9-V������.��+���>�D�~@uu5:�Z l�P��;�G�#C�NѸ�t0�d��A�DM~\4hP%�}>��O�f�6l0�
7,b!��;h=7����Ko/f���m�"�S�����qچI�iǨMg��v�]�G��E�@~��[����K�e��j�hnn_#�i/�����]�Xɑ#G骔�Q4ps��������3���nv�<��ӊ�����0�J.�[����MJJ�i��[/������O"##�d����s`����F�	�����'���J�8�HWab�Z��b������H]M4ѤG	9���֭�imm�&�}�[�3="��������2�ϾC���p��3��)� ��+p��N�NZW�ǅ�(u��n��]��z��6�z����u��fC��vv9*E6��lw]B`��Uݙ���ܼ-�hPeEŭN����yT�qcc!4���)� Q��4]8f̘5n��D�����{-fs=]_�c��mujJ�X�<�^	҇�7�x��_6��3W���6���nGM4��%0x������
��:�@�x��C�::�B4��H<}ТE�L=��wj@��Ψ��7e�B6�[�fO��"A<ڙC}.9Ru~���9�:t�����.<VYY~�|�!���X�x�^g@�u<���7�k�j�<x-��;��Y4psdϞ=��9�W555]��p�I�s:P����čܫW/1�hG��6N�2e�����G!p㋌���Dn�����s��s�/w;�w"	�&�����=<��SG�X:�ȩ����ݬxjZ�&��A�۶mU�����l��F��r�iv@��.�PoLUU����N��9?$�Ggp�?�F�!�ֲ�Á�饴bwئ,�SR���� �����gnoҽ�Œ��"�^��&��6��nz6����<�d7��e�/�X>��N������ؖm�ɒe�r�n����f��H�⊁9~ƺe��ܹsμ�����\�T���1��ر㻛�����n�Ze8���M<%ڳ�2(����!!'SR&�չG�y�6uV�L����A98���sIOOO)�� 
Ą��js��/.:�9�!.����'�ԋ�/L***���,����(	a��`	p��HY�iz��YD\�9?�����Ԇ����}g�a̐����5$���=t�>J�|T.m-�vVS<�39-#ZZZ��uA�cd/d,�ޜ�I9R������j�>B���� ?0�|>p��=�r���}��شi��^��*�sfD*\l��������Z��Ȥ֎��hD�tD7WY֯_�\�q�ͽ��qt1�4yM����\ox�i��a�1��x�JZ=s��*����Q��~�P�?�,DM��M�>i#.���E}�N��۷Ͼp��z�Ā�f��E�"�*��vr�SB��|>��������� 9��X]�1!G(RPPp���-H��":��j#����B\Z��.�Ϲh����?آ�_�=f��^@���؞@bQ��L"to�@p�I�d�\�
��V��ż_N#a�'ٹ^:�}܇V�Z�p���J:�i?����)*���b.(M�q����njl�O��������*
�R���;����E���ٸ���Nmk!D-��q���LFc(#3c�̹3����/�r�����L����� �F�5mۥ�{aORN�KEmmm)}��~�sHM����m�0�>�m����Ia up��.ט ����8��.���p8,���Nˋa���i����b8�S��4���M#�@%7a:��x������F�E�T�5X=f�C�N�`-D��C���EE�Ϟ�����Ϗ��X�}p�>����h2ά��+O)�.��K7WQ;�N��^����C����e�X�XN��I�zAg��3�.)��I�s#G�zu��9�.%�Ņ^���$�H�I��ښma1���E��J	�%学�Z��E�w�k��Y�s���H��<u�6���nt������^��F��H�Ӄ)�юŽ�kD]�ts�v����V�#�N&��j��u_jE�����$	$�&�/��ؘ�_��� ��u��}�6���$��n����ӻ�Nz�G���ןq8��>ZB�:c�/5տ\�}ɉx|X}c�=�pɌ�:��J��Ͷm�g����� 
��}�B�T9�� ��������ܝ'N�s9��gU�vf�\m�m���\\���I���0
�7�������c���5�GQ�}�A��3���x3H�����2�ꢋ.�����_K6`&=�h����\1��bB�n��i�z�V�<_۷�F�{����$	@�����ʐ!C,���0����i��smzB�#�D����?@3f�w���{��t��i	��ず<k�Ն�/F�&���3��x����O�����ohXB�(���fdlP��.8 �Gg$(
�QNgF���Ĕ)�V�_�Gm.Aʊ�{

�jC���5Vl����N�����~�[>��ș����ch�8�����d��m&��ޝ.��r��@A�@���%�uj@��^�w�kt=e�����j���Ӭ�����>�}��X��<x��Fn���l��
�Y6��(������p8|�j�~��>.���?�w�\c����A�����4����o4�D��	MMMä�@觃��  �{�g����^���ٵ�L����E�( i)�??�`��3v����K����XAa�9:��*o�x�AO�7�o3|�޽222ܲ$�#h���oL6.](�eB�q�}�
K����|h�W]t��RQQ#}m�h �-k�̐�2@=0�7@�G��Y]]]h4������}��>�k��9uꔛ�5��tڹi�#Ԛc��R��E݃>r$e���g�뛪h���;X���%���S�1$����𶎶1[S��.��D7WX@��ꫯ�466.
�B�(J㜦�h����Z$����B�����6m�꒒�nI�K�dAQn��f��oP�@���;�!��k��Q��B��x<Px����h;�=+�]񼷷ঘ��[�E]�9A���ۿ�Tpӯ�@�(������~�{,ل<��Y۵t��>4 �������pΜ9Ci[����g�PK�t�it�4��[�,Y��)S�4��w�X$��l���4p���$p���4W�#��Ӯ]�K������
KUU�g��݋c��P($�7_X��-LOU���Xq3�h
�ׄ�W�zLo��tA�ҦM��322jH��d�d%��9b7*�x,����pg�竭��l�F���}n)s	�㐬���5'��Ha�����F:��F}��MvGGR��A���;�&���z�h���~�L�n�Mm�ٳ����9��V>;��hq�'os@C��-��/(E�v������Vڏ��yv�\�#��{����
���y�r9��:�������M��·�!O$c
�~�=�%#���y2��j�22ܒ�����ܰ� �B���2a��իO��+�:��l F@�n$���Ѱ�o!���ހdKt�h�Z��M1:f�I���RT��C��_��l���� �V��;�l�.#��.��ry�n� ȋ1���xpm�� @�T�����(� �����s}~Q
�V�$i'8]kC�D���I)�?���r�0���'\�~����\���iQLl2��v�V�}�K�6��G``�-..n���UQQ/+v�����f����F�������r�%�řv�q�F#:��tlF�ƒƖ�2:�z��K):����{����=��c1�y`!�PC
!�4�a$�Z̐����t��ѣG��=��'yyyѢ����O� 9�^�#5�x���������_;9D��DB�׍E���c�J���]t��D����Fe��"��,*ȱ�~����"�r[[[n0�Ɛ^��r�^������b�p���D��{6\[[�O���f�S-"�
�1G��)6���664��B���+����p���Dl� K<�����'��m�Z Z9c���vK8�B+:��B������4oG�"6��Y!��!� �6��yT."�]���A�́ɓ����^�����W�X���#��,rȫ0�'�\���Pp2��7��h�\`���[IIɸӧO�׻�]t����2Az�T�t@�pH�vK�G�2)�F#����l�������!��+;;���q~���{Gж��ʠށ��;������������N2�+3��N ��l���]f'F�Z��皜h4����H �I�_4Q�n��lؽ;����݁@`0Ri�ZI͟&U���9 �7)Z:�"Y;f̈Z��w�����=7'wSS�(���tZ�~Lfp�h�j��q���3H]�/�̯st��m���-�ύkhh8!]~]t����QM��ϵ�F$&��m۶�C�Mss���M	x�����6�[BN��;??��|��={��j�O��Z-�F�~/o���wi�{�t�J(�gώ�Z��xKKK/��LL"�r�����5�x�`(<��I=o��:S�\A���u�f�4���cQ�!%�Q����ʏ+	��J)7U�<��r89�M�����@OW\��������KJ}{(�P9�B� 7Pv�AS�[DDϵ��<8��բ��e`�9<2 y#G��x����nt��K�� 6D����d��egϞͪ���a������؁���� �k�{�y�hQo���N��˷���1j�)��u��YYYMS�N�`pg��G���9�@�XH�6s��։D��xo���F�:�����c҇L;?���e�	����9s_0N�Z�#I��ȟ�0�=}�5b=���t:]�����O�<��^kse��k���^:Vy��I��W�,V<Vp N �Nx����a=��1NC꫱�+"�o������v{YY�2p����z�N]��ӃE���huZ+ZZ�)i�
�����1���9J���$�dK��^������ �^���~7���d�,�<�mg�Va����}�k$Q�w����k�X{���;�<D�q<�93�s�ݘ�
����=�;���s0�D�.��F7�Y�ǰV=:�.Թ�==���Ȩt�Ȃ�XJ�x�8P�\��b�6N�3����wʔI(��	����5�~o^���٤P&NA	E˾�w#:�Dt���u�zUZ�a������|����1�>;m׮]{%��O]�g@���M���x �?'[�)@�/~��,�Ԙ�Q/�xhx���٬ :�Ǝ�����j����1tY�"i'�smذ[�qL������P�j̘1�=o~���s�Ir�F�������ޚD��vr8�[�qx�u:���r�̙�����c�*���ۿU�`�F��C��v�֦)77w��)S���͕��������w���w�����' ��.�̂�W�!\�%r�����ц�9���Hͭ�n<t,�y���nt���<_����#�����?Hl'O��A��7KVI?a;��x�5��΢����s~��=�������sgg9N�6��/r��(v�T;����M�TUTT\�s�d���я~Zm�Z��d��T[w����|A &#�P�������(Ptps���޾l��|>��1Z��(%�H�Q6�Z�8����L�Y�u"��������t��6WX�;z�ކ��S�����p���AA"��x����7����� �uDw�Ɔ��g�����M���d-**����>������R��F]�!a%}��Y���Fge�ќ�vCM�������?�A����=~��4����O;����ئ��4�2H*�B�T�dɒ~�#D�������~9p����7N��D�Vy<�jL���sWZZ\w�lM��2�"�u�����~MLn�H8�`�/�/mjoʡ�/j��n.���`��u�uwweq�M:o���9����@�-�t�݀骒.W\;p�@�[{�����3':ٓ�V�C��.�xڠ�7K���7@�º�iefN7�h�e��'`����{�ѣG7�:z�N]�!gC'-�|`
��ׁ���ـ !��կƓB�Z�j���I;F�4��6dC��NMyyy��m����\YY9�l�p�QѶ��mB)��6f�·�vɤ��u�L�sC4F�0kSS#6�z&t'���N_���[7�I:::���=|Kk[�X\���v� ���0��mĨ��HYY9)������5q��=�>��ԩS���m����~?y8L��>.��sDc n�::�5��z��de��,Ɯ�bC!�Mwpz�9-����SO�>=���x��t�E��M�Y�������� �6%���N%э<Bv:��N�ɓ'�{��Bs0[�{�)/��N��II��H$%S=a�Dyw��QRWW7��tdq��v�9+l�w����l`;٦�iӦ]r� //�O砖l����ߍm�8��A,���|��&'ɼ���܋ݷn.���X�e��ֶ�;�F��7?���^XuXXR�k�'jm��ّ#G�7n\���Ut�޼�DՑ#222
}>���#]0�u�Z�H�7���^�n?n��	��,�ޔ�q����!z����E��O�m�f&�,�Ŭ-&f�r�0 I�ͣ�M�OKeee���^&shi��3cp��F�K����rrr�dee��)@���}}f"�Vj��@�|��a����9j��G�~tb`��b�����a������m��1�q���^}���@8\��s1[:������>q|^0�HJ ��]�����<7L��F�E���ࢊ��d�#~@��i].N&��ж%ۮ`�7�@KZ�E�%�����.W2�{��&γ�uDo�0������� ������)�Ν�[UUU-]C�.��riB����D1h"��;�����v����f�f�o�J���o���N è��r��kRvN��I��RZZzv ٵkW�}�n%{RD�70�т&(�Æㅍ�"�������ܹs/���9S�����>�~�������1��K4)��J1�F7�(@�[��:������n1f?.q��H?�@�))=[��v�;)B�M�F�Y_VV֨{�W_JJJ�ƍ�����x<����&������Ey�p;����
PP�����Pd̜���]	2��H���m�Ed�m߾}7]_��׃.�|<���j'�.M���o���ڨ�eq��^�%�n�mۖ�w��Yd#�Ѻ迶EZ��JG��h2y�"�жjժ�6q?���������P����|�,x��������q-{.\����}��Q��~�����d��վ�=�_�d�p8X@��tps��P���p����Q����oh
�����8���qc��_�Z-����wǍ��ֹh^].^�ؕ�����<�� �26�St�V}�E�Qs��)� ����#�~WDr ��V�%E���`�Ñ��5;;{2}��͛7�����r]t�����Mz�G�i��Xq����-�$1Z�����}k'7n�8����sd+\t/�bI�O0�o�#�O�l��>�w������_��^w׮]Z�{� �WF�����1���1(�8�	��e#%��o2;t�x��Ҷ���-����X2e�'�^��(]����(y_eeA}C��tSsd��QtҘ���⸰�tڿMF�����N���A�J7�3�S��c�����Jwm������$R�~�b�V����`
>��.9�nph�z�fc�W����źMMM�Æ�魷��u���m�ڒ��.�\� ��裏"�̄�����2҂~�Qz�F�}^�P[[k����g�-a�)u1 v��遘b{�GhA�Z��LЩ[o�5��P����nrMM�<:'wx�}Ѧո��C�Yu�z����2/g�8777L�����sb�s��xi�C�o2�4�)97b�|�E7� ��ط���@`f(5&�)�l�I�8]�&%�K�%3:o�E��xB����.ވ۝�Μ93wӏ�t�؄�������S5;B��Ho��4���(�m��0�^
HA!�5���vl�8HFN�A���|B�y�ap��jUxs�`����7�	Ń�g���@�����;�Z:���t���IUU����m�/��3�H?SJÒpP!`0�5����ȷ����\�6?��φ��ȕ��m�XF�)�����~Tz	�G �V�WM�8�J[h����~����gƺ�n���d\il��`��;$�Ն?�T!�F �mw�M7�y��'/�y$�=j�[ϚL�(�*;lj��I�\c��(
%�o�k�p$�vGm�_�\�����476�H7��A��˗Rx���F��)���D�o���J���9z��t�$]>vA�fȐ!�跽�~�������ݠ�&''G�~x��L�M���@u7}���Q;$�Ş&�b��\�G���vg�km��,[�ׇ��E��$��w��Ʈe'�6h���B�"4,^��=WM�6|�j��#�o�H�^GSk���'�O�x���7cƌ6�v��׿Nhii���pd����;�ũ��M�#u_a�����7\�.)��={6n��[�y�j�G$\TM�m�B��/Թ���E
��+K_�mo�,r70�z����~1;�(6`��;F��qg��]�''L��7;;[�4�ћ�۷:s��R�")v n��cx>�����
0#a��'�R����.���>������O7Z�6)e�+.fC�;dl�oavvν[�l<�{��s��љ�u��
���/�8���5�t�"� D[L��V*X��{^��o�j�ﰦ��y�E��HC�4<4)M�6����C!19Og���K_�R��_��X�رc������BN��?�\k\��C2�x!���::�p���馛��x��z.Q��v��N�5�2c9_zJ9)t��8'��@�n.RN�:�]}�Ԓ��7(�ʩdLBcTJ��$1�C�ɢ<%
�!���v�(�j��KJJ�:���O��fd޼y����k�������<P�=!-�q -.V:%D��0������h��-�t�R�3X��ˡ���H�2���y��W������������g�Z���&�������ֆp�J�A'SAAA���nڴ)��7߼�ޛc6�,"��h�c@��[K�ZZ9�B�0p{��G�>}�6��d0��r���x���֋�����n?��_�2�����\�8����݇���y 7��Vu~�h2Z	��UUU�d���J
�V�\Y���:#Z㱈�@�E���M"�(R"�#nX�A��L��rf %�����Ul�x<z��x^o���������)���#jox���(�+,,�QA�OD�H4$�TѨQ��x�:0&0"�2vQ(�����G�2��<:^##+�3fB]ݹ�_~��&���C�颋.'����mmmH���ъ���`���7�"�=INH`�g_���*ȑY����K` ��4�v���沆x4� Ҝ����'?����?���.�+V,&[1�l��[���D|a�p� pP+�))Z����I�&��Ru}�� Q���}Fj ��z.L�D�M��;�tpsR]]� �|3���]�F�PE�Tӟ�(wI�FT�'cq�I74]\tF�7n���N�kLfΜٶgϞ5^�w!�2�#%�^"-���Rv�G��z	��HMR�����%2r����v�,tD��@�f��q��Hq�;w.c�С7UU�?�����-�.��rE���~p�Ro#P��|pW��l��uW�:J��nr~�����E���立����g�ܹs9;"i��Ǔ�~L�LȑlWDv�؆(=?8y��*M������f6�ϑ�qq�>������`� p��Tx����>�w��فg�}���Or�c�l��\7i �a��x,�����n.Pp1m޼nTSC��tQXcHG$��b�R��RI�h2�I��	ɐ0����F�Ùr:��Q#W�Ŧ�^�B�ݺu���ƕdP�A�u��0�'"1v�U�x����{Q����Hmm-Rv�G��pâ $��1Dk8��948E�-�0H���=.,--Y�s���ի_���b��.�|V����ݻwO#gd8���)��tGt�>�3�m�^����<���3gθ���o�>w��fs��E;�Ee� �Bڗ"@R������;�l|��g�m�V�r�ʻ��h��cD��bP� ���) l�Ώ�����~�[ߺ�NvQ�K���
�~'��e�2dZ�)�M")'�q�@�":��p1�<Y3���{nT��r�HH5�7*���e��	z_U�l��Ns9�Lguy���H�H�\�2���cǎ�ioo�K�c2�@�b<Rd(�RV�G�{v`� N`��#�r)E�x�#3Pa ���e0��ul�!���:iԨQ�C�Y��s�D	�s��9I]t�lB6�S__��tݥ���)"~�힂N�I1.�
�EV�y��555�� ᡹h/gr>u�/�]��Ǩ�9:mڴ�܁E�5��G?�{������l<�J;�I%Az��FU���Zw�ĉ�hiD"aJ���W���;���Gg��1z�^�\i9~�x��C��'���4��M�`$��������"�������s���`��yy�ZI�kVP�RYY��'V�"�455�e<��� . $�*((H�����46��RRR"����Dx����:NfJtf*���dt�aÆa͗�y�)Ú5k����%]t����W^����<�l��6ܱ����و�qW�;^'���k��Ǐ��m�����'?y��pL&=�����5p6@D6�^UǾ u�����e�7��ͳڲeK��+��}�̿\���q�	��a��~GG��-jD��� 9LG����_Q�5:MI��F�plZ�����_��J6#�}�����=���+Z[����O�_�Bt�1�0Z!"�8�,�}>�bWr�h��t�H��fԨ��t�wK�\�#5k֬76l� b�{�0XP+�`y����"���DG�a y�Gw�Ǌ��t`8�Z�4A )|�Yx����5����u����Y��͗>�����.�\��ne�:uꎮ��b���n�F;В�w%A8�K��F:}t�̙,>|���C�M�|{~~�c�s�۴!�s1�Ne@�6i�
�n���rڴi�.\(",mmmh��;���n����~<<��o<F�A���)/}f�M7��t�ۿJ"a������x ���{.h�57WX�y���{��Cbֈ��D2(�15)�1bQ�FH�d!�M`�bIy�F�h��E�xA~޻��&���5.������VWW/'�w�R,��B� ���Q�����X<"C~2Nq��츤���JO�Z����¡cDq��� A0\��c��744	H�����_L9�$�$]t���81uuu�	4Xy����~���iu�.�m���83u��8�@?��g<x�����|D =�	��mJZ�̠	�#��N!�/^ܺf��u����fҾ���M�L����v��#̽��V�]���q��U����|=�G�(����|'H@銞[�)���>�a�.+��WZ:d󶵏���M0E&��u��,S	��Ź��S��21D76L��9]@Ϣ��l�ȭv{v��i2���4�~��r֓�?+++���C6D�X �{a�����X�� # (�`D������Z@��l�clޗ2�Ӓ.4�"�0��%����G����_y�'[�n�����[��J].\Ξ=�q��ѹ�c#�]��ݍ�<$=�̪��t�t�(館�y��'g�\������Y�XxH.�)���?�M'�p��~��t��vvv�Cz��+_���ڻwo�sy�[�x|��Xq
��@
�(��#��U:�٢v�ٺ��{�j�J���.�g��=���aA!1�+3��o� :�� 	��r*)��dB��d���eLI�P@*�.�J\R~F��{�+d�Nw�Kq�U�M�;�%������;:��b��O��D�������������x<����)pR���!���S�4H��΄���%555 ,Inw� ���{�Ŋ��a������5��X�c=8��$-�n�~��m۾��c�������u:��E��S�NM�������L��Ȥ�7�'�͔$ �Lz���y�|;v�(y��g�O�;����u��s��I�bƓ Rj7&�GmHh&gf��ŋO.[�u?���n����j����\��)-N��	�s@��2��i����óg_��?�A�>x�ϭ�(j�ږw�9ն�k_S�q.8%���HYA~*�'��TJ\�f��g7J��O*�vKC=ْ)�R���ƶɟ$��(�������+��"���ԆfggQ&���E��� :Å� 1L��C�bb���b��?�`��Ɖ'è�;�`�`(��a�Ǐ7͘9��ࡃ��?��G����}�^8��������|ggg�	�n�ֶjk��	' %}=9v��C���G}�n��9���nԍ@W��\�+F����b�sY�%E�jm�c�6��0"����o�nٺ�K�5$�8N>�a�p�`+��B�1��d�+c�m���p��@Q�H�g��LӇ��h�L
�p�}.�8upsb��%��X� ��9YR��$��^��IE��1�H޸l���d�PJ���S��pdz�F�(;@/%]>q2~���믿~�ƍǒ�����)��Pq /06ø�(N�;,`�8A�0�<"m%&�+��-.����<|���S[[+RT#�������W^y������^��	"u����nݺ�'N���@�ū��8C�i�d@'�9 ��s{�O��}�g��}@w����܀�@��� ��r�ل$m����p�����Μ͛7Y�ץ$�)h"�t���BĆ`W8m�}����;{��mK�,�_�s���d
������2 P�@B�b�����������Qu��?f2Hvg2&�����R��.}~)�f�8]���+��:�D*�p��1���Q2EI���}��w���4E� +��2��J��^�k��Fe�����O��pdF�A(<Fʋ����	�U D0l0�X��L�TD���������g	���Ϣ�E�������={�����<
t�� ��J��x�$�!��|4�z���@va�޽{�C�% �M�>��E��A���TБf��)Z/ r�{�wÝw�	�O~��/����E��DW&�:�\�k�&��f'=֥��Wد�������T��cO^�sL�b��m�b����I�o�l.}6�����\����%*F��ط'��s2.g�,Ҩ�R��IN�YJ�"�d��a��j{%�䒲\�R<il�[���v���`A$�0ISS�K0�o0�J].��FB��Q!�C HxN(0N`.L\���1���b tO��Y�	i-�hQ�mE�kf�U,.�3��0X<w&H��LH�����2><�޿{۶�P(���ݻ����u�彂��SO=5���z�SG>��7
�kYL�� '���ᕒ�ӑXNZ�3[�Z�nji6[l�2�V��"s�/��X���`�&���h0K��_8;>������3�ǎ^������Ǐ�������,6s���0�,F�mi�> 8T�u�d}���X9%N2�-;Ə��c���Wu�!��]��������b-�
zRKt����(@���m˭�<:�('��q9��}oK�Y9R]�6��IQ)H�A*,&uwI�-�TR�|.�{��Y�����d>�6ϵk�.���D��e��r��v	�S�O7�ܠ\����"����QG`��8f>f�����\��A�9�"8x������_:p�s��ۿ������+^��]w}�E�n�KZ���7�СC����$=wSN��9t���PW��t�D����D��� �!R[�hZ���q�\*��bQ��x$�*Lz�"���n7+���-�{��g���|����>���d�� _eX�Q#l �yᴙJM6�ڡC����|�Uo8������ą�J�N�7e��U��E�PNN���`s����W^Y�����d�:Z�j�L�Y��8%�L0J�q�H�ڑ풲���T���^��V�w��<z��FI�O��r�-�gϞ}q���IYo# cQj��aP�q�����Q	ӘR��E~�����(15:�����s��� ����RÑ���III��#�鹭�"{�<N����涜7�X[��}����ӦM��pt��KKK�EħO��E:g�x<2���,w:A��T@�ىɰ�8򀈄�����`V:�6B�����!�
Ń���7��wע;�Z��}�k����	��#�w,m�,�m��q��	@ac l8�H0���>:�u7�����]Q6⁲t�R�֭[3����g*p���z���>��zA񕐚���g_xᎺ��*r��ý��:W�g���Mm_4�d�$9s3q��'.�������yc�����ŝ������omm}�������p2T&t?A���6Q_EFk8r�C�MwE�P� �O��ap#F9�,�,��7�	�Ց&�1��Ɩ�����B�����嫫W��ii��������j�t��Z��^|��)G���t1�t���3�uč@:�u6�I����p ��A��r_���H�Rg�������p����<�d9�ʪ��������1ޚ��+�t��3�c_���&`5J#�tx�ؑ{�����^�s=v�X#��\�sN�������Z�C�ŭV���OB�@��͇H��i�^�}��'73c��l0�-���K�T"�l��F#y���ಧrJ����+�o���f�;bܼ�|����l	BO���~�r�o�wT����	f�U�����*S~E�;�Z[���c��ϛ��X8C6h�C2[��>R]!���gBG�sWg�4|�pSIɠ�3g�|q���!oj��ŋ��4�.�5A$�ݻw�#9�	��+�M}?�kX�Wx�0�Ӕ *V�Y��xH�<�y"���bpb��*��;��z�D�n���@`�=��w��\x�_8t�Н��<:,ݗ\4��/t�mv�4�E�7m���h��߾�ݏC�kjjL�]�b�sN��L)>_��b������RQQ����)�c�,����u�vn�������LWf4���8f����E�������H�E)��$e�g�2���C�.�i�FY.�۾?Ų`�������{����_&��CRa`�&%}�5y�6����Q����u��9����в�K�[� �K
�<���۲�mR]ݹt-�G$Gx���t��	iĈ��ɓ3O�<9�С���Y}}��>��T�|����*kժ�-����鑋;��c��(NGTDa   6�S�t��f�Ѡ�N����;&u.GtT�����������΅oZ6c܌د�녛6n�ف���L6ۀ#�uvx�ǈ� �p��C�_�
Һo���W������D߷�������_"�fbm���z���_�~up�>�9#/=�ԔM�7K2Jӌ�5�eMY��'3s�M'/k:����Iť��n$v�����6K0f2u�"���R���ƍ{�ȑ#C��ĭ6�|
Ј���9=$X Di�K 
��bءh� ϭao ���4!���RQ�ں��GD�Y�۩�o��fs��G@�:y��s}z�ҥo]M�]t���,�l�tˑ����3RL�*k�*0�@ �
��]T�,+��W&w�
�f�$�Ǚ���p�ǩ09��E�o4�+ڝkF��b��)'��mܸ�[F�q��e7��8 &�E��Vr��HBԆ����NG�ȑe�n���Ə���@���'�G̈b�.��X�!�!��/�	G7� �W�}v�����)]8l.�S6�Rf��+�m��}�������x��0	���dϰJ�]��ϑL�I�;O����[�'��{2\n2d�;:�vx\ هa�������������!�����=���P=�s1�dưM��"�^uu��}�ν	Fҭ�x��/r�Ep�:q�j��e?�����7�di��2�˧S0I{�ƍ�ߴi�wSRr� ��@&�C���3��o�aD�L Z�rf8�,�Z�? ]�* 	��9TY�_z�������r��5���_}mُ,f�,Z�Ɯ8�ʁ�3�8��a��6O�VSR(ĭ#'��E��;0v�؋"»B�+��7���J�Xߜ��3�8�N��6-�W7�C l^x�1V�������peĤ(f����o=���?9����u�f3�9V��M%�h�J�JO���ڒ��9n���gB,X_�~�a����WF�{
y,f�k* Qڼ�Y566
��؀�d�#z��ia���0aNl��+`���a[��y���ؕ���T��ۙ��Q�QM�h����ױm2����S#h[_۹sۘ����W�\��;�躘0�.�\�Bz`y��f�[��K��Pg�H*,�\��7XD�Ox}�� r�3㸨W�Mc:Ŭ�Ce��Ĥn�]�_�=��a=5��
�"�]��-�c�$�/]�ڷ���f�.�s�A ,�u�8O���P����<x�̙s	��x�?������8N�ݙ�����4�	3�q��s�̋�W���F l��G'�[���N��֢�O$��dhPN�E�����F������޶��P�͖���U2fX�=��f��j�I�|�d���;w�_�l����O3220����*�1��a�HOA��.�F0! 
ovv��Ŏ���E�0l�XX�w�6��1�q��b[�ހ0|��\�C��p̘1&S�t��74����O;|���>>I]>�.���W�oذ����]7����; '���z�(*�8��t�!-�HGf�m�%�{J�1t����=���3g�|��`pj��_��캓t8�7|�p�p*=1��c���ݜ��i/�#���!Ö�����QZٶm���s	�C�7�PL,yF���1������:�ߥh�y�;���]\7؍�B�r*�V�e��.��=t0����C2Z�q�M�x�dvɒ��)ٲ�R�"���O2�����Ϟ̝;�k�ҥ�H7���-������2rA0�n����CX^^.�wR���qy��!��B��\�N�%��l	x=	Z��� KYY�d���5uj�j���#���H\�Æ�;;;mmmm��ڷ��MM-�?���7̝{S�^p��4̈�  �IDAT'U0�qժU׭[����s�#���i	5��|0 �p0r���+�u�K��]L`X�Q��N�������m�ui��?$􌹪��h���^�;�e#�./ֹu��5��~��A�@J�i��t�-��[�הh�c�[Rq������3��%��z�{?n�a�5�d�r4�5冀��mR��\� �銊���?:��T`��#��nZ�]wf����t�;��T4�;b�Н��q����p�,�G7���S���%.[�?��dGD29M�=�Fe)b��,s@��:��gTP�K �͕+W��bѯ8�C0�O� �L����b���{
�S�N��I����Ǟt��.�U S2����R� "8�4!�Ëu��"č	�����E�0�<����VL?q��o+W�ܢ��t��	"�[�n�b������ܜ����z�e0��,� 7���0:�ZDC�0Ew�(Ta�s�E!҃.a]����㓘?G���c�Iұz��7ǌ)o�w��*++g��d��̑����-�S��͜;�+���|����h�o̞={�Ǚ�b!;�
����:T��~39�3p�uS����M�>~�"����_�����zk�?�.Y`�;<-�M)��ܚ_\�yɽw=;���w�	�v��g����t������D���PgFB�[#R�KIo$I7�e�)�+V�����
�3ZŅ^Ó�'�]�n�;4y���X���hB��;I̫�R2�FN����2jz8��#��|0�N�t� CH�y�^3�Bw�XՔ��s3>���ݻ��hv�I]�uI�jm+V�(_�r�O���X��l�˲14P����݂. �C $�?��@S�"q�Y�L��x�i�H,M�	�B)��$ up��!MǪN|����w��� b���`D�-9-�S l_�����f��8E��O:�iҤIK������ߐ>n!��O�6����d����tGs8�M
����t_�?���Nd�s_x���gk������&ey<����d4i]6r�7x�O�'M���
Λ�y�d�����L�|�ٙ��LY2�eIr���R�M-R'��t/�3, ˢk�l8l����[L]]�ȫ+��{L����40� #��,p`@����E��A��Ǔ��2p��xc��1iο���=ODo��Ry5�qb}�ŁQG��:������2ȥ���铛������o�}l�̙>��r-
����_�0g͚���z;n&p��� �|SU�Y�$�U)�ō�Q���N2���S��UI3)���}e� 6�;'��o��)�"����ȴ466���'����t;�D[���9q�Vxa�xMD�z{�_��<��)���������7�p��k���������:oƾyR�`�~S\����Z�|\t��gܬY�����޼���uIɠ��d����(nH���Y���E>z�lU=���ގ�/��ri"�k��P�'���c4g��n2�0]�ɘɔ"p�&..]>>QNK$��L"C�}��!O�#��))*�Ƅ�'e��G1�bP��tw�ȸĘ�A�F�,&�ܪD<&xu$������dH�!%�2i�F�!�����8�#�t�=m���t|C�~{��'�6TUZG�����To���{�Z���u�6�S ���p8\�l�����i����PjӠt �-RTL���S�XW�%t�@��6��*�܁	GU�#&��l��s��'��:N3;;�{Dry�
��|:x਻�+��uP�G�-��s�=�s�̹&hH�y�����q�!-�s��m�Z�b�N	��-��{�����A�����i�_�{���ޛ�)�L��A0Gjg̙���������M왶nx#�����[���f�dsڝ�`0�;d���hv ��N:eݮ��AW}H2ڼ��&.0]>^Q�R��֭[�$�EnU �*N���[L��B�"8pd��--m"}��o�m��[�Μ� )�a�[Y�C
��� �0K�e ��>�xMrܴ��Xt���;�ٳo��/��e�С5�g��]>.�H'yϿ��]{v��f�Kzc�kZf���U�@���dJ��^��%n��� �� ��p�u�G/�\�<8��b�t�7�:$�4��R�/�@ɤK6�~I����l�o�!t�;��m���I��0��l��p��O�~��	�\3�����T:~;����j���c�kSV�@����V����3n�;�z���N]�~�Wmv��Ņɘ4�twG¡����r����濔����Ϥ}ny��l��w8��sҔ
��~��A�s'���=vK��`#�i´W��\�&�L���"q����h��[o��$�t�۝��v�I���!W
~;::�ad0#�(JGG�ʂ:DDWx��bw�0�6�EtT��}A������:t�HQ��w(�?�8r\J4)V���#�����A�0[h��x<�
ǭZ����ܼ5��ջ>\����r��}�JW�\�@��#_��ʬv�E8I�X/P:��v���8�J�@|Ks����%��z
�݌�p+�K��lQ�zʅx4!t/B'��"�Ujcb�0��pf,�����tLv��7���8���{�t�c0����K����y<�gn���(����|�gPo3�������(�+��>����F�b��$�XWQQq�䃟p�u�Vף�>|gSc�9�ٳ�ƑE�YnnnY������?�xÂ���6���ğ�0,�ٶؖ�vۜƞP"�XN;�UkQFe���8��>�`�R�S�5�2X�6up�KZ��f-����}��)�=�+��+3M��\������6L(=F,�6��A�6J�TJ,�XH��qr8������TRRJ��.�M�噃C۪�4������� 3{�=E����Ohii޷gϞ�O=����6��*]����oٲ�+v���O��N[�����f�f�;�@���(545�:7��aCJ��z\@��jb�b�x�R��N� �7�9��i.0X ��N���clH����a�'DQ����h,43� ���t�1o޼�_��W[����I׊��c�����߃����@8J�iy�g�c�#���A�t	��O=����'�_z�{:�ڿf3�F8�P'B��7?k�ۋ���ɳf�����W�Ա�o�U������9�l�]�_�|6smV��K��y-b��Jy�1�C��F�@�f�9i���fu(*�9B��k֬	�A|��A���g����e�I ;����(�'&<R&��v����t�Q�c�ӌQh �i�d���R�Y|.3�#�/�Cȑ���l��������������޵w���Ə�R5s�̀��\n��y��9������;v����ֶ9tS̴��ɀ�<t�FL����-^G�7@w���T\�ڔ�e�I8ݺ�D{�b[x��E���S�y���d.���\�,"3.e^�ٔ�9p��a�@��p�#G��i���,�9sΟ���o�_k)�'N�����H�̍� 7<�灇�B�13�߱:77��޾h��7�O��>��CSO=r,�� /��f5���хw��|�ʻn�g�ԹS����׺�:�޹u���0�v�c��9F�M�D��·F̜�V���ЉG�t�He��)�=I�$]_&CP�t�3]�+j��)�o������}d��oj��e�l�aT�>j`��G��G5 t(���P���m�A��
0$=����S�M6�����b�0����*�,Q��=��}Ho�=E�r{{;�UE��\ү�7n�{ǎ������ۛ6��***��8�����Dk6m�4bݺ�w644~�������ź�p�ߜ'&���P ��Qn�� 1 '\�
���b�!��}�����ǔf	�0{0�����v8��z���沲r�ݐ�>��|T�Q��QPX��lԨ�|���k���y���g��Ϣ�g@����>�������y�����R�ۧ�,]�������6��~�N�₢�d4tx�B�tr��O���+��5�ϳ|g��q�������0��,�S���v�L�,�`l-Nz�?�kJL��K�e��H]tOU��5��@J���˗'|��l)�A�x��О�H���p����Za�����p��n�4K��#�J�D�����j�K�Q��M��d(ɂ������U������t���&>z����|w��!H'ߝ<yr��͚��'WP7��SOL��΁/�47^J�m6���$R}���C�3X�<5�ۑ�?�M3���KR�9��y�����	�(�|�(��� ]�~`]�S�����a�Tn�J�2����yl�#
�U��,))�&�Z1~lşgϾ�Ե��7�xcľ}�n��3G�����S<NB��y��A:ߧ�s��}��]��e/�e���B4�3��(7�����H�%ӝ�kѽ�?y��A��GB�ӯ�j�m�~v25�n4���M�&bM%c��8~椷���v(eN�l��l$,C��'ɀ�U2Ȓ.�|��]T'i��Ν;;N�:�MR�2�FY�v�LN�g�� p�#:�@<���[Z:D x�LȝT�	���҄�0�L�	�f���ž�c#Μ9�	�� ���]nmm5�{9��Yt|S�ގ;*++Onڴa���_;g̘t��`����,*�]V�|����8�l�2��������D<Y�n�x,)stM�=�����@���0G�e	����Z�)X��p4E)썪l�mTE��a`�]@ʼ7;���1�B����;���^�CǙ${М���f�葏����|�El?�������t�.�vq��3�;ošs���8hР×:��SnR����?Q�����{;ۿ��t.����Iʲ�>߹)3f��p�o̘1�0]�4Z���ғ�w�c�,/��N�:r�����A;�V�]-�]��u�Vc�l�%�r@�#�d��$rqup��G��j^�b�32�uuu�b�"�`��l 9�C
ëN�]mmm�-#>���.)��,%	r�m�tk�Rg Т̲B���*��x�v)7�& :?�|�
<�!���h���A����(��6�\]]-Ӿlt�CȞ��{�wv��ر����>}��]�v5]w�u�,6]�#��v���'����G���n�ףN���Q�WK�t��g �qC x@�Ƀ+�!� L��K$,��h�Vtѹ���DR��*�ߟ�;�tqR��d�d0I�*"��֏��z�,
#��[f���ۼy��$�l���yy�����p���\S������9r��tl��s��N��Nz�031�v�C���49J��� 7[�.u��o�=w�v�Y6��t�G��rƒI�tf�����+�s�ʢ"O��8־�ρ��{W,�Ė����E��ʊ�׽\8&�Z����J�qD��)5:�>7�r�E��(w�}w��o��쫯��SUU�=R�2 &��8Np��1�cWW�D��!�ϐ'�s䇽�@ ":CP����~`��}�����
�:�_��| ���Y���xVϴi��B4���Bz�M����c���ٳ�r�m۶��_�'�ӭ��t� 
��C?}����Ͽ��št]��s� X/�X�wr�E��'"������d0���Q@�ԑ)�T���=���/t�P�����FIa)���&��s��(�� l�<G��J�~Fd:��<�@$����=#��Zy��?��]�`�5ǡ�l�2�={й���I�| 
Un�tm��0Q�yqF�n'�wɔ�Xp�Xee�}���S���En�d���N;�&q��`�n��Q����_����d��[��/{�m��Es��_<fK1�|Co$�[գ'��c�Ԓ-r�m��n"H��T$)2
�I�R�\T�k_f͚�z�����H4>|��I�g��v��a�%=LwRq�9�<T����X�5*=��ۼ�a
�*�l�S�:,Lc#�m�̷����� �hi�q\ؗN��yr�D}���L�^_��~ҍ�t3;�cǎݿ���L�<���	&D.vp�.�<�]߰a��ta�o�����.��ib*){�@��[�U�� ��k ���nK�����d|Bw��t���ruEŁpz��	����@@���چ1���&�O �c�Ϻ�b �e����4��sbB�xxȐ�3�{/�?��_����Z��۷��y������8�Ā�gF�|)��t��%�\�������&�!����_��fͺ�::�6�m�99�e�"��/���/�~����n1bD�����gW��r;��_�L�E�8��1oo�v��^̛<a�\~�{��T�F�F�	�X~��.!ӦM@����O��&�R�[z{{=0�ඁ�C8]�.�tP��¨�P�H�}��[�� ]��|��2���~��硝��xU�.n &l�b?��)`�6K|5}��qa%GrP��.t������ˉ��d�� �,@����=zt�o�Y5v�؞��2��X@�˥L5����GC���u0?��$G���9K\-��j.���l ������C�Ƹ�9���\b�ө�y��*����\�ܦ�0+\,��<�����v��z�7y�#ǥ0ӱ����\��ְ�IWZ�0q�ė�_�����t-�֭[mO<���m��91s�3��2����Ӆ���I�w�#;�x9��n�D�ׯ_���3��l��[b��D�'+߀���6����zd�����0wM��ٵy�����w͋��֬�����a��V��K��h���?W6m����ϛ��G��6����knt�h!��>}����<�ڵk}dD�"C�K ��S���p��b�J��2��3J[w�t�d@a����Y��������q� �Ra�kxD��$����f"xr���
��`I��w�T�GMY�ȴ&�[i��0�@ѭt����?E�}l�С[^����ÇwN�4��NWJ��t>�P���/{~������#��st�L�K*��Ck"�2�u��6QTڧs�ӹE{6v.PU�J"J�7�� t`@��1�S�}�t�GIA)�Բa����b{
��7]Ǧ .K����(<���ڇ��J�:�)�� ݈�5MK+*F?�����Z���z��ӻ�q6�3oGm ����1�D�0ӋtQ�8��Zrb�/Ǳ}"���m[W��_��u�N�\D�N�#+ϝGW����@0X7�x�����oL�=�ć���#4�ZV�{���9"��[���V���Ǣ!�p�d��'FΙ��<kV��m���D�`��٨��GF��H��r��֜~�W�����k�z��n�d��?{��ue�ު΍�� � 	�Q3%��HJV�r����Yl�����Y�y�{�g����=Y���e%R9���H
� �t��gW��hQ�d1 ��X��]U]u���}���"5f��89�,# ;�tmsx��(��Ch����[��0S��ض�/�혱O�$������SA�8<�o����rtϜ��a �>�
���	d�:J��?s%�c6ms+}~��ݻۨs�M籕����^{�0��ٳg'�+H@at���k�z���_�����#���eLq���Hw\(��=���M��آw��}�0!A/�yS8�[{�}a� 낲�*��'�����X��@���`-?#�h�d���f$keK)�c��i�Q���	�X��q��'��v�kj��4�������777���
:~O�X��}����\�5�hCj�Tyyy+�ݟ],Sƨ&7����_����r˖��Q�"��V��[��RV���p{�+�Z�­���*1���o��7������n��ɀ�M������8ރ����1m�����G&3DӁL¥ѭof�����!r�R�F�#㳟�lܿ�Ж���Rz9�����2��`�Y�=�LX�~0�"2��	���~+a�Ԍ_o׋*
	�+��b,L�H2	ᬢ�(ҫ���Q�k�h@�9p�9:7t���?~����a�A�㊊*�XA�P�m�t!�~�7�c�����蝨J�}���%%�����-|��is&�%ÚJ8�`�O�|0R��o}����m����պ�ZD�J}]I���F�Rȭ�{���&%�Dz)K��vU	�Ⱦ��F��gE��*�v�u�z-hgNf	���v�m�d����%"�Ù]��&F��1����6���m��ͤ�:RYY�#��r޼+^��׾�C�F�V`|��w�;���
:�Rv�FPvS��C��]�>RX�U�����0�}�iN��1*���_/���~6m�损���x܍��>�[��0i��6c������N�}�n��طv�j�m\�י��Ϗ+.�O�z4��D�d��)�:k�u�����h���p[���=���L	�%>"0�#t�y��c߆�Nc9u������t6L�η�qȈ]U��5�QH�M�8��p4�~���`�0q'�BL�3c�Lv�,�r%ft�L����#H�7�B�{��3f̰�� �*��P���N~���ڀϿh0<8�v��{�֭'|���R?���������U�N�~� m׿|�rt�ʍu����'���*>p�@Ž���44^a��t��}WM��������b튝��4[����8��ɷ���294��Q�?pOY$��ɖ&�~�䢟lK�?���w�:S ݈��s��$��m�B
d�3�~�+��g ׈�+�%�w0�{�Y}�����,x������b4�g����Fj�9�F.�|-�p���Q�x�m�[�ms��	=�g�80��45�֭���Ǣ}��\w���Ƣ����P X==�tD&�����\y��G��r��UUU���|�	W˯~~ف�������UM���m �쏧��Y:��M��yA���%J��x
S:Q�M+��G((�8�q�n�W~��_�~�g�c�u��y��ɴ�&�Y�-6���={Ei��B�ftt��%f�4��ޞ~�5�|�c�ɳJD����pqN5�����.��^v �������D��� �A����#9 ���Uܐ@��M��SiO������i�L$⧢]�����������C����;wn�0aұ�7�р���r%�J x��.�S�N�������ɓ�������B��'�u.����а���ZJf]�и�~�`�[�E���l���9�]�e�-�N̥gC�q�a��c�HH$�"w��X"kY��_�J����A<X�ܛx�4�����,)�c�,��s@٥�J��Ne�"B&���������O�������x�h���}�ߜG��:�2:��91���,r��B���\��P���Z�DnΊfuT�0|z ����ݻg�]�O_��x'UW��ɻv�4��ee�{n����-^�d�i�N�ׄz��з��_�������t�β��2$���Aͻ~�����׿�M����"���#47���ͅ6��QS��قS���A3�4�DDd�~���ڝ|�1�ۄ!OY�l�.�(+��J+�
b�#]���t�*x]]�e��*: �x����m��e<f�Lr8���B����Kdu�vx���L���jll�F�tw���f��4ϴa���o�i����!���#����#^��HA��]UY�ZQ]�wժU����1 �U�?��o_X��H�w���ww�]�F/K��3L�h�Uj���{�zj<��:sAH&#EYk	��}i[t��O�Ł���b��ι�lwQ0k����R��p*��t�"�,�>�j�5���A�����n��Zں7o�eK)�d��;�)YQQv��{�����;Ｙe,�駟<x�Nj�)t�����Fv�3�E۲�	�Z�V�,�:�b���a��-%g��������_��~�OS��o�|d(�D7�I5AbܚU�#K%���@p��+^��%ơ�x/m�����ܶͳ�G��tb����o*�yBb�1�w��W������[��ڨ�hHW�-F2mhi�c�Hь9���Q <Vd�"7
gN���5k���:������YB|����1SJ9�a͉�Ѕ�Έ��t����"Lt@�LR��j}�=V89H�=V�Ʉfdh�-��̣�JjrECOvkJ�}��2���Gi�R��ėL�ؚ�?r�����q[��媳f����$�IXQ��ە�x�2�,=�v�;Nw�}�3��w��ֲP����������ʪ�}�S��Ј8PCSa��b�k�&����D�Ν�*��������K�gCL�����n�VР��	�~m����������\���d��[��bK�e�kԕK]@�=C�5��i@�mא����ʉ}d����:����4�ı�4�`�e����n)��o�/L���@!�B���ж�!R�����ߟ+�
R������d<q�������.���9����ۡ�v�Xb�,g����ٻ|��In�pK��)��w�����gY��,3��)�E��ʊj�n���/ejFW �ݽd��7�[��Y��w�.��"b�Y����ꅧ���z��sK��/�2IƆ�'�Zx�Ϳ�P3y�ߠ���]�ۇ�}�@�WCd���.U�VA�,�fw�����Ϟ\�n�}ԁ�@��x�\ݜ}��۝-D�ɬ���a@���5�
fb���` ��18p�7'�C���qN��.J�a��;>9��]U��]^�-�ir����bk10D�c�&��I�k���bn����45���P���7�km� �_׵��}�H`KUUe7�6�՝D(O�l;L�S�~�Μ&"������6Ϟ=oWW��ԩS�?���;��&���ģ�Yt�����d`)C/�-ٍi�┑%$���A�]8�k7�)8tXάͯ�#C�.g`��si&����f�%m��X89\<��)���Q{ �ؖ5gL�x��c+�l��IT�����.�*))��f���W_}���|�;�cx�x��I�;N�N�<I�1Bc'��Ѷ �r�,5�@�}��
���j���O�~�*|X�WrC'�~����6o޸����U�Dj��������e~�Ū��4��U��.�b�+W��N̞fT���̓�������_+0�%�����1O`0T[�j���~^1i�>m��?�)��1��X���/��B�p5��)�s��o۶m��q�Ɩ���������/u̎䂛��/܎<qg�6�sF��SAr�j8>���O@$�u4r����{���i#:C���u�=���cZ���v8J��KK˳�Q&C����x��zaǖ+�Ω�:�::��_BK�HO�^�]���~����	�J�
i�,,<��?;U^^:\PP��
�����ԩScc����ܴi�?��-8y�����Y��o?2-�O�6���bu�Drb:���s� I���K�bR��=[Z,�j�חC�����ɥ��)�|�?|���p�_���p�Zn(G��!?�Lϒ|���K�,3��{�#�d}�|�r89���������=W�v�-Z�h;��Cؾ}{`�[�����*��\3�a�M@y��v���,�}���k�����՛o���g?�9��𨹹9�s�ۓ���>|�N��f�	W�<�@:u:���/�YR\�c���/.�Ն�W�?*>��i��n�����ߟٵ�����[��)��DO"�S}ٔ�Ӯ��巍;�i3?B4٤�`LdD�t[�ka�)��%B�(VS
�,H��ux���������`KK��Q�0� z�>��F�xst<����	\'3X���²UL���N��������3m˳<;O�k��Z���"?�l��Y?�D�u%'O�@���L��˩d<{���ʅ>�.څ7H��"a��8"p�Wo��f��9���.v�!�~���x]�_����������/�qGEEIXz�E�@�?��y^�'�F�����ٛt~���kcc�����v�,����Pۇ�D�"���"��k!]c?�f0B.!O_w���w_U4�hf��i#]�Ieʈ�TQ�R;\.���=�	�,6לZBْ�`��E�+�[�.�l��Q�}aU�v�3�Q����l+���}va����!�L�a��C��V�O�$�db���C\kM����Ρ�<����t�^����@MM�.z��gh՜9sz>��O�����O��ɽ�=��5^ӬJ�#��|p�=� %b8	(����tR�<s��>���sFn��ٻwo�C=4mǎmK��N�H7��QU���;-� ��T����M�,z}�ܹoN�;��	�~�������+/��ڻ�EiqK���0�J�AC�*���TӲe�,��w>zC�.��d�R^�L�e$3%��OYn�9�?p�رW~���u��}���۩�m�g�C�gg�,jd+
:^���N��<\ˊ$tPp�p�2N��fx�>��}���LR�� ���]V<��;M9w�+��[��x��x���	3v�?�����YIƒi�NXǆ���ck��v����gI�\�)Z/u�x+PR�5Z�q���vZ����;���z�N��v%q�����'x3���4�?�)������(]c�|����M��Em�Uɤ�M|�T� �Δ��5�y��)�.��Nj� �/@���h}7�5H��8�T|-�:��XC��� -ax<��6bA:mK��ҳ�E���c�#���>��ʕ-��A��%H�Z����m��Ǌ�(<;c��t�	��\r���{�ݶ����M"3I��S4Ax������ӷ����?m�b˖-E�o����+�-����=���3ˁpCq&f�"4�ˊ�'&	��N��f���gՊuN������.���.��
�R(������w�,))�p�mKV_s�U[�ꦴ�g��e�����"�r����(J��>��C��=q��e�Uu���C�6u�?�ʸ4�Hr�1�z�LӜQYn�&M���s��>۹jժ殮����g6u���
�gW<˵ɂ9b0�\3���R����6�e��9|���<�g��vC� �$��ښ|�r�+K��E�F����d�#Wi�+�:`��a�Z��V�2��{�14O�S}��κ|�V����A!�께�Dt� �2DH���oC����ണ��&�	���r���I�C�ieP��W'rci���ј�$�?�![/������+|�p:	��3�s"�tjD4�n�.l��-u����r�)��`���˶�f+�C��ӕuA�.��z|�&6|�|�;���9CDj�E��?�}��'`mc�o���p��`�z�?�;�*��b��
�t�e�e5p�� ����&Ԇ=�Ph��ŋ�ig9����<4G�6W����ǻ��rA"��1���Ô>~��ms��[�bŲm4�����_}�����+M��>�7���Q��Ti��?L�r�O�o����5�]���9d&=~|hn��hF��Ȏ�u�p^�<C�7n|��_ܿgϞ�#u��1��`�����aG~�v��1�EG��D�r�a�5��3�e��i�}<ֱ�D���%2<����V�ػ��F�U�u��*Y'�;��XW�Y�Y��Be˅7˞�|y�3]���r�3.�bjg{S>��1L';.o��ODX���]�ϲ�9$7_�˿�6__n3�g�[vXDl�_�l��D6�ߵ#����d����eK�|��X��|?�5���cՑbˋ��փ���"c7�/׃����P|L��gK��C�LX#���;���^��O���{��^�������_~�j��ퟤk�R(�l�h�-OR�ⅉ�%I.�K�+厹s箝:u�Y��0�:����.�4����&9r����t���)�8q�+V\�v�̙�i�٧��z0��Z�ᅫ�V�۷�nc_&J����ᷗ�rメ�״��̶N��_}��q��9�J�F�	��%K�Ĩ#���㏷�Z��epp�3�\�L���<6�43b�-[P�� gf��� �.�A_�  ��������{�<@�>��d��p���3������|7֜�V����X��� �"���
a󉏜љ	�5yY�c�Ȥ�Od��cI&G�3=�(�B���91y`R�V
���k��u"�=[T��9#�����󶉠;��\X���C��8��o+[sK��$��LT�<�R�%��sd��0Qg��G�HY�:�A7L�{������4����Ƥ����?~�{K{zzo�kU�.A����Hn�~�U:���{XH���Mz�a��W_}\;9��������������h���y�ʈ��̈́����������x��mS�L���b�;�N�wY��o��RM���H���M�[p뭿��_�&�
]��'8���$���&˽"BG�

 ���s��������?`�ƍ��A�N�ˠ�@�m2�3H沼f�N�3j,	�61@���kTY��4����u�ۊ������	��L&�9��}%!����F!?
�(��o���z�H^9��u���`,��̕�r�Cy0��Uօ��V�x>�}x��xy[Y�Y'o�8v�`Qg ��#��-;�#�F[��lȚKScڪ%"r� ��c����\��]QrI�`��.�Abb��x�.��v��
{��e]�l�a���r�;�1��4�>�v����/������ݚ6�s#=���;w��8��$:o�	�e��������Y�qM��.�����â��Ύ�(�XrZ=�%w.[�lc}}}�\��MnL+��p�M�D�'�;��)OL��g��N�7n�?�X���ȑc��.���k��fgcc���fh�5���->���@"y=ͳ|�(�q��>����Xv�O�9g$�]�ao_F�|�a�����"QEmtHS��.�g-L��իW�~�g�>q��]��,�Ψ�e�ߝ%,��ٺ<���ekk(xP��A��&��1Xr�u*V%g����<�r�re��it�b��_!��[^xv
0��-"9�Zd���{�q���-BUUﲼȃ5��Sv����Hu�\�6c��vfm��J��Q&����)[�d�G=�r-[��v����I&��b�ߖ� �.v�ʚ
��,������W����ʓ�U#�d&�؎�S֪9��'d***����tz����=��O}�ښo|�b�����E���?����S�X�=�m=�����\5��hK���L�"N�<im�\���D(T��̙3���c���&����@8|�<�1���f���^��
�>_oMո����7��TuL��`mCD"��fe~��e��G��%��^�?X(���VU�f�u��η`i�8�H&+S�?�1�GϸQ��HGJD&��Y((\`8�g���شi��-[�|����wR�^�'�pU�S�Y1GL�E#���#���@h�B3�\����`�A�6��ʝ!���v) ���L?�yQF�ёK9�,|ι�@�2#n&[Td�{�rc�+[d+��~&r�s=�b$�'#�'7��)g��U��o7>�|"%�+�G���K��ɵ�x��N����d�;�T���"�2���G#�a}�в����a��հ�`a"dGt�\Ulqcb*[��7H�U��q�Dj�i�'h�7h?�,Y�d������� "��<k��}QTX���}Op�����|6x�L���^ :>@�>��EM_�pἍ������"7l�!RS}������H,��Dj� ��EE��Ljx��؞������"|N-fK�o�S�M:�jpQJxIS3�#<nG�/Y�+�`a�v��;UT虾N}�0�4=Wn�Li�L,��$�\��(�",]�t���_y啶g�}��رcw��3\j��q�5�x�@ɳh�TȑK<X�bPt|\]�-C��@�É�0X���� &σ�<8����r�7�h�[U�s0���0˖�3�[��[�p�|����/n�Hr��y��)�ұ��[���e� o��ȯ�͟��'C2A�;���L���ͮ˟�����-�Vv��ņ]P|��P���>�O���Ä�	[k`)�s!��xar���p�j�[դ�Dxw7������:u����総��P��e��~�o]���m#G��%��H$�nj$�knnӦM�蚘Ԗ�&LxmΜ9g1���xOr�����L<y�h�7௏F���8�9�N.SR:\YU����j���A|Vu4��V���죷��s��ƛ�BO&�SG4w8�r�8m�_k��U��{cr�0FF��.�O��0�I�q�!�
��ǂ������k�����W_���$=ӓ���3�|�TLr�;���ؗ] ��?���5���'�![p�;lّ�y��i<`ʖ~/Zew��>��L<0���f1���'-��F&)��5"��L�@"9A�ܶ�*o���Ǔ�3�*�-x}�t��#N�{�1���$H������F�;�(�>���H;&��{9�M�`��E��b�^,qB���Y��-����uhk�>��i,���^.����I*i�H�?EǱ�ƻՕ���~���m����5kָ_}����z�""W���}�v(���a��5>z��E
aA�{�������k.���\im�"7 5İ�mmm��T⪮���鱨uyt���Ё�T*�UX\����<)Di�|���Z^�zt�'�;N�]�G��N%��nbXw��U�kg̙���i�O��)��wJ˸��J0��+m&�.Q�,7
�(�@�끅���?�e˖;��Y^TTT><<��:T ��e��<����NtbLj�sT��A����4G��`*ko�(>�����F��O���3�7'�������G��P�E�2!x/1�����\e�vV[x=#����!���t��<�m�5F��l���<��ێ-~6M�ЫȢ`��s٭���d{r=�G������\~%�MU�u?ّa.�te$�����d��+#m�@�"6�������u�����Ϻ�t4������������y����X7'��q�e�t�����~z�w,�äNfbdj>VYY�����{��y��d>�R�ǎ���fq*_lf��2���о���-����b�!
h�����{p�������Y�q]��}�]\�
��.�e�����?;��n�W+��0]��.�n3	Q;�E��.8V�z柾�E;^}���w���).�N��2���̃����$�.2�O�f�����Gg�Y6|����L�<K�-A�eu�)�]�y�/��� c��B�\�Mv�v��[s\ZrT��[�Ɉl9�k���q��E�d7��l��m8��-X����]�<#i�u�L���#�$��Ϥ5��>a��eZ��I�\�kb8�"B���.�f�y�C���>��}��e�,E8F�~B��d]:W������{�^�yΜ9{�򕯀�_���ň��חlڶ鮡������8��Юra[vIM�81���N���sKK��;*B�_s�5�m;w{��y�s`b8<89�L��uW-�����}��YZZ��%O�3��N�k^k*(*�����ɔ�,��d
�Ԍ�E��%o�Ob�����s���&�nP���L�V������((| �1���U�+��Y�i��[��[��\ր��'�ʊ�q,:0���䋑g��S�����9�������d�«3s�z���D%��Z� Tv�Ƀ�l!0�B6G�֑����'#,?.mĀ�_D�L���L&�6r�!ٝ�ߥ�\��l�a]����"ڻ���$�ɇ�Ȫ��D���s���_/Y�-�}�ߕ��yc,�ŏKj���b�ϱ�+�����2�qG��G�?���Bm�v)Zz阚��WTT<?mڴC_���,K�}��'.V�=���+z{��.���pm�bj]K�K$�I���I�+¾a�A�b;D�9mk�uܺp��'�-[x^R��O�l�'�`�����c��E/C}�&�.a�C-B)�;TZ?n�,�Pw���:�����|F�c�]�fw��E~������-He��+�t����H�

c ���Q�v^}���W׬���ڵ�\�E&PD�Lʶx=v"@+�͂ݚ= ,����Zz���2)��"YUx&����5���8Q6֠��G��P}�4!�������bM$aQ��[Rc��Ȋce�k2���V�u�L.�0��	�מ�r��\o	�a�����&ߵ�d���L��&���z�Bd�'郕Z.3�ׇ�r�9rdW"SY�#[i�y~��h��1+�m���A9Sl+MNG����.��I�|��Be���m��Zh�/ѽ�̹���ַ�A߸����Ŏ�omnضcǝ�hD�U�ˁ�x��5B%p��ul�����|��~��>KD<{�l�2�k�v{��}eɒ%��s9}&���Kz�[��E;
|G���na[2�ɟ�v�����t�@uM����xYݤV�߯T��=-��\�c�+�.-ԙ1�I]K�].��z��"i%�;O�f��͎r����EK��zc����9���ֶE�Lf��I��ј��5��hAa�m�%�������n�:Ea[!R�ܼI&<�l��08ꥰ�~���x$�ɑ�;3�R�������pe������[������=���!��+&|l�� !W����3�J������2��B���������l��Z�wr��k��β��� �� ��>�9��50�^.`)�����^9k6���Qy\������Aǐ����wh�����X�p�N"7aT�����-.�_���ч~�93����e��b}d�&�A�.e�g���e�������H�&Im���k�]5cƌ�6�w74L�:0T)�j�TwT������t�{���)	�B���u�v�U�
uu"���23)���߫�4����[$� km={]6lصvݺ����s�鮮��`��&o�x"�|~+↉k#�	{�dr�5��͉j���t�\��&>|��+G���f�#�,��0d���!��X��p;z"���9a�`9��]�3���$'�d0c���8̙-6 [vd�
'X�������!�~�QA�9��L(���e�\{�ޑI�lIa�U~�_[�p��?�6`��$�>�ּ��ӊ��1�E,Y�,k��RC��IP�w����7VVV��>}��o|���%�|�'}t��֓�Ȥӕ�ڰ�κ]#��d�������������aO���>��<o��N�&����Ŧ��{RG���t�\ZQ�ZTV�����E;�QZ�f3�v�?�r���h��{Қ�+�0��\}�����Z�f�;n,���5�X�ʲǃ���g�I�T���!5<h�ˑJ�`�g�l]����L89�	�J�œt�+�Dg��Q�c�����3�u˿��W֐���s�0X���]dwkkXD�v�9�[�d�5���ڿ��(��1yɷP���Z�k�9h���m��k9�w��2��-4qK\�$V���l)������Ӻ��~7�/o���n����?��χ1�~����ݵ�����;v����1�~t���#ϰ���F<��R���wQj�5W_}���γl��<� ����q���_�3�k+�*��K��:_~�M�����t$KM���J��>_=D�K��+\�hҴ�o1[~�r�5��{��]�w}r`phv"���	�=OhV��1�L=������UnV�k"�����F���̛�~�בg���N��ͦ�灟I���)@�Z�.2�/62�w}' �; K�s�]]��0W?+W��������$g鱉S:[ނ�.��Ax��㒬T�^vw1�6/[kda4޳���ܑ�9���5�n�������m�HĲ�O��Ḙ��w�M����c���h�mDz_���ۻdɒ���v[^���[\�صkWɋ/�tG"��>ed�.����\��]�y���h�����}�B��޻'O����˗��:���܀Mvv���v��oS���jk�VTU���]?����j�;�6�����̚��%e�����hP((\DhҚ@rNn3͎yo��y��o/8v���'���fhx����B?
V�i�\g 7�ylF�g ��v�:Wy%G�v�)�:�b����?W�0s�yd�#[N�+��-�~>������u�<�#��������/�p��.�*#[�d���ؖ�3���������d�d������t����5U �f���:�������d�C�1�9A�q���Vmm�Ɖ'����gΜyA�G�m<��o�vM{��Ϲ��*�H�	j޺g���l�>���<ɠ�����ʕ+�j �zT�hl��;Ʒ���m2��)TVv����w_�FME�(D]ݍ�tL{��#v�)*f��'�(

!�.�VzVOoٲe�m�^i>�ε�m��M����9}NTO�f���-cds�p�A|dN�0�39W��9��`�À�� rX���p�<,T�Ů���V�Z��9J"2)ʞ�q�B�m�I.��C�����]�4g����2L��D��KR��.3�\�)d�䂔����ĆCѱ.��g�[W��Y#�km��mMbD��,�t��c�p��8���v� ����n�3���3
�9��G�^�a���ij�E�<L@-m��m��rۼ+���v2A��$�����@���7��\Q���g���|�Hen�(�h����y P�25ܨ�kR8��Eon��y'��h@��.r83�6zn;����֖;ٷ{��mm�W����4��:;��-9KD.��\z�-��`Ɲ'���S�c��I��7� p^+�JOO6�Gvkq�s�j˄G�~ r���.���|��MnF
��m����E��Q����N���D/�.&>r�q@��m������Rp3ɖ-v	�Ƞ9򫦦&�bw;���ȑRL��kϮ����zo���1'��>z=B��}�ĉ'M����+��?~L��	�ٳ�r�k�ZImh��о���rP�w���W���H+�	���>�����ܹs�\(O˨"7���u����j��<*n������E��fb�(.�14�~`��ӝ7���~�PP��t`���8�s蝃>�k׮�\���l|����i� ��3k�G��r�=���(���@�3�N�57l�;e��$�>�B���ph6k_X�*�8���ï�@���ɍ��[�΄kz�왏����욓�a@�`�%[��U&z�o;�%s{c� �U��l9�k�, F���p4�6�{c?�a1[|�b�XG.� G[���$�������)//�Z__�qѢEG�uX���DG���G�mmm���Wa���κ�kJ�g�?IG(�ף�v��{
���n��K�Ƹ?B�P����D*7��˅:�QCn�atDE�<���T2�<TR�YS3��M�&"� �8SG98�Gӆ��>��K�����l�X[[�+{�{��[�����6������#���C���2�#}��	��҉�#yg���ʷi��K ��\%�Lz�]6Lv��Y��Y�kH��2����2�Q^��kw�9�[.�)�&rR=YC��H#&Ol���|ȸmpn /8'~���a=v�9����XL�W���ꒅ�r۲+�-M��Ei��}��Զ�'�#"�άY�:�N����ф��7��ܳ�.j�&j+]ֲ��kf�+���Q���<y�*�p��	k\ST�v
��.����/�\��Fb�
r���GO�?��V�JC;'O�����Wǂ�FFA�����?���S��O((\���|�?u�78p�|ǎ�>|��g�`]'�QI��7�1i��59��=�9B�����Zx�PpΣ#kJ�u�d1�Zs��,���#�k#C�}�\i�u��r;� ga�E� �2���+^�H7�<���!�L:d�M~�XJ�6 HvO��4+�w	���2�}AZ�f��l=b���%�%�'�_�$�]���hG;dܗ=&���~.�}7d�v��s���&L�:}��=�g�$B3��N�7o�~�W����p�:��
L�����bK��91�g��d���^�d%�����g�V��N�7���k7k�\�'7pE���=~䝯P�^,�466�gAAɺ�Fl +!�[?F{��RPVrD"��}���ٺu��������*�"�O�N��?":�	��6�h�|1�&R�Z9C1��$�i ]�GF&%�k�Lb`@��ȳ_��@��Wdf��,A�&t,9LJإ���u?h.���
R�o-b�����[ܞ��-3<�I9bF��aKg��povgqrR=&F.�6v�9m��ߋ�w��]���{���illl�?~7��/� :�������~v�#Gory<%fڰ�#H9�[ppmQ�kڴi���ò�! ���`�(���A�Ϙ1�{[.(��ņ��䞞��q��[<>O礆���yk,�n���ñD���+(H��|9����>~��Z^9|�`���������4р[C����EuiK��hL1h� n�z.�[�
Οɢ[y��g��6�|�)�Iޖ��QF@>�y/ѱid]-#,5���a��bf޷���=�	��ɉ�q�����=v'����uH�8,[�d�|l�K0I��g��p08:��t"n��1:�!�K[��뷌?~#�C��I'����J��訟��'�w���j�Ɉft�����aٲ���C�Yd�ݤ(���rȲܔ��f�84s��?е:9��#7h�ӧO�8u���.�~3��'N��EQQ��Jl���ܗHDƅca
��p8n+<�ǅ������k�@�<xU{{����x��FF1�� n1��h���X��L�d11o���i����9t��1��r�H��u��!�b#kJL#="����dR�,& ��($>/�I�&e�E�-�	gt��$�%D�xem�a�L~�"9i�_��;_�Ġϡ�0����k�ޟ��O1;:nܸ��f��K�$�TWWG���X�zu�Ʒ�ߛ�Ǘ~���UVAҥ�8\�3fX�p��Wp��j�kd騘��+���\s͛�%��������*��}٭��A��he����ޤF��u����ܓI��D�PPP��p�*�����|���u�L������5k�o`V2���>��4ܦ�Ӓ�+ ���O��]�@w�d����kn�Ƀ �m,ב�ǆ���Y��.jd	�P�� �Y�qs�)��>��<xq�m���J�����ے��li�&�F�n&��d���A��tޣ�PhCC�>���r���6\YY�T.���m۶��_�00�������X4-�����n $d�$����BX��E���ŋ�Z�h�y+���pA�M[[[iOOח���ʒ��}�5U�.-�x�b��� ڷo���jH��z�n̴3�8|�/���NK��C-3�;�g��������D"D�\�V�9�j���$w w�2��z�wYv ٵ�/8�39�9ߪ![Lx[& ����n���a��̎��'��� ��ٙ=������e�|����|Q����n||� 8�\"�p3�xE-'�,�뮡��`{QQ���ښ����{fΜ�5y���4�B��QQNg����>��sK�?�%�^���s���vU�$>|���Od����=;*Nd�^;>~��ǉ�M�３j����cI3�ϕ����P��@�x�fW!�(��ܕ�FA�#@z�`���w�ɷv��<q�DQWW�����Y���S�i`�D����._4�p�.�|u{�AWآd�rgy�A����8�����}�Շ�����������xg�H@k��&�%������AEv�q�?�����Z��	����ed��֕�^��&Xe2�����ޟ��(?J��!"0-��2t���Ƹ�`L $�������7���/�Ѕ�A��}�6ҖU�]�~�׉�CT��D�:s��iZ{�`IL[��Mz�����ᦛnz�B�9�+�A⠎���d⦲��S������͎���(((�;8�],H��A������e%�zZ��i���S��p=�0kh�Rꀽ�x�J�n~S4({�i��B�+ ��Ϸp �Ȍ��=�E���X����ي�D#?Kr�o8픝���Iv����]��,�f�?r�?�v�+1���@  7S{UU����ң���?E��'N�WWW�4�j:�X��3%��}��T�Z��A�Rae�u/�D*���@r��Z�P�<�cǎY�m R����n�C���d"I�Ė<�hѢ~1�p�-7��Tf\yE�����������QPP�s��X�4֢s=L�~��!{{{�6KN�:��뻌�o���H�d�K�S.����0< <v�a�4���roy�d�6aq�ɸr��R��E�����ɍL�dKo�<犃�q��"�d�G�䰐7_ă�W0�a��.˵��e@d"�ް��t��]�E��Dĥ����dEEE/�?XRR2<c���%�0ؼys��~���h=y�3D:����v�J�'�1=>o�]�{�����s�l�
z�������� b�B��"��+��y%7԰Qj��J�o`46������U�n�!�n�������ttt�J�=ZC�g|��D"5.�LT���D"Y�ɤ�il/��?@���e3$9����KX�i�L<X��ODdݍ���31�*�2�ב&3�؏-H�@YQw�T��k	���4��x=}��w�w�n���u�B�'�k�O��ֶ���;y��az�766�T>z /�<��ĉ����za��H;+�xX�p_�]��H���Y���JB�r�S:�����Ǯ��׮�����L8�䦦�&B�
�SPP8op�aA'�G}�qzu�>}�}��O8.���,������bhh�&�USGϯe�T��02�4@x=ܺ���]��!�<����#�`59�^��$<��ɢ�� �	�u1�.�Ö�l����aA���=LJӵ$@�=�}�N��🢁�^�%%����q�K���啃�'׆i L�7β�)23z��/N9x����z^N����r ᢕp�qM"J
�a���\P��Ֆ���O =��c�i	P�{˼y�^Z�|���8�bEl.$��,,��~�M�E���۷�Dp|��i0�������Zʨ�/�����b"<��d�"�N����P��M���.�M�a-D�<�A_�$�M������D���~�rƸi�l�(ٟ���ٖ*"2����N��bE���5-�r��t*�v�<I��`������@o�0�QPP��y{KK˺}>�@EEh���x���,^^^�1c��.2D���`�{��{����qC2�,b�X�E�X4�������rU!�4t9����D�{���\�ti�h&��������3x� ή�I8i�Л���D\���.�ٺ�q�'���D"OO�0D��@*+@("C�t:H��T*W��02����dO&�v�������NjXs4�@O0��z�谶X�䊡�%\.w������DVb��'A��Xiii�f�P(4L�'��`�L��!C�SY`."�_�>��g>�D��
�q	d��^��5UUU����a��Q����[��%
�Nxx/�GO�q�oM�4iTG�)r�������������,�����͎����O���АN��,N$b��h.WBK&]DjZ*��<��E��o��":~��N.W(S^�����dL��DX��t��llL�xQ��K ۶m�����_��y�����#\N�,�"�`�`�A%��ޞl>DB�İ��+N����=��E���={v��P�FAAA�,@�R�P ���~0�؉#�J��#�'~䄏x���,�=gن�ٗ�>\X�S:#988�c�ܹ����{���@�EEn�(����o;����'�&R����)�?G�q�,N��8*46����k��i����ꏷ�v��E��1�={�_��[{{{n�z�!�H㢫���l�Ć0-�L,a��@�7¾!���\��I"��F/�X�b��i����"7





c����~�����_�x=u�%�#�F -��pAU�$�H������bRÕ�i�m���ٳ��;N�%�"7





cȭ���tƮ����x��!�6�g@Z@d����X���p"���ʬu����p<f�������o�y?m�c��((((((�1<����[�n�"�����dJ�pk�½\�].��ua���:��p2Xhh�NZ���;^�a�g�"7





co��V�C=�W���'|>�Kj~�(*����WXft������K���L@��̙���ŋO�1En�P7���V�v���!̚d"�YD�!2��a��h)|�e:��p�7 ��a)ZOSSӣ��sϑ���Q��1�7�xi���{���zg(��a�0��	O&���P���OI". -��ư"�@f�va!��)G{c�����Տ�q��ƚ�F�"7





��g���/׼�j՗�.�R���ȈBx=^���*�
�D$����w���uP�V��u\.W/��ԕW^�jڴiCbC��Q����k�\���{cUUUq�4�H,!�^;Q"�`�QAo�����»���Xp8*
���-r�u�@���Z"6��r�-�b�C��Q
Xl}���o~�����_!R��u$��I~���a���`������>y�:���%��֍J��<}����c%��A��Q�5k������_v���O�>�L%'t2��]*��&0a���3s��={�d���a��rcD"�V"E�q��kkk��"�"7





�O<�D�?���=}ݟ�����W�q�*�L����g�k��	�k�2�H��ӧ�}�zd��\�U�vE��m���bŊ����EEnF�~��гO=��hl�ۺ�O7twA�4�h"n寱�P	�=�S\b�������EEE���5�@h ,�z��!J�ٺx��Go����"�"7





��7o.�կ~u[Oo�W3�
".^X\�rJ��H'Xj\n�0������E/a�@pt�ml����.��I�'s��{t�ʕ�N����((((((�@<���`NG[�=��5���#�@b4���5���	�e'��	�0�������-2������`l�ݮ>���+V�XS__�QPPPPP�� �y��'����7�f�GA���5�`�IeҖ{�#��z��)**�փK
�X�)�	bӟH$��0��~���>�QPPPPP�� �ٵk�ķ6���Cᾕ�`aa*�Ҹ�Ծ����}��H$bYt ,������ME��h4:L�����_�r�-�D|2�"�"7





%/�~����֏���r"�G��0������;V���	����(&g)�u�D��{<�_M�:u߂�ly�?En.���^Z�zž�{�%R�H�ą�
 3YR�kB#��u��������\ ����RLx���js*
=6ujӦ/}�K-��QPPPPP�  �oݰa��V�CĦ���-6V��S�[":��ȋ���+�cbN5p��̘1k�����q1C������E[6o��dk�B"4�d,mM���h.���LX,�#lw���'p�b ��*(��9�N&�����cW�"�"7





�DT��>��oo��9��W=8<�!�����~�0�/\Pl���4Z��Ȗ���+��S��'�1L��'6�"7





���ڰaì�_z�s�Tf��pDKeL����zuy,댮�6�9"c��f=��gC���F����x<.�H�,Q1��&d$�(���ȍ������yD{{{���^�\wo�b"A�V 1aR��D*�˺���"c3�Ñ�����7�� �M�6��F���" %�����:x��m�T��H����0)�*�E��b���3��E�2!rB��������aq	@��� ���n�:sㆍw���z���/�!&+dK�"~��˖lK�Ơu;��ݴJ\\P�FAAAAA�<������_�|__��D"�O�Ӗx:��3X@L�.�EN�-6��(ƙ�-�ﭩ��}gŊiq	@��s"!x��ۏ9r���PV�,�aXv#��A�97�L��;�	��~���G������>q�@��s"!�u��-X��ͻ��ĸh4�ЗC��n&. 4���-7L��j#�_ d�Xm]��p������?}IDJ��((((((�C���5����w������� 6�A�!R�و�t�ܰHمe�L�[J�� 2Ir��%��[�P�����K�j(r������p�@$��/~q��#G?�C�Ġ��$����E0�Y���iY+��3X���ٵ�1�'C럠��8q��K�j(r������p w�o�1w���(�I��͚��Xa�.��n+2��95��������7jkk��{ｗD��En�2 >�rrº5k�i=qbF*�@&��hX�vbr#縱H�Cft�`GU���߁4�I�:[�n���������_\jP�FAAAAA�l#���O<x�z"Ű����(�|��l�9S$�����b�WX�`������F�?;o޼��B6�3A����5o�={Æ��E"�q�l������[���n&3�*c��G����a]'I�\<�L&�L�<��{�'|���K��((((((�%�u�����=�%R�CdG0qaK@�K�E/���r爎��������`*�H4���G>����^�V@��������7�|������E��1�d2)8��c]yW�>�a0�a��{e#xƤ��}>��.ܹ`������ȍ������Y ����뗼�f�'��xE*�ғNeo,�XL�Q*���a���Trd�lx= �b�yJ�~ޮ��x������ .e(r�������wԩS�._��ٯ�S�9�n�����t�!���^Z�}f�Chi�����ә�M\�a�lW����墨


�d2�����nѢE{/ewC���$�{��>��~r1?�g�G�+�LĂr���P����#"���bdd w���Wf͚���oN
En>
Ps�ߺ��L$�D6t���D:��ڸ�i������#�Ɍ�h�%v�[����p�DX�F����丱�D��VVV>��/�[Yml(r�������g�ȋ��ĉů���_���N1͌ni���,�b�n��B�9�$y�B�G$�c�v�����z�R���{⪫�:@�B��"7





&b}�qO=����ۯ R��"�H�Dd(.R3�`V��#4��!�шp{=�5�䴡�l=�aZ�5�%L��t�6��6Dn"�t�5䴹��B!En��(��5k�ؼqݭ}���X<��R	��W�rgú�J#�EQQ	�V��D*��q��/+��>f6jJΉ�Xn��P0|�;�8��Q#�ȍ������b�ڶm�C=���=]��XD�x\bʔI���N����â��Ktt����bh�_D�B�xEQq�pytKc��nYj�(��F�l�>��x<>��q���.\����)!F@���}���Ly�ч������S�Lq����X,"&M�(fϞ-�~����X��CQq��I��q��Q�7q��{�N�Io�DMq�����w���+**^�뮻"B�]P�FAAAAA������?޺}��7������F�~�[��f��IDF��/E���r�xDaQPL��$���DS��v�S�صS���"
���"�J�Y�uM�TJ���Τ��!֣[E1�ؤ��_XX��m��vL���En>�=Z�v͛7����ؠ�]��H���L+�����tҎnvHx<����4{�,�l�2q�5K��O�A4�kS� !��aa�:�~%Rc�>={��3g�T9m���((((((|@ �{ÆMW\q�䫮Z�۾}�hk?)��b�����ȍa���-�zQ����03+GMaA���,��α�ϯ��7���KTU�XI�	�̸]����V��'Ni[c�Uw�uW�PxO(r�������100P�N'�]�re]ˁ����7���*��8�"6^�wk�En��I$"O�t��}VR\,��).*�dB\�l�hok?�����U�Spe�����ܢ��oo���w��d��{B�� XmR�TS \����]��QVV*.���rE�*\T\ ���@C�1��@|��C���R���@O�H$�b��bɕ���u�ĐwP��VX"b��a�i3,��~v��y�;�OC�������X,r�if�m޼�
�l�墶����X�""��5�@l�ߦ��<�4TBd(dE<Ň�,-MoO�(Œ%KġC-��o@������O䆾K$�h4�qҤ�g���/�|�K_
�En�L���}+O������͡C��ɓ'���"�}��KcmL4�d��UO*� �cj�^PTVV���r�s{,b���D�֏��`��5c�x��5 Q�8Tf���4>�p�fUb�A����ڄ������ϴ���k�vwA�/j�W��	�E2>�W��(�i8ل�"��{�HJ�(/�e�x]n����^+�q,���jV���D ��T\K̴���{��fΜ��+�B�A���Ga$2pSO��%{w�ģa1c�TQQ^"�a+�A���v[.(!4K�L	��@�W���Z*
�����>�HFD$�DL$3)QTR"*�j��I��;ﴈ`Q1��)�k�++˟��{��^����ȍ������{�4M___ג���/�ٹc��֣���QW?N�<�p�Maj.+BJ�M�E��E&�E�E�4T!��Bڛ.�ɤH$���>*�>�O��.K��g�~$�3LMk�z\��7o�v��pP�FAAAAA�=04�3����G��y��!:���z+����j�^�Gd��0M�.�"0�)


-��[�2	184d%���H$j��z�R�}��q3cd&V755m���Utԇ�"7





g�i��������h�qǎ��{w�#�]����ֽ����f����ǳ0���DD"��M$@(/	R���׼�,)�%a�	2$A(�3�ͳO�L��6�]]�v��ί�G(o{<U���KwOWU?���;�s�j�B��34>>F�Dr@����O�w四�9��M���2�p�1ߚj�`�ju8����7���dP2���LӴR�4�a���(}�k_��&V,��!�   ����U������W�_�|�����LM��dY�Z�x����@������(�0���y_��� �p��t:��P���&Wl��:َ'W��}MS/ۖ��G������  �o��Q�~��vm��k׮}��=��������0��y�STl��x���d�qT�T�/����_��|�^!�r�e2��,9'&Z[[[��'�O���^�q�o	�  �7T*��5?s����ܸq�	_��y��<y}��j[�)��X�о(���.g��e�����uz=����z8��>�q(x�_�V������OO~�C�}�����_'�� �   ��������n��ŋ�����ѥE��?D��b��Η$�\���{l�b�GL��D��8�"��n(7��_�~O�uɴ3��Å�\6�\�{�g���7^~��n�8�w�p  @��^�:ӨV�p���W.]2����I2E�I)��1cp%2��r�E��_���qWm����R\�	��#Ӱe ⾛��j��{e�ַ^xᅛ�>�lD�;A�  �oԶ���Ξ;�z�K��89�MI���r���*��*8�*�'��yY��{=j6[*6��܆�����V�x_q?��������|�ÿ�?�=��O�;C� ����4��T�;/�={f�R�(�?y\Vm8��?��-�����Q����<o���\� �/�l��"�p�MW���-*�uȰ3$B�������lE���م7�����p  ��~�qpkg�s����v�277K���"��){mTyŸo������'dՆ�3�c�3m�(��w�Á��8dێ��$Z�t���|���sSSS6� �  x��@�_�{��7�;w�t��e��6\�15CGɣ(E��N|훛�y�0_��D�X�۾�-��:}p�uj�o��0�ER�t�����?����n  �%��Y��~����s��M7�M����O�ڃ`��^�&��R��r��w�0FI��@�'
y4��V��u��EAG��T�85??_%x�!�  �c�oG5�C+k��_�z��{+��9V&D�1��ĶR����~s0�*�����0���7�W>��`c;���-�?
Tո���`��+���  xL5
�F�Oj՝?z���._󞟟#��ɶuR)�����{m������нl6O��MM�P��Q�ӥZ��`�_�#(S���풪[�3�8U��i�]�PxC�W��%7  ����Q��}�^�~����鴛�SO}�,S%�TD��I�J�@�y;*�)��:w�r�"MO$7�Q"�N��&�d�GV\�	�W��xy�y��b���:)��f�srr�K�A� ��
GU�թv������}릱�0O�BVVj���j$oG1^�������(�.\ȗ�X'M��ލ(�����c^���`��/>�u7�~qqq���]7  �Xi6��f���{�w?s�����gg��f��l
z]rL�e�z>��M�Q"��y!&ߎ�-����<���(8���h�!�+7rD��(�""��+�rU���]�p  �>����������gμ9ǡ�ԇ��l�Adp��0hE�����J�t���˲φoG�A�`��n$��9�)���o��Q��5�G�B����{n  �Q�o���/^�|���7���8J��+����R(����5\�ID��.�K�r)&���AOC�[RQH�>�:�iP�� N�_d=�G���<7  �X����Zm�Oo޼�Ǘ.�ϗƋ49U&�[���ǐ��
��	��\r�Wnl+CA�O���b��;����NV��8R��a�ߌc����  y�a}O��[y���xn�ґ'DhQ��(M��12�p�aX�ʷ�H7-*�'�q��e)�"���;�jS��˹7�x���E��I�����}ϰ��ǎ�q�C�p  #oggm��[��ʝ�O����/���,�$��)�7\�)
�n�FE��95�2�+Ɂ~�z��@���ߤ�#(F�.���]��?l��ɑ#�Z�  ��4��]�t��۷n|���7����b̬g��Dr��(Je�L���}�nO�&O�������nˊ7�o���<�r9ٟ�$I����{i��M���  FV�����[O�[�Ϟ=3��r��4��M���ˊ�t�K���H�����l�^�X��t��^��Z���>Ǖ7�TUO)U��0�A�4}NQ���C� ��$B�����X�W��曯������DyL�c<y8�&�FU�5� �)?s5��lxw[�z]j�[��^r8��lx
q�$����8J_�m������{�  FS�S�ک|quu��\�d�L�.(^���E��n�^Rē&�q������)9�O�h����+6}l|9�/����c����a��UM��ɓO�c
�{�  F���ꝏTv+�=s����!33Sr���$��������{�"���"�X|U�?@ף4�d�M��"��Q���y9>��3���4I_�8�m��-�  )�;�R�X�V��z��['*��v�*��j��},+3�<�Ӈy_T&2�p���r���0�{�9ӦߑUn(��]T*?|����W='����l��=�p  #��Mowwfgg�K�o�|r�����4�r�<�ҹ�8�H��8��q"�`�^.[���*�'����
ro�9�2�%oX�܄LjE�E˰�{�x���� �  %��^�����ϝ�x:�dz�W&���R�$d��¡F�(I)I�I!]3�P(Ry�$���0�.7�P��Q����v���oWi���)��������yE9��Q� �  	|;����g��.�?�DmwGY:<O�lFĐ��XcȞ��X&5�M�F��T��Qs���ˎQ"����n��]��)�"2-W<�x�!�P��@m�^��?>z�h����p  C������T�Z�ʭ�k��|�^���R�Hn&#+5�C�O��(*M#L���}ʘ.yټ\����H)(����hP�ݡn�=��*rw��ɑa��$-���e�E���8�zt �  �(pv:�Oܽ{�gμ��O�r�\��V/4�r�M"�n�E��b�uól����O�>�E�i��ko�����'+��������l6{~nn��!7  0�DP���V?����/^��Vw��~��MC�,̕n"��?Fq"'
��\./������H^��a}�=6l�s�j�S���#R-��W
��)lj��  j���|�Z�ڵ�￷zG������tE�G�̲�#>n�Ex	�P^�Nb���MLL�kߪaP/��Q�8�p�ɸ�:YY�	�$�(=c橅���G�  �4��޾������?y��y�TW/�Q���y���Ã�zj� ���2�#�l&�Sd9��e0X�����&����"�����q�i��r��["8E��  J"xdVW�������ŋf�Qxqqq���8̏�*�$��x�7��%��M�8|�;�v�M�N��"شE����Lۢ���׋@�Y��i�)/��G�  �U��i�j/޼y����*�<q�,��&"n(�d����f0����}P��\����~Wγ�	�~0��0d[ٶ3��D	UM�`�Ω���
�#�  �N��o6[�{�׿�ԝ;w�'����x��)�X�Pu2[�MH��}��o�ˢ��irrR.Ŕ�Qr)f�|ߗ2#�ic۔�
)��a(���5J�Sf�<��G�  �4M�۷/�s_��pb�Ȣ2??O�f�P(P��hcc�՚��0M�HQz�T�����&�A�W,��n�)}�J�ee�Ë1� m���J13����\����p  C��on��o�l�����h��m�*
y�K�ؘ%�{WEp�I��Wq�q��͑�q9�P��2���A���� ˴�g�F��T�$z�5�SsG��0��чp  C��:�O�q��e�f�O�1����Q�ѐ���x���x���
�.���ǆoG"�Dl:Mj��z�ˡ~1��E����&M�DX�U�;�i����� �  n"��^_h�{�VUuB�����E�O�v����)CV���l,��*�&D��Q�rx���5�FS���p����QT�?�����}nn�E0n  `X(��_���ǣ8��W!tZm���V�*��M'>fj�[�yYf�s�L+C�l^��wz����j�j5�)�bl궼��q�8���Κ�sjvvv�`h �  ��0{���(�ƣ8P�B�af�7�
Lw0�O7mY���ܤn�O�G���+�P��ypt���`c�yn�L��$U�4����4�N+܍C�  �B�V���;����?s��[�+��t�}Vxp���Ŀ�2�DQBq�R�Z�;w�P��h|�H���đ�Ǖ�te�Q53�w�u�2,�ο--��vԐA� ���I�p�Q8̤a,Y�c�A�C���+ݝ�\��;.�8&M�hss��/:-,��N�J�N��ǐ�dȰ�tn"�L3sAS�S����7�n  `(
~���� � �D����&�8�lV^��pp	Cn���a>��Uח��nj����q��qrܴ�&��"��������<E0tn  `HL�M}k%����i�$D�L��2�.�i�lnp[�9�8�GSr���f�M!'5�1sق\��I�����k����T*u��  ��+d���J3"��"����*�j*C
Zrr���9�p�f�V�n��u\��dl�(���y��KKKwQ�^7  0x2p�Ѹ���+����%�lH�����$��T��vF�4��}GVp��]��=�.7'���(���B�,vG7�  �\���y���x���D�Ħ.e뤩�P��p÷�xj1We���_�g~8���*]3Tn�Ԇ���eL﵉��6�PC� �������_Lf����:��F'�41�C�J�-|���
ٖ#�WpT%�$�����0��GӌP������`qѿG0�n  `�LMMuvvv~�h�)�����i�8ģ���d��7Wh8�p%��L�҃�U2�Wx"EU������T�C�7n  `���V�V����˝�Ս?���㤨�8���LۑGO"����QUK��CWs<�M�0Z�����E�33�z#�  �R�X��i�^�������nﳶm/��isӰ�^�R{0��麞����v�iY��������%7  0�E�E�9S(�o//_�e���|��O� s0
����&�W5UK�$I�8��tC��d�:N��'�|rW���C�  ��^0��*έ[�.m�n<t��D�yJ�IJ'%%QU�oA�X���m�o��{�رc-���p  #aos��9�ׯ_���������iZ"�=�<���neii)Đ�хp  #eo _k���   ��   )7   0Rn   `� �   �HA�  ���p   #�   F
�   ��   )�z��gApˈ    IEND�B`�PK
     �8�Z��X��&  �&  /   images/9c69fbd4-c376-47ca-8b4c-793dd402431a.png�PNG

   IHDR   d   M   PA��   	pHYs  �  ��+  &�IDATx��|XTW���^�`�4i6P1�]�gEQ� `CEcԈ�%�h�c��(�h�%�XЀ
�� �O��_���o�/��D�,��a�9e�k��]{�3L������������������������������� �.]��Ap�HTTV�B^�,+ 	ll@ ��zw�'9��e��дiS��� �._��7BXx8dfeBYy9h5�&9�Z=�Tj(,z	�%��]��	\�\���������a���'���+�.à�C �o�h4�'�����K��3��)��sK*(TJ���o���[���c$F���Σ7d���|^GG��Ԅ�Q������Zpx�BC�Ӫ�lV���gs8O��v3f%���Kw���79x��΄A�!�c;�l����Jii���tHIY����
/�
F���b1�!'I��}Z�-f���d2�h�z=M&0�f�X(������i@cЁ�d ��6�U��������«_-�� �Wܿ���� '&Bt��ԩ�{��
2�֬�Z�/^��_�11�lllz���+���*���xR�4J�Z��h��C��7�1��j�#�3�j��jBPh#��l19�z��dq�X�<�l6K��rZ�16U��a7�\�A>�wrϞ=�.�ΐ~�,Y��K�!��6�^��� d�w����P�A(+-���Ҧ�X�TF��SUU՞Fc���ժTz�!����kg'y�,u.ܵ{K%bnР�;8�� `1[0�=
[�[ûrᖛR�����d��`��Kp��	��Xt[:@��h
���J����l�lw}��،�}c�((,���1N)���@�.�`����d,�Q@N�<	Ǐ��������!�mk?��iL��GC,&�QI���k���/��� 	�]�~%/0�9�x<x�<���cGF�u��;\,	�\�H�P��j���b���
8��;�Ɛ �\������E�����耹�l��g&p8�	���8;;]�������3�'KZ�n�eU���b�� 4$&&&��1�G 1�����ŀ�b�ê���dm���kjQa���,4��a�m.s؜=���O�K���3HcC�
u�N����O=��d�0br��[c5��Ӏ���+�r�f@�¨����|c1���H'y�J9�'��&��d�ف.3�+cW5	���p��v�ؑ��^����`䨑0���вe�?56; �.\���" �ys�ة���{zx�,++�ǜa��o5W1���b�]����2��C/| m۵��e{��QVV����&�p����� 0���x;�V�3-`�' 9�V��@1[��<���: �����ނ�C�Y�3l�K#�W���#�ˉ
l"�z}���4��b�߶=5�e��P�E��%K`�ܹo=> Z��m;�C���;��;w��{>����I&��I�сN�{��������˗K��{������D�Ojj��a2)�J�F#��>�'��5��ht
�7�����(�0)fs�j:�!����	)�.a���I0�@�Q��oЛ	�%f��m0� *0J�z����u:'[[�q_lÆ>�	�/7.������?��_C�M�o$77�̙ФIc�? ���W�t� ��
J�Z���
�(�����xk��pi�ڙ�a,{�,/�(%�B��2+�ǧ���bfQQ���)@��`0�7�Dj���d��֢�O��=�$#�����+����$j��	:B'L��KKt���#(Z�h��\giUu�Vo�uC����ӛ��f!U�,��1���$uJ(*.�6q�ҥ'z����?�^|�������~m�t��n
;�A梜�G3p ��C���	�W��
�6�~b�7<�]�]�r%U��z���k�L&��X/�cKhJ��#�Ӑ�x8ЦL���{����{���҈����$�	Z����p�@.S��S�c`K1JJ�{�߿��SǮMUJ�p�F'ٺ��j�ѸU*�L��ʚK;}�T_ԏ���H	 �Cr"	�%����n�����&mݸq�Q�`ڴ�o<^���7�,�FĎ 77g���nS(U]�x2��i������о`��|�>
�z{�<��Ѩu�ji]�Fw�&�,[BQ:��n0�
;��Ao�^�(3z K���W�ATT�����&c��Y|2y
���C��Ci���u�BQ;	��S[[��b5olָK��t�H$��_�߱c�o~���<|=�u�I�++�4k֔�*nE�N��'��/I3� ���?��Ȃ��aܸqp��Iprr	�v��~�Q��r��*�c3F&���9\,>z����^���;�JK�T��jͨ���X�
K�3�t!�O�D�S:�n	�ow?��D gϞ��BBB��у��G��~�׮]K�O�:F���q.��G��}�e�<���L&_#	������%.vv������>��dgg�iҤI1b)b	 D�?x�fT]K�Z���r���g�App02�����������/ �op��t��yx�f�8�V���)-�[�x� [�sf&��6G�0D�B?�![�*�J��ѧs�N����C��({@$U�Y��M���q�.hu2 �"-ZQ����Q���kp��� ���;v�dEG��q�ж%����ݐ:����R)+������sߢ��N�� FZ����'O�@�F�@�R�4���������~�����:�9 s�̡$_��p�;|\T��0V�b��b��铞��n����
����Bǎ����[Ԁ�^�Qi�4j�#ch�������L�����!������[7	s���̊+������G�M��|��_�p�XRR2��ӫH�ҬA1����͋x����Mh8��oyhH;?.���Q���0�_:�����*�7���v�v������w�^6t�o����x�W�ł��Q&`��T]UyĨ7ۡ��b�W-�>��.a��+`ذ�0v�Xx�"�74��L&��bѦӭH�>�������|pqv����W&��b!HQÞ=;��Llr�7�{���w�B�v��Ν�k��r�Z��H��j�Noo����rSX�^ u��|��igz�N���5���p�J�l�eeй3g6�(;[~������K�q���������p��q��������Ja!fg���B�hHUU��n�{��؉#�F��ԩ����k�W��O��K�+���ˣǏ-E��Ә����%���J	O�{��iй�2�t�
�������뜉�d����EF�a^۶Ap�����n�L^{��a��d�A���(�����]V^�]o4�����(a��ٿ~��g���:�;��ٳ��e#z�#���eA��`��DM�XZZv<j@<�~q�8�&���EPTR�c�7+/-�H�n�ް�E�@�ʊ�Ta��`g�8:&bz/ �66<X�f���k����0xp4����k�R�/��,.�w1#��Ŗ-������k��*�����O�؀I?Y�3��
�z��v�J�?s�Ӟ����\��#��U��['֡�Gv�� ¿R�tnFFƶ�#GB��\ؾ}���>}z��7�o4!f��`���|���f"�`���cϳg����x�Jm�5��^0��i��'��Ν�H�ì����Pac�7��Nƨm���]�Iſk������	�)�)�����d����>#��߹{g���I�r��6��_����7o.�H����v�Z��n2�Q9Iw�۷����Cee%lڴ	6o��������2���-�<��h*rv������d���k�@ �J�޹�)�ݻ;�޽���B�T�44���|�` �X�H���2����Y��4:��l0����ڿ�4��	2�R%��3�v���ŋ�O�|��)b��%@��[�24kڬwM�,�d�`�4p�$7Wg��k��>���[SSϞ>����d.�T���F�s'�P(�Z�p���C�V��B󟴘�
�NX�����T*U�>�;����'~����N�{q٬�LF2�I�e���Y�f�'�"M�Ģoz������,U�応�/r��ޠ8:J�sr�WP�a�*���N�>�"0))	�����d�������!��E���E� 4�@߉�`�b`�������l��Ũ�!22ҊJr5��HϾ</#����'�Ffޫ�ݥ����uJ.�I����VV�����iz��Ցr�<e�]�L��i@���
��ټyxz��GE�o���<x�y�.<Q�V�~�� {ezr��E|���F�V�&��z�����`	�!�͛S���Xy�8�{��\��#�v���z��d6�$���x�hJR��34pK�{�'���:)埄�����ز�.��)@��ǎ��ԛ7
)))N$����w�ܙB��l$�wF�@��@��.�(�ju¨c�EM�c^������B��,!a,�%w >>^��+t��s�-�ˑ�!��ҁIg��`��c0h�-Ŏ����NJ��/�In�V��s��M��
����I���%� r@�ύz���Zz7\0vl��&I�H@�F$ߐ�l��x����Z�ջ�TVV�mݺ�����Mt�Dܜ�fݐ��f�EȠ3H��+��^��d?��ju�޽���޳�@�T{�۷g�/�,���ր��4$�0>Ď��*/-#�I%i+�/��k�nm�hQ���`ggG�m�o�\���*MF�X�=V�d������M�8�J�8Х���he2��yl���|_��Ն�b�ϾĈ�^������qY�R��}�]�hA�+Ed���(o}|}�k�n���#*���?`�)S!;�*��ot��730��d�?:�o��GE�#7��P�ա�/i��ŋ��!����/���1tBΣǏ�}��|�l2?s��!g�%���Lf�i�P
_B6�CfWUU7C�*��㥷� �>$\�@eu�<H�@do/ٿf���G�b%-zc@�1:�1[�j��J�[�����b�QN�Q��

�'��>���8	fϞ	K�~�a�B����p�i��)��#�ސ88���]I_��h<I�������{,�%���t@@��B�6��E������-�d6���c��:�()ܼ��췺��/�ƍ����yϞOBY(|�$�j�#K�UU�cCBZ�_�p��˗/a֬$��z޷͜9�M''��4����j4EB;۹ s	V:�p�\��-~^~~�%Yb����R��̷���ܹu�� ����s&�2W����
.�^��͟�q��Ih����=*�*!~Tln�F�S17Msu�R�V�� ����`���g8n7m�S�M���bᣏ>�¶l�B�W������֛pFC�@(l�T4��O�Z�=~4 �ik+��=<<�?F@���Z�.5�>t��)dr���oȝ7`���`�(�����.Xb���q#���s�7��[�\�ƍ�����������k���|��BP*d���AQQ�	��~���5v�l}�|t�6�N���0iR"*,@��i�	�.��H2��ec�0(ʓX�̕H����ee%�6H[���@j��huݒ4�{u��o���k6�g7W�
a��~6(���b7-��wl�����o7��S7I�zI%^VV^���2���䤗�� ���� a�7�UT\tNlg?���`����cʔɰh��Z{�v��MHN^CM�c�����X`1�������H�A�X�`~�N3��~}H�������`Ϟؾ�8�>TWWp�W�@CZ��g��E�������U5�^��w�����v6�§D���S���
h��o�U۲e˨)�%K�����H����h��%�%�G��i����WVV�C0z�T^8p`T!Y.%`L�6��6m:��02?���oI��0 r�� 86|����BIIi6*B���[o{{{2�z�u%/��ς��c��ի$2�x?b�a2YYW���ܸq6nX�*��l|�"5U�.�D�C4�=8�02%FUÏx0�.�����nx֬Y������/ظq�ʮ]��X�#�]S#���R��B�|��v$�����qW�ZI����)..�C��Q-��F�ӧ�+z�kv��QH?zJ�J��<2�+�? r��`D�X68�:R$��K�"W羮�.đ�Fa����t�de�j���Ҝ�dR0bd<!��999�	��.�m۶�����`�h]4V�Q(\?B���l#��^Q��4f@מ��]��M�R!66RS7�3�^���()\VV��[;�[j0�!O@��op_z�Qp��9��q��X�m
�٘
M����:�7�m�&8v�(�J8q�{���lw�ڵ:���q�,):��b�y/1:J0�]xyz@UuU5�y�F�z��� #�3���v�ޝ���O��PH$�,"bX� B֎��1kV�9��.����d%0Yl�گi⧹7�h����='Y���Ԍ&���:v�H=1Ecܸؿ��v�ڗb1���dqU*%�J:1��+I�"�+�E7�e�?����{u��l��uf��,X�%��� �|�ͭ��6T�iE%�d)�<�PZZB}��G�B`���d� �T�Fs�\��B�X�!X*(,,����졢���3X��ܼu�.�#F����жS{8r��D���XD���_�n 0�$S%�/aE�*h�*2�e��l����{�m8��%yBs�	z;��:�z�]���4�X4x�M�َ��LX�|9�Ǐ$�f���4���v+��𫭭���M�NI5@��416����j4[v�qv��Bs�N6��.��t��5�s���H��VTb�j�&Qx���0f�H1�m?<f��}z!=u ���B=$�d��l��TR�o_�K������꧷n݆�c�)E�A�{�'�*U�$r>�XL��&L�`y�D�|��dd���*��͚�7i'�RRRfm�jm"O׫��yKV$��Y�@�32�i��Y�E���y�����S�����c�c�6j��1/��
 �p9R�B)�f�I�KV�0�(/%�(	|��V���x��h2�5�ڊ��J�2�^�~T��Gj3�s��r�NĞ.8�^������^�X����h4��E���uT���ԉ�1�Y��!����M@
� ��6�@`��m��OG'n@����l�f��^O�21���L����o���j��M���+W����qP�}/4��0,���[?�B�n��/f���*���j5?��`~~~�C餆,V�_�r%��	��-�Z|� An����
��Z���"��a� ��d9"@�L�1	j���Y���jukKֺG��ePF�)���'�`��α�ѣGW�c�5%r2�:�O�h���s+�J=��㢢�#�8�]nҤ)�5nu�0����1r�\�%'J�1F��54Z;Fw���9���U�˼\���QH3�\�=�O��o�y���t�^��>��B���)52�xL�����XPґx,y��yHG��L�L��B�"�E6R��Q)��tГ~ ��C�K��Rό�hu�t:��yM�p���1Vc�O�ׯ���	��4T�Kl҄D �v����+W/�3h<�l���K�
9�]�r�ܽ{��ظ��A�@@C_�(%'l������d�u �ʡ㸩�D�4�6d��\�F�����,I�FYY%漒��¢ym�t�\����\�V��� �"@����F:婁$#K��zd��<�N�nq��	��Jy?������	-��l6�����x�mG����2f�����@{��6b˾Z
3gςN:��5)��.<��:0-kP@d:#\+W��d��) �+���22n��pH�2��� ��19Y�B��Q#<�fx��	o�}Wg�{��¿˖/O�� �g̈́��ATt�K����wŃY��>�k4�Z��S��P��
���r�+�T�%{��a�!��{&�U�y@�O�cI����o�ii$u]$HGʙ3g~��Ǐ��5k����(��Z+՚�\TUt k�D⸌����L�C�1]\�~�#��0��\�)

>��,s<����5��%@ŏY�t�����e5Z��ơ�T�q�э���X��ɕJ���<<~�D��Or�*Ek�N�)( �+z���j��y�����y� ��f�h42��R|7����������v��ʮ]�����ɓ���B�ܹ3�iO~��9ސA�T���m���6!U�m�D��"�Ӱ�T�^R��
��z {LHdٱ����@����h�y!PRa����J��?a͚5��K��v��?�p�鐕�#��L&�ZPP@�f�o��#�L���HB�)n]~��0j����fW����={�LJ�`lF�
X��+�x���ѝ�I&c���>I�@����i�C��k��v�b�yEt�U/^��ҥ3���[+��<;�f�H��d����T����C���Q�� ��N�IO�� k�qq�f�+�d��/UX�T'���3�U���J�ċ/�xT��gM��嫨M$612@�ⷌ�{h���!;�YU�����hj<�"o�'£���Ra�n�������k���O��맜jkk '�	5?f��(N'�q���$���r��+����Ml͊��64�\�b�f��k���ku&�:'�ɓ'"H�����o���2�nބжm!�gJoa$R��>��NL=����YYYE�w���j���-�?��4}��'@��ѤO��QN�&��l�4j���HMݴu��ϩh#���Y= ��V'��ZjgϛK2h�Z����d�0g0_Ik浘�X�r0̈́y���������q��[BX��;"w�B���D�>Xk�c����7d�󏨳��`�*��x, �Фq����$k#\���aa�  sjjj�IO�����VRR��	ļ��w���U�
�1�o����[���7yr"U$�I�x= �5,Z0���rc۴m�����?��{�F���c�X�)])))�D�Y= ����	:w�N��;?]NrqS� �R7l w2���=}���G����O�˂<��!&���?d�H��!S�Ri(.� _��Ӓ�n�<�u�F-ᾩ�򖦐����:4!�Fӌ�����7�&c�s~��9<a��m�T���૯ެ�'V�[ڭ��@ǎ]@ �8���Z��f�+���^]#�s���P۬Yc���3��&oc����=}�E-`%MC�v��x��"ptt�~����4ꔏ�j�-M�D��V��LV��z�����!,�)^�烻��Y�`r�d�>�%�]$����s�����=|�cF�������Ub[!H�=�L�*����]>k�&e�	�[���z@���BՀ���k�\]��|�*'���|��Me>y̛4ʽ�o,����F~c1���vV�)"�u�!T/��?���ԮF͢��&�KA�<�����g)�4}��V���+|�2�4Q�4o�:��ae������z@��|�Z���>f2�Q.nv��A@��g<}�]�fq����,���VT��������s��Ud:q�0�3�����y�yCk׮3ܺ}����7~�2�t����E��F���<��-B��҃B    IEND�B`�PK
     �8�Z���*6 *6 /   images/a1588c66-a70c-44df-b30c-55fdbd854069.png�PNG

   IHDR  M  �   [���   	pHYs  �  ��+  ��IDATx��i���u�w����ֻ��mf��=�YD9�IKeI�l���Dސ/�cdB�I��$D�,�4����}n���pzz����}�yοn���&�83�7,�۷�ޭ���Sgy�K��(��(�DE��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)�됶m-�rr�W_�sĿ׎����s��D��Vn5��Ͳ��EQ�M���7�/�����W7� 
�N��2�.-�	�n�g}����tY�8�n��ڛ����&i>(�6�\�s�N�n�nӒ�{r꺶��;l�j���m��~S�V[���%�M'Ek/,'�n$��mf�$�y�P�;�;�U@��R�����*�S��]-�vՈ������1EQ^�hR���� ��q�f���R@�y,|���֡˥޸�n�P�n�ϒ�ǲa@Ԝ�j�j-�S��׎�4yUU�n�uP�,����~Ȣ&��x,v�D���&���ݲ�Zf9M��Ro�A�nO�q������)p,r�?ê*j�\6�ZN��N[66+��IK�'�*+���Òl�t�p\*}�)l��Y�-Y-��vIv��Z����u��gY��عeQ�_S�rRr���q>�ȟG�n��%Q���x����EQ~�QѤ(? )F.�QD�)�b�i�̓��`��Y�ͨ��aNְm���i�ږ6m���u�cLuy[r���)Y5%�O��zȨ�
�ꂪ�U�������[+�9m��a��R�_��P�KvP�"k�x��izDA���(�*9>yA@ESQ]��[��k��u_ٴV�zVZ�]�蚧5��;���)k����n���6����9?k�����W��vl�����q\�v��v�̥6�mg�z֡��ǁG�=������n��ޘ/���(��(�DT��RE�AE��|4G,���"����l�ͳ�uK��}g�Ԟc�q���������Ϣȵ�iX`���b�a��ˢ���?F�'�w�Z,�M,\��ڪee�PYZ��q::Dv�B�O+��
G���D�G��ōGgΝ'�&t��=�����x�"uz}�Y��I	1�A�̢�1���-���#�N�L:���vl�"jW		699��*�Y�V�UU|�1ǂ�\|�QV��<�/+Un��Ǫ��,#Ǌ!�����3<�(��;/y�w?����N�������VB��(��hR�T|_J͙�8ʲlT�VY՗X\�9N�ԭ�x�Z�-�}׵��u{u�xeUY"xPxd�dȲ�y�)��F-� ��-�u�,2�D~$2��,K�x[���k%5�IL!?���4�[
Yx8o�-Y3񾠼��Tp���yA��M�bFw�ܤx���pDA���.eɂ�F=�+;��*�,/E̐�S�ʬ����UC�|I�2��dB�2��c�"���uZ#�Z���ß����?����+��l���Ǣ�*��z�ucUM���nQ%�{�,⼶�`���g������զQ/���u��6��������5_��+��}k������`�$����Qk픢(�*��74,���)���<{p��T�����ES=J~���G���h[+j�l��<+ X��Vc�Y����q�ФˈD"AT@�,� � �����(��+���*M)��%"=��c Xl��f1�9�qL�k��԰�i�U��Ssi�$r��/h��K*o������JRjx�|>��ҷ*�m��J���Y�5Hӱh˫�IN�(��<r�2��$@��3g��%���sj���ҤQl*D�,�7��q����m�xo��ӊϟŕ#"Z�e��mce[[M�vi^v����>xG6?*��;�|�&g�Qܱ����������{�ng�tn߽{�~����Tk�E�a��IyC�H�d2��v��X��Ǔg��y�n��,t�������~U�~Z�.+��l�b�8B�ʦZ��-�O��TF� �e���JDP��R�%sI*�J�CŚ�fqP�QKd��E�>u����M.�.����}��R��[���F,�n'5�+v����z����sE4��H����!D�\�Z�N�m4�9�Â�����V�oס�g����mZ��ΩiE4��I#B8�|J��󊌷YJ�?�X��(ϰ�y^��*��kӔ�\�$3��@�i=������З4`�׬���F�3
���:���5�ٴ�O�o`���c1wӏ�ݵѷ�]?x>\w����,�*RE�K��Iyݲ*����Eq!����ٻ��]W�y�n��8��؎c[Mc��cy�/E�I��t�F�x>�J���߳ȁ�ZEr�b��J�&�f�E�ϑz%&�"˖��Bı]�.�V�XD��>�w�sX�����1��5�_��,r��,F���W��wD?E�8F����(*˜
q�`a�ؿ�I�?���ő�)�F�X-P�}����㴤��sZ*2�C4������,�}�o��4�H�����]~L#���w�'r�2��)-,ʊ��4��(d{K)�SC��s Jے�ɔ�-�)���ѳ�e��x��E�e�Ֆ�HR$�ڟ�ٝ��w^�{?�wo�d��;���ϝۺv�K��z�.]���抢�BE��b%���b��r�>]��墪�V���-׹�yްnk��N7�����ےR��#�e�p��e{R���P�Ȏ�(U�s�|�֬�H!��\�>"G�FA0!EwR,a#Q*~.���J���V�w"�+'�l��j$�TI6���K��lV��b붑�@���#���" &z�T�vE+�Fz|���C�9�_+�����O!�[��D�$5h�t""N�T��7)�.����3O^,W%BMT�".��r�@y��λ@�	������2�x���H=N*ʌ�;�����O.����9��P-��򪴜 ������ʝOg�׾�¦���n���O>qeq����a׿vv}����������_������v��P��� T4)�P�4���yV��)�w�"��?E��E�I��鸑��M.���(��h�g�m[�%!���.�DY%b i'+[J���qY8��#m�h�w��ǘ(�I-�Xl�f�G�6�Ǣo�f[H�!���B��c1�&�>�CD�N�{��:��^u�5+�os��W-��_8nD�X�ER��3�	��&bK�X��kBtL����NRyHIB�5&�'uX���)�����k
j
X0�h�����t�{�����
`I�HJΣ�|�z1��x��-\��s.�û��|PUԾ�2D��2��%+��e��k
;>�_���KeA��cv�ֽ�R��z�,+�,)�y��I��r��YV~�o�?�V/������^����>ya�uP������I��d����r��K��Gi�S,D>hY�e.}Ǳ���l���o㼜�b��]B�ͱm4ҭ&)iDjԔ�,,�"�[����ػI���C#E��*b�HQ8���0"Ƣ ������D� 
��+#B��՜)�^5š�Bԉh�Ԋ�����W������{�uS����4Vdߑ�E�K',�Ƴ%-�s�v":��A�4")7��H�����s����I)ġ�{!j�����
B�aI�P΂g�bu�b�m�B�*]�]%��L�4�$Uhzc�[l���>�UdB�n�h�hE��6pl���gʼ�b�P"���Ţa�� ������|�=~�QӼ��GA�.���ݣ�/��꽻u���~?p��c��������|���B��(ߏ�&�G
^(�������k� /��i�Ǭ���e��'��֪���l��>�>���}��^(�"i�G�)�n$�$�ܼ�bA=�#�߈ ���u��Kҭ�J�5�[�t���!�5��pO���b-�Hy�>�xa߭I���(,�
��VoD���W�$2���iQS[��;L��H��a��|�,NTBT�G	WB��nܸA��ܧ~/��'�}�E��@Iv�5�1��IR��I�Y+�ym,�Z0��2�6�y��.��V���d�2.�*R�hm0���VjMMJe���+�X�L���3�7�"�K���J�ҩUژh��\3��
�,��<l�_�@D'bn�k�t�BH���,T-*{񨂸J�L�T��-����}����֓/������矿�����/�?��?��+߽���+W�Z��(��&寜�|�./�&�u^7&+�g��:�j��r}4$?D�B�i(A��x��E0���s��M&����C < J
^�%Hâ&˒Uq�$"AuIIZ��\�D�����H����|R��{q���Đ��pJE0�X,��z�.�||!�Br$�V.�K��X��\ݜ:l�)'���2�$�&��*���U�,Q��?�J��lF�GGd7k,
��c P,{7S<�X�H��/�!L�n8���U��1�&Q+����в�(m<ڛ��_z���ۣg��g>�Az��:����,.;�J���li?��CZ�l�8�ԗ�q�qBY��*�2~,�����Y�͗�Ԋ�,��6�:I��"��l곐�X�E�����XJ fc lZ�j�p4�f��}��Oz��w��ݽ��+������S��ξ��#�1)��EE��W�a����������g�ے��u�b1M�bx[`I���L�F��a����"
�#=d�G��]|/�oي��x�PoV�����@F�tX�ث�q�DH�ȖH�I��=H�I h�`Z�����߲"OiooOćw�n�XԦ�	(�#JS���Yuǯ�P�ݜ�wkҍf�Je
�[��_�X<�KD��݈�o�����uBH�Q�dZ)5�$[�]Cȴ"����2BOA�DD�1uZM���Z�|=����2a;���{�51Q�B�D�Te�PV
)M�^�A�ʍ������J�T�"���`��,��_��T�X�Q4�����m�p
���m�zþ /�O�_�V�u{#\?���?�N�v��;{��}����3۟�_~��}~�7�}����+ʛM�Cp���Z������GM���(֋��$���|�x��ql��Hʋ�"E��*\�����r�ˋj.�R�$�a��������I���yfK����j�I��������?��j�W��d�z*l �>��ٴꛨRS�"z�1%���U2ϓ޸�]��1i:�W�7�"i�JE��[�(�t�EgF��:�6��E��
|�b��*��'٫9S����n�_'5��R�$={��x\I(O��~Ki,�5:��cQZ�k2g��`��{"�N�ݑ�D#��E��Z)��C���/U��O�+��8���T��#�����f���f��l���{%�4^P�`��P�ﲈ
�cq��X��R;���M���R���Ʉ�n��βt�ʍ{�q�޳/���G_�������ҿz≧���'�c�S�7*���
��RzWQ���W�O�Yq��l�Dj��\	'"���<G���$�j��Ѻ:q�n�τ��!a!ue�h�Gg�')&�M�HT"+�v+h���a�� ���_��W2C�������/wY��:9������a9��8+����MIa����N����X&��T�DX�M&���u2,wu��)l�ds��)��B�G��DKb�ލ�8����ܠ�\�ȡ+ή$݆a^���Ĺ����ϑ������V��r|���洱֣�Q�z,�l���_ϖE<��6��B�Ƕ�6r��j�:���HP��$�)�y~em�xwv�i��]ڿx���ܳ���s4����1
X$&��Zf)�YPMSQ,��,��	�|��7D���`0����Ή���ߧ��]�O��z��t?����?~�����c���׮]k�?�U��(oxT4)����ޝ?�U���u���j�i$Ǔ�KI�dF4���Q��N6�$6����$��K��J��?a����9�.8K��d:�5�W��`������]�j3^��+iUk���8��q��g��D��˕�)���O�ӡ��_u�5��j�}���v!��^Ti%�Z#��?�1�k�{�4"ca`�X\��VE�(����9ƶ�Q-�c:�Pp7r�`�@p_0�*K���٦���f��2��kE��E
f����೐c�X�#~`=��:_�)��6�t.�
_+�-�?�Ңؿ�V�J�}j�-CP�G�����n2_P{�6m�Y�A??���)
`���N�V�F|��$�N�\����ir��������c�=F[[[���h:Ӕ�S��ɲ|�/��+w��~�������y��z��)��FE��P�E۽?+~n�f��E�[y�t����tf�a�Ð:aW�;�'B tY���S�	B�nۮ�x�+6D�I�6�J���(W��JCd&/Z)̞������t�!�VJ�Tkăc�ͱ�W9��:��HO-r��Ԧ�B�EEe��$�E�4>K'h��i,uB��%����JA,A���7D����o։��)���B��o�q��)זk��x�Y�+Q5��n�,��R&������,�#@=..�;D���"ڄ�,H�)�ײ����^��VE���״�Brc9`��Z�k�� �t6"hZԪ��my;�M:<�Q�ۣ��?���:�ﯦ5VEB: �~dal�زX�v�����ԺeKqPOҒ�gsZf�ɂ׌��+��h�N�Νc�AI����c����o}���C7��}�����������3g�%)��DE��P��i����M��q^v��2"�mr��An7�N'�0p�x��"��Ը@4��&�}i�����KNĒ)Ҧ�H2&����͏�Q�5B�#<<���(_y'����b����Z)�F�K�#�������&1����8�,��n�B���;MF���}҉g��QlnF�H��� ���d�"3�k�m��ý,.<2F��rM1�O%� �ء�ώ6h^4���5uMR���NU�GR��Bxd1~Px����(e81\���1��,�
�w�<��I�5�Zm))Q��I��cg�+����E�t��:t��UX��IAQg��ٞMs4����)����%��HG"�s����)%�8�!e�פ���ĎYH/$���Ⴗ�\�Ģ���P�\D�a�.\�`���s'��ٗ^��7�ˏ?��;�����o?s��G����PѤ<r�׋�|��j_�RV����@Z�=�Dl^��ܤ�l��M;>�~�|�^ENj�8��&AG��M)��[b;�*s2n�0���Q�?�^w$.ܰ3�L���G����q�.E8�V|�DIQ�IJ��Vs�LwY��~ו�D�e!��~��p`��ʘo��ZꢈR>�ZF���ɔ��)\��[v���	|��6u�U)z+���7���Pp5߾y@GiM�����[B,y�1�2o�����{���h��K-T��"b��๘����Q��(-��,|:=���J����4���~
��e�S���Լ-?q�G
qԔf.���|��D� ~�����B�_o�̲���Z��Z�C�M�Pٞ���{l��1Z@�y]�>b1�йs��<O3Z��Z�}�<\���ll���>�G�ӷ�ӟ�GY������?y�ɭ)��BE��P����U��c�i�.�����Ն
�!�x��X(Q N�A���8]d����~$���0VOf��*�$�>�>�'VG��eCE#K�&�a�&�jH��qTi)�x�u"�PH�ȑ�X��X�t�/ܞ�3aΝ�r$�<g�]K�)��J#_%��D�@Ә��N8�1t8��`���E���#+k91�si�&��.	��������)p[��q��JRfR�Q��	��q����=��2���hɪ,���:�`��o�`򈞸�E�y�2 \YHG=kbuX���	�}c8��8Zߤ��ޥ�Œ��t]�H3�a��KM��@�ִ��ǂ���Ad����Te	��-�W;��@�w��\�\ҁ�.��|�Z�Y�9|̑�ɹ�2h��t����$��&�����^D˄����{�o~�&�	���鱋�i�X�1����&�1�Fk4���#���&ݺuә�Ɨ��g���G��k_m�O��B�KQ�7
*���B@���9Q�����%Up��Eʅ�d�H��7�lKt&p%�m��5I7���y(ڮJ�\��ߠ�
⩱V)9�A��96����beܶM�Xk�1w�WWKj�L��F�5"� Z�)Lw����a$����i��+Gk+E���6x�!&o�e��yvH�I̤������b��G����ʌR��X}��� ]�
��wali�U2'�Eh`�n<�`�9"R�-KKā���sJ��9�%~j�,u�ŔHCy`��C	�qV��VS�H�G!;R�,.S�'����N���;�i^�,�BjY�5��3�[��߆�C?��z���:H�j�Xf�AX�XlOX�N2�g�S��"��X4�>�zCt.��{5�!�*����iY��4�!�Y@���)X(0u��v��oݤG����B~��1��>��ٔ���T�s�!Z�Е�\��l;}���^z����_���}�կ��y��U8)�M�C��식N���e���O8a�O(�\6�IY���I�D(���㣉��ц�k R,�$]�67�8����d{�V��ޚ4�D\�Z
�1�Æ%���"�����0[�þg�(Q&�2��	��&��R�p�����V���I��Y���-<椛�Z	={eU�s'F�(>N�yv$��G6�;�F��Ll��5�g�ᕹtˡUNR��I�aL/J�a���~9���Œ��H�/b��^@���uNn���$������s�aښ�.�̒EU�y��o�Geˌ�|��Jg�C%5K��c[�#�^c1�b�*!��Cj���C�G4����Z*�ݻ�G;�5�v^O��X�e�����B����!9,*C4 w�	וN<$TS��mB�J}� ��hH�?���R���E*#\ tע�O7i�ץ���'{�',�豋�h��r���w���K��G?�s���`Q�7*����I9����w��%>��.9�@�=-��
�J�>р�	0Hy٭��������DCp�h�W�&�h�[��vR�M� Ja���"�P���P�->HU#�a=�e:f^\��R")8��vc�su��4^�Q[��Wk\˥�]~2�Ε�����ӓc�*�϶M^��R�a���T��@� Z�1O�B1:�Z� d�r�F�")�B�lpLe[�bo����?��k0��<�p�X\�b�Qds��"B%��Ř5
����̫[*Ft&eq[�u/��"Q��-o�-m�$V_7Ȝ���P��ū!cQ������Ļ�%o�U��}��©	z�̐� dA�KJNC#~.ml����v~L9�b>�"��z&R���)(1�O�$�(<O�1ᩫO�tm@k���&����Z���7�QH��E:����pB�]~Y*�]y���s���_��~����2� EQ^��hR^s��|4^�����I1�E��Ȫ����2�)�\k� 2S�1�I��.��g��Ɛ��׬U*-�DZlS��"D�3��Dkj�"
�>�������*����b�|����%͇���0+1>�xe�(�օI?�U��8�u|jx����xO�I�8���E!ͅN�͍y~(i57������$����*2M!_S���
����>��Z�9�<+gt;b\/�3, 
3�,1��'Dbp-�_��K=���I���������8��m�
V 9k%��-�?�F�_��!T���;�q��J���X�Z�'ʤ�G��1�]�͂���ߔ�5+RJP�����bBz�EVEM�҅3t��E�6�d�(���͗	��xD����8�2y�O�У͵!�>��k��K�[ͯi�����>���Ǉ4[,i|�K��1mllXg7�Dd��ws?���^�o�{��R�u��&����2Y,a�#F�X�jV��<VK�D��� *���ot-�ENߌ�#/rY&�`��[[��m�'�B�3�hB�Q\�V�i$x*�f���$�ī����z��d`�Iљ�I4�]_!Ѡ�.Ă-�N�c��MD�<��5#^PkWl)To��i�7�	�O8��d'��j��8f�Yf;X;ާ(�k�y���hNS���y�13�jn
�!Q腔��.�b�A\��r� ^�߇RX-�ْ2d8G�2�J��U��D@D%�<��6:4l�6sX�ՔI���s�C�ۣ����\�iY3�J���m��,`�n-3�0�i\��x? =ɯ-҄.�Ǐ��tt<!��)dQ6��t���}��>:^�����ծ�u'�R>8l'�/i6��Zǣ��e�혱5��#jW�x|L6��n4��ut)I2*���^D�0
�����^}�s7o���˗/g�(��M�C����h!$\I���|F���_Z�Q�CF��&	!,��xjk���\��LK|+f��8�cJZ�A<�]�fU�BIm�+
�tq�P����y�=Vk���Q$]����_��_�3O̔���.jnx�'��f���5�`<��j1w�<��zI#:���d��(D=��wRծ"@����wz� ��E�i��P��#;v��DA8���H��UW�笺�m��M����/�b�]����/�'©X�������c�,�|�n=�xImp;G����$;N ]���,��\D�+����!�n�pN��1�ID
�5��\�v���z��{��ƥ��hg"nas���t:����#xM��E��ɢ%ߋX�w)�� ��ʽ*�X�ш�R}>��x<>���	�|�||�4-8�ta�5�.�=��H�����~�4t�bJ:�0�6���_x�����?�C���nQѤ<,�(�C-	����0��݌G�P�G�WV&�#�^�2���ˑq��k�tٝ�)���-3�P܍�%���Uj,�1]�j~0��r����f��ڡ:/Y��"~:~G"
��{w�TRtn�%yA��6/Ɲ@����+�NƂ�[���bQ��J�"b�ω�0a���\n���"q,G�Nj�E�8�P�R�O�4�񢝦tn{���F�h��B�������I�'+��-����Y1y�6�QM��k��?m���%+��`|iWUi�|�����I��ϖ�|M�Y��Y�v���XdE,Y���m�ő���k��I���:n�{ve�ʪ�Y8!$��u�����Y���+m�b���$��X��y7�C�T�7��Pp)���f�E�w$��$��㲐l<�{���gc�1���5D��YVI]Z_?G�ݻ4�="�/b�ב�g7t�,CXb�?�/�l��Aߣ(�I��I��\�_����ڵkןy��S�(�ST4)�c�W����h�F�Z�ő�ʤ��jK��DmD �	���6R�T/��Њ�Te��-_S�,8<c=��i��K�)�֋ �݈h��j|�Wjq�F�9��,xPP�dRb+�U�xġ
��nC����C � xPǅ����I�U�VG,p��L�ǒbq m�D���v#���i��m"d9�PS~���ڻw��ަ3�V/��lm�<~���s�}�T���*�7������a������$]i�r����4�]/��oiӸM];��˓|����2�Fu�w�"���Ӫ��_�u�r�.+�^`�����OvP[u�Gn�^X��WE_V�k|o�SO)p�_mV���L���+#S�v�}��O5˙y��)���m_�LO?��wi��t8���Ϩ?P��2��cu�(Ƅf�E��#)�j�,�r7I��7�f����Ey]��Iy(�v�p�2�@��˂"�S�� E#�D�M�&�� �� �dy�0�R�˺���KR��A-���^��h,���m��y���)�t%��HP�R�Ŗ��*,���s�B��<�4�%R��t/����(�E�f
#K�>uB_
�Qo��D�˸���*ia�q���buG"li���;<�CT���c�4�ڔd���)�K���hsm$c=�_�N�����6O߽w�?���/=��������O�;�?|-^W��1��EY�b-cbn�y�������|=��,�<�:iY��t���.��A��ϲ(y+Y����aA=�Z�ϯ�S�0dD*�Uw%j�|��,�IA�/\ �ь��H(���*�|9�����g6i��ѮM[gh��Β%MgtoL�NA��y���@�`@��1|���5겈������?I*��u��&�P��܂�4>���J|�l	�@(�?ԅ�42�f.YǗQ&.F��_�I�eYJ��LDOo0��Wi.uR��BA.L~�h5���
{+�A�N�z,BJ�1�ląF�^L�<�1�������
7aB��+����
�xH�Q+F�R��_�*
D8(�^���QǄ"n��%�ɩH��P���f�
jxlߕ�b6-�|%p<ˬ���}
��66��ɧ����ݿw���w�"Ͷ���{����}��.���7w��'.�����E��2�|�~��Q{b�η�Ydmܺ���|�1Y�kղ����ۊ2�)���*���f�Y�+t��0T��������|��YL�U��jX��lK�ѐj��6nX��!���HY �z��T���is}C�o����$�Y|�k�/�cmϒ���]��M�)��M�C�u�$/�S��9GRTQ�f�u�����U����G���՛Lqt�唲�p;�&���=_��m�9H��bD��&�Z��BQq��i5��p���UWi���!z!���M1�́�;�ҝ�4�Ni��'&�[����Ɔ�bq��BWiwU�$�h��ד��մ<k�lޢ^+��1&K^�m���y��M��J���M�Z��F��}��h����[7�x9�l˺x���_���O������3����G�:e�Z��J@ri��ڵ�az�����{�{W��z�_��q�\���	~������� ���ݚ��f�<�d0��>���:�Y��@�6H������
��-:<:���]�?<��l!��F�����
:~ӉgŇo�f[��&Ey]��Iy(�m���|�l� P�#g,B?d���@As%]a�bA�����-�V3��A�J�1�����;\#���H
������\�+����,@J-.yn��NW��,~*��XF,t���z���O(z���"�)Is^ �t4K�0�D�-�8=�GF�`���P�Dƥ&���l1��j�`���y�B]UR�b2��A�[bItx�Bi���t��K��t��y�/hkc�.=�V�F��s��Ŝ�c�`<����_?�{x�ċ/��?�|�ҝ7�K�3�X���6��=;_�����8�L.����b�\����Y�?[W�E�	����g�SV�4 %g�)�(���� dG|�\����}1"={O0����]�$՜e��]��Atu�7Ӯ�.��CE��P�j�#fS֕e�fو?�[�E�����ŉ��@�+�<�h�ޏ��ؗ�E�ܝ���Dg,����E��t��	5F~�z�@j� @Ę2Ii6�I���P"�	]���C�Cqx��(�2�Le+QV�X[F�D���ြND	���M�r�;�)����*[q����Â�l���s@��x�)��d4�BBR�a*�k)EK�d*~Hk��y;>�=�r>�Y�nD�3[���I7��BQ�|r���������f��S���q���/<��S����7&���[·C,/�urw�����Ņ�������]�8{6I�KV]_��`E��{��hjL|�FFK
x,��}I���ۣ�lL��]~�Z�I��xrDݰ#���C��`8���������x���*�+�����k��&���K��ݗYi��v[����I�7�Q�,eDLiBT&�
N�4�V�a�,�d>�f,�0|����(Ķģ)pL	��e�om�{�h�/b��_Q��(/Q���F<a#i���hY������}�Ytu�X�k#���y!���{!K�X�����<�gqF��R�ER��?k>WfF&UȢΕ�@S�$�a�6����wD7o\�jxϻ�����������lS���x���;|l��X��V��eL�3�,�������'�`o���<���|8�-�×^~�'wv��c)��ݣ�s7:{�%oxV�����&/��~�z���r}���ɣ��C���S��?m��7��Fs���S��Lg��+W;�][��|L��C~͉�l��#�\���1�,�i��G�T���뿧=Z�%��иֶ���z���O���e��_�����7���s7��p8U��M�âr��fe7E��]��V�!�e��QLk[�|�\��\ƥ��7M-��
��,R��[N���[G����Wj�i>��l6O&�8��ʚ\�g1㊠�ՑuE�fҟ�"�D�̗9M�}r�&,�R��eQ�Q$���D��x�>�,�N1ˣp�=W啤�d�0<�B����$�#>f��ӡs�'d�q�,�s.���������)?gF�۷h4R��%��,Ҏy�����M�<\����v����Ȯ��L��'�g�r���O��_��|��՛�@y�h�W�[;;;~coot���[���<������ng�c�V�q'�pD�t�=�Ai|�����?�Y_���-��p� ��,S׮���"�������^{>ݶ��Wv���a�_e����ݛ�������~��?��s�󉝝~��y��)?M�����n�(#����7DW ;:h��8=$�([�0��I}�\R�2P��|1<��F>�Or�y�XNi?NEX$�X�Y�sA�8=�y��b����(c?��`W��l���H�m��]���XȅQ �&�?� Y��(��뱈��\F���A�Zߢ�׍{�$����Ik}��"���W%���Y ɔS��ztt4��=��w�����T�"݃�B/�ud�-�9�A�a��$�L��qF�3OK
kK�{|`��6m{uz#ZL�(Kbh�������kW��������?��~AorΛ4aa����ï]�����я���/�I�Ζ�A7X�Gԍ<�(址��k\�c��Kg�P���x9k��A�?����i��S���l��7�Çm�=�FֱU��xc'�/���W?x������g_�����0U~4PѤ<,�*v��r�kN�ҨQ�K�L*�-�wyHYV�\8�T�LfR���%x���߅ߡß�1|uN�w�D$IG>·i�������0]�BBX!m�`��x"�:]c8i
�=�GB�n.	���,�����}�G"E䖕���٫�k�c�=��墔a�v�K���ƋL�4�v�ɦ�^@��'��祸�C#�UCw��������c9��Ęd��@�/��(����ޢ����x|H^Еگ8��i1�ϓYtQ4��!��[4���x���6u7�g�v�O����k�n~��/}۲����"AK����ڗ�u��;��?<>��R\�l�v���z�Ne�O�<�H&\㓄v��`mD~���躴������3H��ۇ����^�{��'��ss7�Wd��̘�׵�i5�^�PUe����7���|�[���?����헾���Υ��S�"*�����',H�>/c�Z"f�<RrI������ӭ�|�0��н{;4�)^$TU����:�@��b��b��t���
$��q=?2T�qetKM��̈&L���#�F��C!o�s]h���Q�������'���kEb_�c%��?���G�3����)^�T��10v�oS�,�|�<9��=��k��W�hclL�"����P1ڌ\W��ÎC]O�ߠ��[�H�aU��>D�,��h��h]���>t�F���r��|��_~ǽ{���+�~����o�Z��J@�����˷?gw���&���Ko�&�`��7�p/�#t�\��xn���6��PSE����dB2]~�k ����8y��$�{�ފ������OE�P���p�:�3+�ݨ��ss1~z�k��[߾���?r��~�ڵ�~I=���CE��P�'�i\��旅A�u}�p%Z̦��[.�N+ВMAQ���G�ٜ��ә�&�$D|<k,�I��u�"�}LF�X( ��,�1-��$ɀ^˖�n�5�m��0U����G["��e&�M��(�����w)�:�6�����(`�`�������S����VD^�ɰ^���������@F|`܊�s~\�Q�PJ�m�-����(��T�ce��2��V%�7�Xб7�'4�-YTZT�"��0)k[������{~(�U����r>�����{����o�إ��c7o����˗3R��A�ͽ���m���͝ۻ�����߷��bv$�b�0�����:Խ�IJN/�k���}�drx��-����9��=����E���$��y�Rޘ���⭐���H�I��n��'�|i�xtgv�#ߺ�֯����Ý��}�#��ST4)��n���N����V̖C���x,5BgϞ�#�+���8�����n�/"�b��HSV4Ҳ�&�G�}�)�TRo��(� **]23�\*-#ǘ_z0|n$ʅ�����Ӽ���)��b_ ��A�#��h}M�p�Ʊw⻲}t�]�r���J����և�F���{�E*���71p(�]�K,vBϓm���&�p<�X�M+�D�_@����!�`�������X@Ř�WT��)o��n�P���B���ˆ���yz&ϒ���^}��3�q�;{��-Om��O-4ea8{֊�}���G�kw����l��/Ҭ|o�6��a`�M�~��,���>]���]�����+��WH���ն��vӟ�3�q?�`¿�3N��Rض��5����| ��Q������;oQTn����Ζ����ƍ�up�����>��<~�;˫gǿ���7-*����O�a���i��CU]t�ʍ���!����X,��ξCg� �"C-�АrZ�HMS�;��` ј%g�歌��ba!��RZ6�g!���M����Lf!��Uq�nmy
��/�Y��2�*�����F]��ޢ�W.Q����l�bш�9
Α�)x?�[[RWu8�ҫ7n���=�_�D�.?�����O��Fgl�%��,�� �Z���Sw�I�/�u��	�N29'[���禤2-��}c�#��vP_5[�!g����
��tAY�HZ�	��MrÐ��DF����Lӷ�W��w7���W/�_�WY8夜��0��_{��ݻ�w��e��{uS��:�=�!���H� Ҭ����Z�doA
IE�k@F�v�G����q�ЄoS|�j=�!�V�o ^"J˿dQwHx%�ILv][�`��76�t�3������|���_|��G�7�}��ō�w0�M��&������Q��"���m����"����/Ӎwd�"J�k��7/��ؼ�G�z�tō�ϗb܈$H�cL�	 ��֒���Y�HҪ[β-�Hy~ �i��8����H1#� VP^Vm�ߦ'�^���p��<�<�Ķ�����f���0V����uYD�9#f��oݠ:K��O�3DŬ�$������xK!���qf9f�%b��8��b,C~Q��38��bK�ӡ��1��j�XR/rXxi������O�傖�ES��n@k�.�]�Q�?_L&T{�6�D��=G����W���[w�~coo�gϞ}��?���+�t�:�m/��n^����zD���T=:ع'׼�^��������~���y����i��8oiQYT٨ej�����1��;��߭2�>9H��>�k�]���G���ry���G_��K�~�����]~�O��������:�̓�&�g�I���,��B�|��ZGGGR��O���Џ��>B�,cS���T����;4�e "1���ɂ�H-�KH=����C�T�Z�V�4)��&�mV?��&�r1LU���8�E&)=��j��z�;��3��4����r�tC��iLy��z�C�����^�u�Ξ�@��:��R�{��K!�x����$E��� ئv�m��uB��B�����s�q�r�2�N,J^2z�+7�_r'b��2�CД��ˀYuH�,��ɒf|�{,�����]����%��}��ʒ�߼�s�LVTg��<�ͧ/m�a������
kя[��s^��y݈�Fq��re���L�i�_�H*�~�|������e��3�[�(�d�h-#��ϿS.���wF>$Y�G6��1����l��(�_p��So{��V}�V�x��/��3/�x�g���ؿ���?�����.��QѤ<T΍�{u9�_˺|v2=~��xl�X,�9s�:aB2��D<َ��	uYZJ�͟�B����RW�ѩ�d1e�;��$�A%7˖�a���-�J)����e��u��˿!�Ɍ66�hsk��MX|��aa!�x%�]%m�T~��{����ł�	3�
�����HXj�<p5�+�=>O>%����iN�,�����r��[���Hu�"��6���Z�|}ߖq/��_T�'|��0�"4�Y,�4_Zb�׹���@��u\"�t4�9s�R�;��l�����������;��7>0=���������k�IR��������"���m���L�� ��Rq�/-~>ֶq������a��=q�p�SK�{�V��Ob��>����nV#��JŇ,��y�	׃_[�K"�MeY�(������`��W~�Kw�~�S���Ǿs���Om���M�C��{m�����?��Q�w�� ځ?d#^�+�d�L2((�F��e��T�q�F�	�HR4��Hל���@�ء��+YD��5"�d�X����_��忍&�A���)o�ӊ��-�N<�W���`
|�������8[��෹�AϽ��9Z��O��R���%Y�U��C|Y�W�s�H�O��S�N��:Z���sC*c��X�\��n�̀��%����$Y-�X�T��9��G�k��g-ፕ�r}J������yB�n�x������S�O���q��������?���~��,Do[o�ł�ߙ���mn�t���X O�1��T�k9��}9���������)���{��P�ý��ݽ�?1o���?<5��ʩd�Q#Z��C�d�-�$�I�䴪�leP��a�|���s\�V�Fg��Rz�N����o���o����ߺ��O�<���?����{�`���:l���;o���ݘ'��P�H�E�$%ي-Y��ĩR�SI%�T�W�#?�5T%�3���hRIp%�Sw��@��7���y�^��Ҏ�")����.���;�{�w�����^k��<���4-�}lhZpx�����&���
�7ٶ�Ky�%��ʑ������$?�X�t!y�U.�tY��� ~ `��X�^6��+t�U�B/�J�?�|#)/T(��R�������iB�'�|��]��9�(���� 8���R��]t��vMJlX{��;c0���i*K���&?����9]�;����h�2p��ɟ����$�8D� �3�N��hYb�a�
'h�Q�����e��1@�&D�c�����:����d`C3��?���a������@-
�N��Vw���߿w8��3g�v�]k>��Qmeq�4]��[w�nђ�)4�0s�uOʭĘ'iZ�����ywv���w ����ᛮ�
�9�Ȍׄ(�e����� �\��Rqeg�)�#�v�i��+)�)��Y%<����<]�5�+����~e<<q�o�y�c�}�[/����]�<L'�W��vo��M��#kk��U�o��>���?�O'�Mk�s��mYH��.)v.;t��ȮO#u3����Ґ�z�ܣ[� �BGL�f��*���⿣�_��4
�=w�rM�c�肎����m~�p<��h������?�|t����n8§B9v/Q��^3$�o[��QBU@��1�#�\>��B�,��hB�Yl�ۊ3d����R�Q�S�b�Xɤ1�!>Ou�V�
  q3?��`6�E�%8�%���:�,�I��ŏ�d�F����)�����O+J{S~?d����6���E�^w�4M?=�~ҟ�?��S������'��aU5�����<�l�靲05��{�)-���׏��4�*m,ô�]������Iy�-��a|�(9um6��a\�s���`���#��iST�Jt�@�,��s�I�M�L��Ha�V-6S��=*�A���̶^��'SVM���jZc����/=~��=r��������߿8���v��;{�/�O��M��#����3�ww�����O�0�`��תּ�e�mC3̺���x�^	G@嬼T�m(둮�K(�U�&�p��X����)�����o���lT�I���մ�2~���� �"*�Q�2��ŝ��s꠭�q� fKg�e�B�6�~Y�
�	�m�S��I+B77�r��~@s~x�k�L�?�tFyR^�m;�3%���*WR_@�Ǡ��e�ԓψ���N�Z�G�Х	����`���AH��A�֚45u!���`4��?�7�����@y�n����s4�Z�D[q���_z����g^���;Om^�gQ�Zړy�����#�~�d���k�ꔵ����!;�,��Qk;GAР%h�;���ʻpn�Ã�|�4�	oL"��$!K�t���$�쑦2إ�(�!{����Z�:i5�+����ʍ[6.�I���{�FЦ��8��5z�Z�*[��o�}���g�����N|m��֗U����-EM_�c	���G>n���b��.M
���п?���q�~s�kz��J$!X�2�� T�;HC���s��v� o���vR���n�\�Q*�'�)ƹP"�g �L �)�(���'�����vMz��@�� cI��=�O�Wk�a�����!��|,%J]c3ML}�7\Z+�RQE.B���Zߤy��8ȏ#q ��xC������� @rq�� ��]�J�Q�l6��÷��A�f˿,�9A�=#��KW���Ө��8<���$��i���
��.�	Ɵ���*��5k��|>���t|��g���f��������A���,�'���`|[�	���'�[r�����A����R4�6A�6�L���]Z�x̮On���͍�ҵ��x���X���Ipǽ)ׂr$���=���n������N�!��J�<��6E�aIy�5��@v$�1ߛs�@�^��z�8�;��w<r�c�������+�ַ�<}�R��u7��i9^c����"�-��W��x�����zZݟ�M���1̱ �UD��xd)���*(?:��S9/^(��6Q��,�t�2N�s(5�p$���?�J�M/��6���o�z�腗�ʵ]2m.��[����2~��Y�DG#�@��Q��Vs��No��ZIU�CZ1:���(]jv��A�ƾO�`��-��P�Q���)B+�#̂�� ���i~^�T�pW"���{z���砆g�J� Y���D�{H�R )���I#�<��;�)�HQ�+E��WY�-rQJ^�km��K�=��[�Z������=��zፖu�%��0����dE�W��T����g�ye����R��T� r�a���v�}���Gw��ك�����[crL��(�I7ߗ���'�x"N������蚢4�ŕ��"���0Y�̖�p��B����f<��_tk&eaLoxl�e�$���Ԩ�Hk:��������K��鋳��߾r�~��qj�}����xy�_c	���55v_�y�^����˃�0��H��mi�ݪU�	F�i��a�Z��#/*��\8ObS��CIIB��Y�H�o5G��^��B�ːL}!��Z��C��~Q�^�B/�d~�ͧ�Swx1�,�d�[΃���
p3_~My�'Z=�[��.H��D$0N
jt�A��J�?��5x��h8:�Ş�H�I������WKI2�e(�ٞd��zo�O�z��M)P�y(��܈s:Q0��xV�@#J�����J��x^���ίt� ��98�"�`ۼ�9vZ��:�z�����s/�����y�'��fh;��MP�UՋ��?1,�p��,�w1�W����u���nCcx�[K��&��(��/]�ݻ?�>Vv�b��4�8	��\Tk��R#��J]��T���7�Zk��^����i�Jɋ`��j6Ņ M(Ж����S��'�ry�d����$#K�k^�Q����o}��?��k��C���g�w�kܺ9Y����4-�kz,��{x��������&qg�M���2��d��S�f�����TJ�@H�����R.K�22B
v-B�^,���P�h>�{Nߴ%
�uע�;�T�I����vM2��Z�m�O'RV+x4ZMlI�P���cc�V:MY�d�R���#aF�yFe�J��}�����^w$ͩfU�`]�N���Լ �d�@�	�!a{�c�"��ƕ H���lh���&ǹ!�qKN���@�b�����q�5e$�����X��u�̓)0~ ��[=��٭N'����MƷ�y��o�^;|��K_��ĉ�׫D�Ew��5��(�b�T'M��
��J��֬Q́]�6�
K��4�J_�%h�A�>��L�O���#7���&�IF�MapH
 �rO�Rz�!�2ѢA�A���@f Y$E'�����G�|ŋB�
M% ���q�H�[�%��t�M�13��D�kK��	�TC 8���*���q|����SO\�?r���7�������KK����X���x݌Ev��WW/]��W�a;)��8Lo��i�ߗ��-�{�VY���E�+!���^�b�T�"gK�Iif�x��l���j�g�a*rP��"j����	��6��0T��I����As8�z{k�N�EG �tm������$�KW��K�wx�Z����EM�Z�hm�KZ�A�f�9�y���Ç�ĥ} i�R�L����nq����-�$"�Wm�2� ���N���  J�lQ(�X%�|���M�04�4 $*<yE� ¯��  v�s��C*�>u�=��[V�վ5	�����G�;��W�����vm�бc��멣�� ��[��?�J�2MC�lg����`tH$�yX��d���L#4ʛ��h�f �j�����`~�j����?>/���o�Y��x2V����5E���7'o�P��D'�B���d���� ,)ە�3��L��ec�,0����H����HyH�[����rKJ}��$��%��:��\��w_{~���]?x��૿���z������e��3��i9^�cd�����"��rn���Ma�5������-I˝��^UV5]3mݵ4@X@�e��� ^����b ;7�+=WzMP+�E�?�Ȅ$̬JH�j��R�V�.@+f`��o�ק��K$ldyl�p�slMF	㒌h&��ҵ�t�E��K��r�n;�M�Wy]��6���į �X�����2��xx��{�yr����u #tV8�|a�bppX�m��D�T݇�T+D�fA�_��
:U5ٱ����5�m�#��g�\�3�~�ik���ը����$���}���0��t:��:xB��x^����QBf	�8[tjZ"���Z�F:� ��dY���4�[��������\N?~0�O���A@4+�� nQ&|ð�X���?�)+ C �υ@(C�����3	v�$I�-J�"�d,Jz*�
R�λ&��#!fټ`�	È"�@AޣwR��}�	��M��1%�*u����6�,ژ_:z��+{?��k_<��?zj�:���F��<��i9�0CS����=5�L>7
� �O�q~k���f9�9��m�ݪ*��2 R^҅�����&eq$Y�z͕]k^�td<]wų�h9�F��,)m�C��g��sL����ɥT`����d&�W�;��}\������&������]t��&��]�K@��֔E�>���:2 �����u~ϜV9����d׬[ ��(��QA���O�(-�>q��;y��$���Y�|��� N8��BF�Eq�_oB4�0J(
걐ѓ���8�=�z�u=	�������:;�����_^�|��'N��5:��n+���)K�%mȁ��1�/ (�jY����|�˗3��W�iJC-��5���è���O��tD�a���Π�ᙔ�D�㪅m�&s���.Fi���Su�q#���'���T�	C��*U�F'*:W�3d���:<<��� NC�������-�W��1 ��S	"��k�X(�gV\ew����gZ�?�?����[��_~���c)�ZKдoȱ��LHu��~��lV�"}+��� �O'i��4)�,�j�0�>/t�nZ�k��n7^t�ӹ,��^C�� b� q[�N-�&��Ż��adb��0xOU>C.��t�b]�x���Eղzrr=(s3��n����F+}�NF�n�R�Q��`HU`Q˳�8T��i�MVU�B��A
vэN�"^�xMZ���{ԮYJM�wt��wDF�m�l-�uɨ�S�e8�2D��+K��ᡇ��c��ɟ�4���h(�S�~_��a8b2�5�.U�ԍ����N�g�ǂ(~���/�~�m?����kh̪j%���2��T�V�����J��
��
��:�(HYh�T�
�ʦ�4TɓASaY.�����V�y����gd섺��i�s=�s�o7Ăh8���g;�E�e�𮔦�� ��؀H
�"/��u�BT}'ZQ�^H�(��5���f����m����'����5��[�%��r��0��ESD�p�Y5�7��e:5g�������'�<0����7��2��Ԙ���ˮ��X���xÏE�'Y<��z�A��5���Zy��(�3
��y�ߤ�MF�(�xcx����@�����d6���C�1����:9P�ƣݦz�I�Z�פ<7$m��D�2X.I��L���N�l�J�Ɠ�c_D/^<��V��h��$�%L�$���2��v]
yUF�p	���$"�A֚W���g����t4����j�E�mIY!H
eˢA�I[�Ϩ��&�7]��aC(K7u!���
_��PV,��!�Ҁb� ��_�Ѣ�ʺ2|_����W�=��D��7�?��F��ܿg��?;���x���}m�i]w����(I����ү��%>M "�S[]���z�ҡ)އ7���r�	%*���*p]s�5]�|��t8��(L?1J�f��
s�魭-��M:�L�<�'��AcH\��P�@4N �j�!�L��9������8�-`�dI�`�f+�R�N��2,�A0�=�V\���Zd5�B)��7�<����<�Z>�)o��iL̴u��9����{G�G?i^��uW��5��?����~��_�:q�uZ�x�y��%hZ�˱؝E�8Q�@��d���5�T�go7M�ci���Ҍ��Յ�����J���4R�Ψ��Es�R�������1D]�u��%�$��H�v(ED8/�Kۛm�Xi�p�|2��y�נ�imv� �R�b;�#���j�6��e������Z�ڽ.u:=�gs�����^��xDk��.�i��8�R����e��ECJ�8�~x��K���tF��͠��>��ǻ�X�PM�����C 
0��s��k����@�gp�5�}T:n���O��c�뻏;���$��&�:=�z�x3�C</jAL?����{w��R<�J�8j�#�	
d!�s��s�g�*�� �E�IF�A>Փ��j��Z�{OTU����O���� ,�y�00Ѩ�s�5 ��&�K����T�1o*���_�U(���"��-:�T��ʨ�]�YV�f5J�B��*�v�Ϳj�F�~1�?2s�ԬvWJ�zi�}�%]:_K����ͤ�Dq
q"C]V�H�X���!��fߚV7l�ԭ��VҌ�Hf���l��]?����s߸?�;��ީ�e�UKд˱�՝7�@y��|d0�zxx�3?�d�]��ԩͻY�t���yW�n1�
]^��0���t��y!?���M;�۴��Jud���3xG�ky�
���QPJɬ��G}ED6����\Jev�.;`���<�1����������o�'�y�=���$oT�V�I-~�t0���#��M�@�R�HdJ!&�(�� Ú/���~��/��"_c0�LZv�i:����(J��]d� 0��W9�<>^����ʟc0�j,ts4Ad��9f�w��-�L?0�Ӄ��Bc�?5lz���[U|mee%|�3'~��A�����U���7M��.xŊܭ���:���خ��o�b��>�:�AG�W�r|O��N���S�8o�|�g|�鼡X�ؔ�3Ox#�Q�dTo��@"@>���?�9�{���2�����5��� �$���*)�X-�������a�i�̟χφ�^�t��{M#_w�}+3�\���`���
��m�:,5Sx� ����d��k���Q'�Fߓ��y�Z���&�W���Ń�3�͇_\�<�дz恶6��xE�4-�r�'ƍL��<����x��������ukB �10Z�-��k`.ivp�:N���堙���]e u��!?ϓE|em�V�7��lP��@�_Ӱ$��Y%�9�,+!dd���D��er 6x�*����� px���n���P�ۤ�hFGGG�@��6�Nݡ.��f�&?�!I�ib*�sj�e	O���A4gH��~�[G�Ǣ~m����&��;３6�{!a��9���"�4�����.�{�C���R�������G3m�����c�<��Q�5S߭;��#����տvM�yP�+��7��;8 �����eX6r|�
�*��'4ǵT� �}J�A9���ex�d��B���N¼�W�e�w]w�;�=��!�����:��%��f�dm��.��I��)M�7	�Y)���8��6_����Ì7(|���5T�\��9��$�c���u�1ڈ<�� �|�k����f�Tn2}�������'�����݇�?����n2;����Xk՚F
>T�s������T ��țd���\��(���3e��	�5u��>Ҩ���y�<����<~_8�嶧=���z�����һWj{���+3��i9��?3�/����s���J��]�wu��-Ev��8s�D�Fy���Y]ِR~ps4���Ч���:��x��w;�h7ȩ9��7h�ې�βD:�4i��ȳNq�s��i�6/��8EhΝy���Zt�St�x�R�F���QH�~���z�r�ن4Ȅn���`Ï�`��*�[�pA��O���=����n��$����+>�m��:<ׄ��n%��4e7��J� �/��ik�rs~��pD���VWW���h�~M��خ����a�һ�0��ĵ=�	���]�y��pz�4��n�j?�@ 2c~�</����H���ؠ,�i�6��炫���R%3���_��Se�2�>Mc��n~�2Z��u �~y?}�h�~p�U�Y�@�0D��S��ep�9ፀ���jd��z���)g�)#GA**��jk\��L�[�&��T�� !k�^8	�K/��m�����ַ~����x���^|��3gy���ώ�����Z�l��K�2(r���I/S1.�b����7 �C�Ԕ����*^}�c`���ưȽü���'���Y^�=���K~�Z���X���X��a����W/�F6��I�~����մBSD��	0m���[ͥ���_Mu�i�#�YV�d��l�t0���!����wj��ѧ^�-F��V�Mi��S��hɀ[U�;�3��!���h@�񈮼�<�'}��ܠUg�">%G �#b��e�1C�۵k�-�:�d�R��.�Ƽ�"��v���55�P!���;ٚ"��`���n2� a@����Җ*o��г�}T�?lo0�yZRs�˹X��Ro����|Ќ��f�I?�q@�P�͇�i��~v0>x������������$0��;Ҭ��9�}��M��J��� h������� K������wL�U��x�UZU����?�F��{��3Sj�M���|g��Z(�"#��
�z��4������9 ��Qě� ��'�{�i�mZRJw���0㍅/�+E��d�yj����,��a["�~5h���ܐe��k'���o?�r�u�S;|�j�{s��c_{�����t��d�-nw�]�n�g�x��d��Ζy� 7�7)�Z]��L�D�L�jր��?�B�c�U�d�\�y8�S}^�[�������h	�^��M˱�� ��W�����A�����FiF�(�q�4J%��E��0v��N@H�09��B�3��FT�}귛�l7Ȅ��gϜ@� ml����&y��"��*8CFG�$�[_��αM�1FCEF�gB��Ԍ�#���[����n*%�Ȅ���E�S˨Qe��P�'���{Z���M�vG���VK���J�1����C�����P]w(�� q����M%���:<�&�	�oG�%LJ
F4O�W��
�^{��`�߉AL�YeYu��씤���9�M��.����|���_��nWܢ������Rya|�%�=D���_|L7�.� �I��(.��Ȯ֬K6BK�1']�<H��@
�Y�B��^�כ����uZ��i����Y��q\xAS^M#�N���\��R��T��� Wt��IBa2�I��*���T�y�%�Ϲ������'/��-�(�	@6%�%�f�Jw?ǰ�X�ǹ]���OHG<�#�'����\z���<�⇟�������}�[;��2-��bx����-�� 
ɰm%\+��n�A���JJ熨Σ�.�Z*�\3����-uq�\�W`,A�r,��1][������Q;��,H~�׮��e1I3���e	Lzs1�؝��J�%6˰��;���@�p�$��j�w�]������@<��_�RxF�`;;�h�ĶdwlYT)N��b�os@h���\��1,4�/*�R)�9h[�� �䘆�IY��� 	9h�g>��[��A�(��C o�i�Q ��5�}��C�@���p�@�)tŋ��ad�J,e.p�x��)��J��YLo�T�+XN(��$λj��YD�yD��X���ٺ��8�̣L3�¬y��v���k[�V��'2��x0��/L��� �t���Ku۞�y*D���|�k���J������&J�%aQXg ��T)�>e=�9�@��[��{�<pM�8+*�zf����7�q�c<>�V��Ma�'''a��0iI�v�l>cߧ)��>Ü���锁���I�V�3C�t��_�g-V��_O��c㒡\��z��T�\QYd��tA�n;�׎�M�t����SƗ�i����o�c���O�3����������_��#�p噟.������N��tBJ5����1��sҕBy�������֔��Xo�OHF״乨��((�iֲ��o��y���Kд����-���Ӌ�$~����]a�YZ^IZ_�EDa��i(Jl S��)V��mnm�,��h<����++�f{C��1�E_�7�	?���t��3��>����~�G�z]�KY��(~��.:� -`(n@T����@n���E�1�)I�У,�l�4ဏ.�0��LL�F[qx�5#gA�,E&����u�(�/:� &2E�Eg��0  �[�q:W]L$i(�� �ٯ׉vN�!����L2`�]p�3@�p|���:���{�l�y�s���`L�V�<K�j�U�\�m9;�ޝ�i��ʟeE��ı:<<�޴,��#��:������% �3�cH�R��L��*�d(�&�>W�28TY*������^�<G���˾r��h6o�WvĈ>-u�-��-*yNM��b�|gUٌ&4�#��.E�M�F�j�\��OF(�[Ҭ P��Z& ���n�!�z8��k%R:%V,���5������<6N~uw�^�xg/^����v6��hU��6M�8k�V�����}��#_�����|�g�z�}�����5�HCcƌLޘ��N8s�&M��Ն�.
0ir��3(�x��(󴌧�Ko��������˴��X���X�p����������^���S7��q�1t�"K���<�e ͏n*]|�`�q��uZ���h���c ����N5�CE���T��$9ɜ��:8�N/���{+t|g��WVɵ)?���
*�D�F%����v`�R[��r�HE*��0�YB�C�/��^YH��1lT|�6��].D�]ras���35%�k�߹A�9�)1�����A5�*90aG��"Cg�A�Z���.����#�f$��/��z��Xʌ��fɘ\+�n]�Z�Z=�7���^T$|.M>�-���;�i8��;��T�d�4�凘#`��g."����!׳�c�n�wt	J�q�H�n()A.�}"򙦕g;���"����0���}G��x��<�t���8g0>`�4��7�?0��b�<W��fEU<J���F��H�"�E�C��=��q�E<�]j��Ik�E�i�sv�Y�I\�Ś"��"�cp?�96����y?�}t���z��O��܉��3�/|�����O����ܙ�O.�?��CO���s{�Q����d�r�*}�EA���0�)>H%�� Kͣ��|�m���[4-��xE�4-�r��"��3x�ǩ�`X�8��O�Q|*��6uWZ��*'S�镀 �X�t^��E�:l�w�����nI�VC��A�F��&:��=���n�`Z�{���*�*���v�#�p&HKy�?ԸQDC`A�ᭅF9~���(J"�9��@^O$�|\xm�і�� �)�ndfJ�OB�քǥ��K��A@���Jq��/[Y*%f���Y)^\HBM�un�=P�Ä��1��	E�w]p �vs�3D6�Q�fK�`�ρݴ��%f�ye���N+�u��;���� i�*+)}T�i��RA���v�9��$R�y�^�:J���BgW�He¯�s���eы�N�_�qz����o���$�wo~x?k�ң��4y|����<Wc��xP��� 8	���6�L8P�/T�\���K�&9^�|tC$�E������S�76ߋ.�+���O!_�Q��3��2(�|ո�y�jQ��IA+VJ���;����3�����o=��fwm������KJ�/��_�_���_����ˇ��T5�}��!����M�o�l*f��j�����S�|,�棇o?�����{k�h9^��M˱��@ ��bY�������p�˓��]�6�4�H��X|�uR�q��%(�h���;��=��Q0�v�Fz�M5��P�5T%<�,j2pi�=]�wzqt�.^�&�l�펟ؖ`����!�<]dFJ9�1D�F_��?������&4mG|�逃Hv'|�NL� e��Z��B���(V`BSR�o��Yh�p���Е)�nH��������@��d���p�B��@Y3��v)h�4R�F�T��t��DQE����`S���9Ԭ���6(�����4Wd6>W,��@EaX��0�<��ߖthY�&)&�ps�[�5p��M����Dw����;����`h��_o~��B�q�����_�3��GФ��Ъ��d|��T�XXz)�?	|*yn��j1�^�j����)�&�|c0{�O�[w<���X�lb�nU�����"��I��#@SͰ)���ƙdRh���m;���N̇Z؞M�\�_���k�ߵ����z|������]��m��<�ͧ~�z��7/��,围�#�S�ͮo�4ː�	��$Veu�a�	S��0�����|��ew�+;��i9������«������x�s:��煸�� <'��T�BѾ�sP��R QtF.-��4�D|4�(��=Z��g������=�j��rEΜ���K�84D�Ad}}���V�PBe�M�d��F��:�tr�����*
��a� ��ڒا��/嗣#����n�Rf����V��J�z�-)q��qI��̅��]���Dl���6
�Y�~w��X�d�4��b�� 8'9�׃ќʘj�2r]�u���- /�":/**i�'T�_ Q\�R.1 *��^��T�Γ����D���A�JeΠ�3���?��?�3^������kkk˲��8.&�FA��A������up���D2���ɏ��,�!�*�BYRا���=]��1��5�,
`��)�&56��s�!"���\ǫI6I��RJh����Ű"�Z�!L2��JtS�:�6eE��Uq�A��޳��������_��������o�. ���C����c�3�_����rNZ�	��l(
�)D�p��	�Cc�ek	�;���}��>񶭥�+<��i9�����,\�<��$��?����n�,�ɋ����;Y�AC�A9�^��$��l7�^������I�@���A���C�]�)�.<GJC� �.^�D1�B��u�-�hssS�[�;���ޜ%)�\5,+� �����f���`� N���HK�V�2(��&�L����u�i.��/��A5�XT���r�'��+�d��j�b���!ZW�쵺muV�GO 3аq�k��x�hN�a(]�ݶ"�#�Vҽ��i0$�A[3�����n�B~Up��	�_�@H�(M����rd��+��4�8	*>��z���8��$�~��jUy_=s����'F��d3X�x�E�)�2��1p�J7��*��*R�Ff�v(�xT���@��f��4�)�t�9y���6耟�3H��	��'<OE�<7�K|_��TX��f���R��{��M*t�Zg�p�*]��Ұzm��������'/^~�[_�WO^���'o��kSpȷ�����p?����%���gFV�FM� 9�l�w�L��*�{�y���|�f����-�+>��i9��U������u�g��I��8�?E��(�ݘ|Mx�\��=@E͵x�X�2C��@�w�E��2@��a>ץf�% Iy�-�߼�AG�Ĉ������')�tpp@�=���Ѩ9~�mooQ���R��2@�a30s�#ٵ;�:��P8W��qL���6'K�J��рQCڻ���?����a����C������|$�	]?�*!��A�Eyf���OGGC��Z[�:�#��y@��kz�4j����H*�!)eƊ~E>�����4�Gr��V��i:|.:���s��f�Z%���� B�TD~s�B2\(i�&|0h\��eB� Z��@���փ�����|^�%��??�e�ʵ螃��3�8�b@+	|��AɄ�<M�|����̅�&ZF �|z�3b��2�� �M��,M��P�.���-jw[�1P��}�Ǒ��T���*;�
��ՌJ�wpB�B5>�d���74��TG�Uc�� ��.՜��w��,V��p��{���կ�vӉg����{?u����#�T�5�@�H�a��s߫Q�:��x#�����ԧ��X-���s��?���r��c	��c9^屣��=���o�f�_���Nf����9�t�D�m��#Kee��mY * z��WYu�N���A��{˂���DA�fp�l�x��k�޽��M�n����*�<��E��١[n=� �+ �&��o������_wMr�|��r���ذ-�c�]<tb 5P拲�g�t�� ��2�E'���8���8ēu%�'�3Cy����	�ti�B?�͕������4(�1��ug2x�yuj�=Z�]��ш`�����0�
�|d��i8�ly���x�� �$	�k�T�;���;~%�:4�P�bz��r�3��0�F||�������_�̢c���#�����Fc�P�^��h<9��5��aZ�>C������0=��Bp��R6E�&�\t|2H�b��'T��f���,~/�Є���`� X�u��9& ��ᾈd&Y"��a��_�,��e0֯��Fw'�����~:�t��^x�.�]����ұcd����m��"�k�@�{�\���߁a�� �s���s㥽��w�=��|� +����A������ 5q�	��{=��Ȉ��<N�j��������zu�4-�r��"�0e �%Kk��]�o�$���y�&^�M�44d0�$')����<GW�N��������J?%;  ���h���}Cl���T�QVC		"��FG~^ԧ�]��O��P�&6�V�����j�%��l�R��e��l�;�R��A�FW�Qh!���8�]���)i�x�R���&���ҕח�4p�p��Ez���D�a{mC��
�6g��
��ۮ���BH,��p8Y�:q�ASFSީO��` q��:y���Gϣ��#�����T��c0��J%t�9h���a�l�@)��qQ%�� �b�q�#���L�heI�M���ͥ�p���q𭃃��L�8��z����t��xݿot��@��-���H�����^i��<U
p���V	�) XYtkfvM��Ȧb�aXx�Z�Mݵu'�G#���R����lb���2�� �ϛ��^R�ߣ���=���������uz��st��*��!��.���<��b��-4�t�>��{$dؕ�ZeǨ��KӴ�G1M�J�J��2a�mkJ\5�cNѠ`��7)��)i6���73a>=:��۾r�m;Z�We,A�r,�q,� gѣEU��i��{�v��^�Z���ߡD-���8C���j���� #!�4Ϥ���9�$ت�W�A�Q Y[��e���j-���R��{6�]6��hL��K�^Gu�5k�.� Իs�CQ�F���%@�R�E@���^�σbs��:o�{	���E0c��c�.:�P�A=�)� �<����I5�|��+�5�j�!�>�3��?�4���׻�th4��h��l�G����@���L&�R9�N��u[}����bXS�du+�k\���JsG�e�	��R0����_�v"��E���m���7UeqwV���E��ʨ�z|����V3w�f38IgL3O�Կ6�?y&w�BO5�L�!e7 ؐA0�Ȕx�b.�|'NZx����NS�q`��(ۀt �h2pщZ�uW)��|4�K9�0Tc�00�A�n�&b��P��˿�9/S� ���Fo��4�<�Ag/\��.\��{�)f��ء��MJ�������N��m��Qws�
���F��>N�P2������Bg)�#x<_M^`���Գ��|k���7�v��Z*Ϳjc	��c9~�b��Y�/����q}��͟1Ms��*_�C�t���)��E^JWUU�����6��(����F�	?�N���O�ĐJL@񳵕�8��x�<g`�ƌ���(�������F�VS)^c���@�B���R,���`�ֈ���#��9u�G�䡌�A(�f&�ʘ� 7y*�O��]���b�� ��kh���|T���i V�F���P_��
syG^�`3ӡ��G��N��uR�I Yqp�%�'�1�l�mZi{|Y���OӉ��hJ�e8��\�l�� <|h��c��9��1�+sS8.5�4�aةL�i�ܓ�駂4�P��9m�_�d��/�O�7����;����Yz���|x���y��«���%)�?|��楮t�p�Ea_�q�3�
d+3���*�\|�,F������(���M��}��{�	�{�L̪A�
f<O���̇<���k�!�*D�`>;$~D�V��u�mtۉct��5z��:ؽB���T[ۢFw�ݒ�BY%�KV�vɭui2��t3PGs��Q���P���	h4�8]�z�Yi~�]w����w�}�k���X���X��Xd�3�9`�󍑟>8������C�ev�uW�Lf�{��P�eKW%����U9  Y�:Jx"*�Q � 
�'�-�Pf�������w������0����\?��4�V�%]x 1uޱ�N�Rq��
F�<������aF�y$F�:0Ea�AJ�V���C�Kz�+�:��a�|�բ��*��s�ϳ,b.`R^�s���MI�qr`j��ۑUҐb��s�������fҡ����{B�(����P������69h�� �4�5ڤhcO� e[�l����h����..�ɔ��K�tH"�k��v�v�ZU�[|m��4�`?(��bTΟ?��O]�z��kx�����ٯ�ܬ�?|m�Q���s����sm���K���6�����W��@��D�^�\閔M�$��\'�C�B��>!Y(��M��_9�y� |@ͦ�?���_�)m�:�u
����\x��lV@R�1�A����2Ze�u��t��q��'��c�_��KN�d6{d�Ɓ
��"���[%]�CJ�>O;��q���u
�D2c:�q �hLp "ˠ�6�ɝ'����?yﷵ%��UKд��#��!��?�V�����G"?�� �޶��m�qd��X:ِ��4e�!���>�-R�cPeZ�YC@:��=�(��t$�$2�E1���#)Y�4��c��'���#<����d�fAHG�	5=�n�٢��9�W z�N������I�t9!q�rLW	iF8슃ɘm���[�Zc�g4f��;�=t� �r�0
�LMv�P)�dR
�����S%�O �9ZX^ ��}�_��J�Ǻ�`P6�2:��4�w�c��U�"�;�#���>����9u�z�J�1�T2m*;��Sp��z��)�R�
�Yb�
O�R8.����Ʊk�a�n�|��Uv�����G����(����<
�tu��3�9Zs��k��?��q���ׂ���L�̞�|n�d� �2��p��	�/�ݥ$:���ހ����]���R�u���P��\j(	�"#�k)R|mk��h0��t[<����3�n�f��{�x��*$5t��P6���������7�~=��%z��E�8u��M�SCӂG:�����B�x�7v�t7P��TR�����ɯ[�۩��ߺ��?z�M7-;�^�M˱��� ��8 �ѵC���?7��?ڨ�w׽Z�Ɂ\�=q&���T�vS��;� ��B�w�{� Q"��LSف����Z��F�?�&H�����䝷��������ke���=Ck�6������fh���#�����g�f��B0�+x��<d�.E4���֮�Z�ͯ!��@V-��R |%��!���'�:("C�G��̯)�	񽃙�n�N��$d�J�e�ф�E��eԣ�dJ���qn���I����\������;J��A����1L�`�g�j"S�߱�9�s\�	�* )�9�lT)�-SS�/�g�.:��4�w�4��k��(J>��s��F�׮=�y���L������g��
�r��tj-��{p� ��9_ D�d��"���z#�7��ϫr��0]���t��}W	�5�*��T�|A�B�RS��*��6�	�6t�2�� ���+���siϒ 
�?�s���;ik�OO_�D/����=2�J�1͎ed��L����T)<������6W�����}��y���UKд��(�0pyf<�_֌��4�~.M����Ʀ�o�qGADK@I&�i��- �H�����\e�d��;d��yj��T���~�Z8��
�(��_lQL[#�4P���/��Տo��h��\�.�0j1��ڮyB�8����M�d��6h(MGCJJt�9�y՜�E���2I5g̄���D_����d*�� �D�u�{h��'WHp�S�ҥQs�4\
���8���l��oӯY��V��ui6��n�Lty:���H�єϹ���u�s��E+d 8ȉ5����� �ViIYIegUV,PҔ�'Jy���J�݅����N����*wF�H/�����`�|����#q��r��ˠ���gWF���'<)�`�!~n�(��&���B	�"�j��R%s@B�Ҍ -.ZxVҊ��5E����$��
�2�%�:��Z��1����u�NE�QK�z��Z��\�K@�LJ�Ȃ�jk���cd��Q*j淟X����t��5z����<�9|�9nC�*�=ŋG�{��T�Q}����_��y���x�۾��;-ǫ>��i9��58�K������YX|>��2�� �c�i؞Wh ��l0�E��]1i��(U`@�v][:�?��f��!�&�X�8�{s��.��������
A���[�b�#J�3�>�B�[�D<3
��t��Ur<W��k��[���fr�y�V�M��'S
�B���lj6�g�娸a�����;|Xb8�:#�%ӄ`���$�T6�Tmv�⩷Б������2�m�Z���B�a���D.����U6���t�\SD8��Oa]�.RV���׺(���D�"��I&*��8b.�T_����]�T��.��� 5-�[��aif��B��l;O��se��/j����]���Gt��t�3�}͗���;W��?1��YEZ�ױ�ԅ'�1M�9�&b� ��$34�%$& ��m�x��3 P��KRs��G�C5�VR>b~[J���sB� ������Hl�6Z�C���C_C�Ra����I��#Xs-�MN��1пy�K���h�+���]:8��'��k?�9��ŋuɆ)Ї��yΉaex�����'?�K�YZ��X���X���X��9��}��p�#�O1�y��7�i�u��q�����PaR���Bo	�& �i7� KY��Ȟ@$�B���a;��%���@�Q�4I��t@�}�\Y��v�.���h��e2�CZY۠N�lϤ�ں�:-��i4��`<�ס$���b&��h/�h��8Æ��-�5�pٗ��yb�_(K��7E^�DKV�t��&�ĀXB1D�fåzդ�?�c:<�Vn�-*H��ҡU	��)ZA
���	xK�X\��B��{��f�qn��s�ȧ�ħ���nU��z|g^�eٶ&�P7u�,WʼX��{_��ȓ�|8,N�'/\�{�&o���v�Z$�_=H�ޛ�$��qe�g(Rv��<���wӔi<�Q�M��d�=2x`����� )�Y%¦$��nPJ�$*#\D$� ����eP��E*B����c��*�x �IN���ACMS�w� ������'d6�ا�l,�b����a`v�;�ݽ!'
���I�Ԩ�̾�%]��᱇��箞?�����OkK���X���X���Xt��x��ώ�����Oۖ����oڎ����vВAiM�H��)K%sфp�ա�t"�	�s MuP�<A�F9�-x�)^l*Y��Ex>
�R&|����t�0��X����h4K���� �_Y%�q���z�&
��q;t �(��-R*=�~�9qe�d������F��\4�	*r�)�Y� G�+��7 ��1���%�$�T�).�<«e1���9�Pb!���h&҅<���Y��B�)"R|�c
���n��,]�H�Z�:�`��*W��}���~�u���`-Nc9�B
�ӽ	�<�b��`�Ϗ��e>�����LΜ�0;�╽�l����vk�Z�@�9�^|��8�e��z��,
 � ��\��,yr�X�@���u��3�@�&d��)�1@1�\k5OeIA���<���#\7p�ps��A��ފ|P�|�O�k�l`�G�w[�l)��@��A�#&��������	�&R*^i�h���'u�զ�w��^L/�t����?��`�sO����a����{�`I��<��Y{����m�g3�0 ;I 	\E��It(,G���r��o~��R�ᰬ�� %1`� %�@$ ,��t�t��ךY�/>�����LJ$������[K.f����|���x<�go}���E�#c�{�ߧ�M�?DC�c gaH_>��(Z$�}]��Zv����$�(^�r�	ϩ��:Cn��6���iK� f:�S"���'h����:!0�Z��˕T�'b�� u�A@�pؗ��^o�w���f4>9�����mJݹ�-�B���hm��<� .�*k. [@��?A린�T1�O�8� A-��^n�o�B�JJ���4��#�08�D1�DI�mQ������D�*�$ۖ��p��'���f�o�꼂 ��dj�>�F' ��$A		J��#�5��!J��F�t�D@�q1ME~�@6�R�:PY��P�W:\���Q�s�|��e��3��`Q1|��G���8~���o���`�zc8F$r>�ϼ���h���2;Ӝ��K4�;��A�L\�83�e�mh:'an]��	^^Bi!5]Mp!���IH�d�
u\�3%+@�(�A�x �\~|���N4�����-�e-�'�Mı|:�u�����Z5O`;]��9�YR�;|�"��b>�,mh�ݥ+�}���K�ݤQ��QRced8-�t��\ ��7��M��>����h-1�}kд��C8t��L���ϿMf���a?�
���T��J͈ �ǒ;]E���#�ێHW��ze<�PgR��C��,��T"�dJ	�"l��F����M�@�1zpt�A|���[-򃎀��<�i�4Z��Ɩt��\W�h%�ɷy[�q�FsxM0��d2-	�Ȧ�.���BY�t���xPq���8�$YEyaQ�T�@���Q������Fܥ�YJ_�U�=��#��oPe�{6�n��;g ��ʢ�1��Ќ�[��\�t	���g"�0���?��5�����`{e�Rbl�3L��`C�a8��h����uL���-I��ia�52(R�YjV\O�C^U��</������Ƴ{�������_�s�ŭ~����+��	]y�x���M�Ƥ,��hg� ���6�H3, �Hu
��?8���;``3gP>�&U��@3�,Ҝ�Og0�<B���A���\u�)VanK)��'\�l6��bD�G�Z|^�Crmd&�(�@ȵ�j̳�� �TAM�%Ci�bG�a*�&��\���1��]�P��6���z��]QOΩHk���7$�d�x���>�Sz�UZ���X���X���������8��,�>���'j��vl�)�"x)$岑N2��p�F��3(J-\��0�{B��di��!��RQ-D���VA���d�n0�Ee)]�&�}^���M�A@F�g���� � �+����T���i�u�a���F���dΏ��IN.���Ma�8� �1�A�������Ĉ�%!�IGV��(f$5[,�_�pJ��ik`S��\�ҡ���� ��̋��]B	���K�^��oʀ�b4@��B!��|��5r�_�]uaբ5� ���e��)��;�'��n�6���u�R�jx��	_hK7,�yBG!��q<G��0	>e����N��5��G�X���<~}����>?�����7�hooo�7u��l�k��9��:�b3D�"�_HY�hkW"�橴�)=V�ȹ��S{8���GyK�3��Y��=��*�y�>����`{.9-W �+��%]x�9�.�sszvA:���DF�B$
H����k�
����U�Y�2Sds���KXT��˞��C���BI>r�����u:4�~;��.�޽{tqvB����>��z�����=ƴ�ױM�?�AЂAɗ\�z)��_,�_��_-���c��2]���J�&I��F��DI5�2��R�&ب�u-��*�	����U[uu��Ҕ�"�������+ I���[/�R
�T�Ŝ��]jw<�81�vm � %Ġ�[�l��IPH����-ߥ����xJgSɐA�i�%����r!1Uq��cO�V�^&��V~����EW���X�b`��
��6�S�nT��ܑ� "�'!��snks �`��E�����Xh{ؓ�-��;̚.�X`$�+�3H� �����3���Xּ^s�B�����5E��fp���1`4�]�u��^�!�#�v����=�|l�]�x6�nN���^��æW�G?��l�2��廧���'��$���)�lw��'d��(��{%)27�PFS��4�^�+=%�T��	��BP_@CyҽYAɝ�rlit0���N�*��S\�yJ%�N,�Ђ��d�j�����M�#jG���s��*�]Cu=*�T�g�τ_3E�S$?�E�tNu�E��F	�05���/�ѵ�]�O't��)���c7�~���y�?N�:?(c��c=~D�&�O��E�ڝN��+�&������e�=ϰlh�T����W(����P�X���0`,%8Х?0�@�xi��Tf	�i�e5�q � 0ji]�E��4�۷���$j�e��R	�H%@X!�t��T*�_��'��(�O�1ER�����E�7{��i��o������E�`�P��2���3|��.��lP�G2*��?82!�U��3����H(W�[�(%�h��e���������7	�tҁ��<۵�,-��YڒqK���Ab��O�ov���4\�x���+3t:Z�-���m,[uvY�qb����/Y��4T��]���i5u}����"
�!�M��W>��7�`�o��7G�����������/_D�Ǧi��)EA�'e4dgɂ">G�$_@��H�p��Ob��:)2��nB�g}Hn2���!�D"&ώ�����:O(�A\2�]����o'����耬����o���r5���k1���"�ˆO(,W���w���n=u�e��5je��	Б�����\�D��&��;�޸�l�������>�5hZ���0���z��l���<��$�?^��{�R>�m�r��L��`Ϻ��a*�Fh8�y�H��P��R���2?�$bp��BVi�ㅿM�E�	|d�@�w��'<�v��&R9���%�K�GB�@��� ���.� M����� [ڴZ�/�tZe�3Hs���v�-m�F���)-8��q.�&pSv���ȇE��M.�Y(z�l5�$2
������r(���vJ��kA�<�9M
�J���$�xUR\��֦1��;2�k�5bdF)Nҁ�[|�
M�x��[=jj��d��e؂窱�$opeJK���X�j� ��dᎩL���;�Љ�l8Ou>���`z�w������+6.�� ̮�<:��q\lNc�A@���d��4o�[���TF�]��C��5�/Ǽ�K�F�D��hS��R4�RF��"����ūQz[�6�n���/�4]h� e�Si�(7����oĪG��ie���?�dJ'@wCj���b�҈���f�l���8_ϕ�V��|�����x��_�u��q�5�4�Uc-9�}kд��#<4x�u�4��s:��(�~)N���*�ǚ*�E�]I�Dg T�2<�v������NkI� F�/�L�V���W��/�r�y�yB��;��\� ��I(O-�}j9"�,Y��s���6moMӂ��t�M�A$�#�^�'�������A�C�W	�B�9L� �TuJm�P0�Ei&5jGH� m���R�R�*d-���'���M㉀��nV�$;�$x#HC�@:��	�=�X���gp+��hwO����84�(OBzp��5-���H�Y�9���fc�^�,�	��st�"W`�68��`S�V�V��c�NS�I�7��D6å�g���c��_�$��h���0zf��V�������}��C�!�tjJ9x�譇�w���<A��a$2�)�ʛ��ǭ��Rg�R�@���*�(�$�� T2����xL�(�t6���	�Lu�)�_K¨�y�`@�	�M�n&�Mz҃g��l)U7���e��g�
�U�V�e#�ѥ�Z��Ё�3p� �d0K3����qs�?�'ݏ�O/��+��r{;���kд��c0.���]���ɿ����Ӭ�Y�n?U�N���a�T�b)n��R�h4)W[:Ԇ�L,��Rsr*�9�ܒ8cPRpB�N:t���K&Y.�2U�u�D��ZJ_�`U�
jh�Gpw�Z���;&u��n�֦C�8���f�P��x�9D&Ƣ"�Ds	�%0����o�T!n�����=W۷ɬ��]-m��aQ�7ȪT�f�RT<є9��VrE&��e�������M��Q��Xp@c	�T�^�-�6�b3���Hr:�%d�2x�����L����}�l��X,b
Gcr8��z�@�G ��R��<Mi����
zU�QX)�(��/���%FЮc��=7͓��b��Q�~0_��Z����{���ʕ�ӿL���p�s�>�ŋ��9N�KAC��t� e�̉sH�L��@+�a�.E��05R�T ��"8�L?JJ:�[0��[�.?&DY,����e�|��<�Q���Jɒ6o2�U�m��Z:%���h<�V0����Zi�����wl�:��)�l���LY)�Y���d��U��8�\S�d3܎��'߈�g����o?�/6w������Kvsc��c=~��V�xz}<�~��"�̟���mEM�|'�����Ȉ~!cÀ�g�Cb��p�Z�eǝ�΢��T]r'''�:=%�	Є2ײ$�������0��96VR�hDż �]'hB(�L�0@ɰSQW�������b���90n�i1����H�z�l�'Q!�@և�o��vz���S*�4� J��˴|���V5b��J�x�vuD|(5K�������3�x��(G����2D)Ҁ�9�窬��t��a�@�`}��)���2m��F&����֠��T\(P6ˠ�iS:17P7��5V#��_�9���+x>�%<'�%�h�c��mf�]��i��$������(:���h������_t��yg��;�w�>�x�()��p�{r!��R��B�J��*���Z���F͛��͑K]6�D��5-R�i�^@]�!��S�� ���'�,zcPo�\!���e�D0�Zs����X�Hg�Ѩ���U����|ɯE���b���7APU|
a�S�f̯jT%=[DP�>�l>� ��h�1f añ̓4M���w�q:�g�d���;��u��X���X���T�{���ۣ�>���������Piԛ�c;��2% #����TxF��3�(�\�i��)�2 ��ζ��`	6��h?�w��Q/�I�7T�A�.�M;[;�Zb^2t���� �&�e�����\�Hf!h[����:��ȭ&�2.��]|mK�1����Zh׏���YC^�G��'���	���A��./;��"Z�mU4��'�jP�j!ڣ���u5�
���7�)� ��b�+�Bi�P:�T5<_��|ۡ��m*����<�mA6��N�)�M�,��0"�����G��G ]Ϧ[H.P��2ϚK��䘸�@�:�|	9	Ki`�/[��׺.&XЪ���E<�.���lv����ύ�{������������u������k����$k.E�I��`��o�fbr9���B�-в���
�2=*O���F/�� ��W�x�--nPF�ku��0i�O�|J5<��J>΃~��_& k��4"�4�0K���XJƵ��C9��5�� ���p�pb@�A�~E��@���p٠��xQ�WB�(��k�/�q��\Adtќ��5�n�����~�[O���_���O?�z���5hZ���1<�������t1-���gD|���[m�4�ű�0�����,)nR]��?<!;�W>v�.m�P9!)[���d)�h�D6�R�-�iBP�=�GX.2KJ�Y�n#��}
Ð�ڤ.�Q#��y{Jej]��)IY���/1%� [�� �i����>���|j�\�:}�ˏ(��:�E�A���r�TDx�8���ޑ�\#� ?�D뉤�-��բ��#����� -��Ȁ���n�G�=�rP��Ō�G#�Z0X:c�h��Z�8&�YB��
8�q��q�C1�H��y�H����ө��~�3�%${GHIx���_[��89hɶI� �]���F��w�qx��|�����?���}��e">�?�����?�d~������OIV��7d�\tr0I�W�����H����b��)�l-�LM����h�����mG����Y�.��-M� ����U�Y��!�A�|�%C�$%��c�4h�iB�m�i�U����>�*&
8�K�
q_$<�h�:W5H���]���!]��������nY�>O������gkk�˗/��d񿞱M��AZ��T_8<��N���q�}�/�����u�������R�'P�*�SM�hy����,-���A�	��K�8�2S�6���v���x�plP� ��s= 4��R���Nۗ6sd�~�o����"�Hh��H"� �;�*�J�r���t2a�����z=��ܠ�A��^�AE���j�P���8(BE��}�Y�%@�B�G��g��Φ�iJ��ʷ)��-���cx��6���N8���|�#���..m��4�&�B:<ӄ���հ�a e���>a>�ʘ��L@=����6�o�"%���D�ܛ��5�0��(�V�||��Pd�pl{�@�1a�v1X�r��Z&�a����(2|����_�c_��w��������If^o@Q��8�\@��P�Ķ�̭�G4�4��F�yt��L��Q漵��Q$lp��lA�g��k�� �q _g�A/M�G��Q@�~IvN5�)��ʘ*:ʷB��C4���MJژkS��$ &�?,ǖl�j����nT:U(�ʩG������>��J��cI������h4��x<��ggg_���>_�����M���C�#�sz�Qn��Q�8K����TW]B�Q�%x{)���2�J��(�"�WW�RNhZv�!\����u��v���\U�"�)\����*l���$�e���8����3��a����	��p�,�PQV0��`�T�4�ہ�b���`���G4�ЌIZ��m4�G4cz��ou۴�oӠ����ÊE�)[D���}�Y8LX��Zʌ�j�1Ed"ޟ�����g��%M��IFֆˁ|@�oJd^��^�DJs��`�E;��HLg:��A�xJ ��a��%�	��R��Y�6#Ǥ��f��hQ��g.`	/�<7-��@)�T�<������y^ �)�As����x1�|���.ϫ/�x�/�~�<5��a�6�a���(��\J� ��˵��`�F)�c��.u) Q�ƺf	,H������Ju����^*D��CG�����ł:pd4UIy��b�Q��ejTyP|���F�H�O��d�F��d<j�Dƪ��l�xmC	�6�R�@��ƪ�Nm�IK#glL%|-�	��5?M��C�/76 �=��۷������wv6~����Ϸםv��c��c=��{M$=�����i6�7y�������U�apV�2�@'��N��Ɲ/Jn|�Q�J�U�� ��X;�Z�u!l�3KJ�Ȕ.. �RL�3)w�j2������=�� h��>��L�@g<��%
Z�MN���N2͕
z%�0�E�I�*3)����b�Ԏ��(�)ͦc�� C���i0� �ף�l�D6y�J*cb����/Y�&��8�i6O���X�A I���3���d��Od ��An�1�S8C���|˥�ݭ=�9���>_�<Mi� ������Jg"�V��A!���,�u0h`P��r|�}(��J"��(cVj����nT��	�:����m�q�(�J�6��̦�ܾ}�>�����G?���߾�����G���jS'�q�1��%���h)C�KY�e����B�6,���@Cuƒ�dHV	���b!Ә��d� ��|�����7 Ȟ1X׈lw�[P����+J���|֍Z�VF��\'�e����'Y#�PUi�����/�v��R��"�
�aK�#C���K�o�Ѻh����,�]O#�,�p]����#i��w��>tvv��^�ֿx������c��c=��?9�ό/�_;���`켨��k�llU�h�_�2��X(���@��n����K;;�Z��Qdld��G�M	I�Jq��@S��jz�3A˥�x��>]�h�Ӷ� ʍ"��c�AY��kd�@�ɰi+��s���d�-��%�?��Z9(�p����|��d6��3�����mQ�ߑ�a��= xǡ�h0`���d�`n� �mϡ>2?�I[�=^N�`�I ض���"��<wx_{�}���bJ�"�0.(��Sr�.������E�vEY{4;�R��xDQJv���_�T�,;8N��"�eE���]�����C�l�is���!Dd��My?F��1{�\ɖlm��iL���W���U^�~��O�;�h�V��������<^�.S�`T�+�X� ˃� ������j����C�F'yS�JW	���U+%Fʯ�<��X��&T�v�Gg�\��!x3j�%2GK,�l�j�ӂ�z���d5�Mt%�6��<K����8���|U�DJvˬ���jl3:.M%�������Zʀ�>��˗j�u&�^���v��L��[��}������ܹ�|>�y���3Z���X���X���OxgD�qD�gޟ�'ʢ���8RV)�AըV�%��Hy��\:�p��ؤ��-�j����@�-�Y��L�(a@�Q|�j������m�*�f��¤h�� W �wdFP����N%J��b�TU])��M�v����4e��o Z4�2b�%]f�61�g%�sGd1�@F���tL'����X�a+`�(͞ǯ^��A_��3(�Vx�R��F��${Q+���Z�7;=�v�ÅhR����f�K�f�����е�C����AԜ�� .���q�P��ڿ���b~��s�������S���	A ϭ�Χ��1y�!u�qKL$������_6N_�x�+/��+'�� �}���ۖrd&�����2���ڐl"2�Z6[ ɒ?$����0������J�ےҚ"��ݏ�Ԓ�:��o3(K��'��|����k�8:�)�&�T�1�l�ТTfI��:�d�:��5Ow!����g
-=�ձ�ֈ0�e=�V��"����EG���Q�e) ɀ͏��*1��䷈29�Yd����Ͽ/���~vss��ݻ��+W����N��c��c=��{�Z-�vGa��$.?V��3e^=ZT��8l��Y�?V���h�O�X �t�9���v� ZK|q�n�#$�q��=�y(dlC�i
�s�¯5�������A����@`��-b$*��d1��� ,��Ȓd)߀3�#�E�F��� "����ox4�U�n�A�M�G�h�����9��k�zM�6���A�A^z�>-�/^�<Τ��(��%��6���{;��lڼ��iL���W��B�����b0mLS��^�:AK�Y��tN�鉐��%�Pu�E��nѣW�(a�9[��](a� �a#Fz�R���i`���)��EJ^���T��{%X�v�6i>��I8����п�5����O����%��U���x�:�L	F��Z�vV�(8�u�APʥ���@�Y�D3���P��f��/
K�آT�Q�,N�t1�P5�Q���]t�A��>��k����\*Y��&�Ç:h$�ʐ2^CKG����<2T�������bOy7֔h�p�{(�Z�2Y�4T�T���>?�Tj�dg3�0�ߊ�;�v�H?q~~���d�G�������/驧��z��c��c=�c5�"��� I��E��,-~1-ʷ�Y�o8��paԺ�9�f�ܠI��&ߓ��h$Y ��?�t�P��p���*h0!�Uj۴���|����ї�:t�� W8'�,�O�MЊb��,Ռ"��p�)^v��~]����W���]�ǀ�Fօ�?�S����4�ɲZ����������������� �5���� ��t��#�i��g@6<%r׏_M�*S�Z��R�,Y;��1o�!m���C��b�QI�!�ȯ{��[B�>�y�f�NFs:]PeB6a �B��]2�l�;]�JJ�x�f��Eq(v5Ý���&��?J�a���Ǣ����]���sxܜ_����������Z��O��7�49�ʙ](t��a��߸J$�2��@ �RpzD5[����@0ţ�� $��6/�F8��TNs�Č��	��� 2�\���=>6 ��d�?�%����� A��XJ@�qh�^¿�Uk���V�.�%i�J�]�𦤬����/���u� 4i)� <?�,�+`9�ضZ�y��:��Q�@�d%�2 �{�7�w�0���7��x<�%����W�����?��ۻ����M��!%8��Q�$)������"�ҞR�E>��F	�XZ���e8P���r7@߽����Ζ��#���IДvi�kr6�� K fK����z2$��k���"/� Ä��Ԙ�G M���6mmnӝ{���+���ɉ,����q��PQ���4`�TE�.��踸K�����}�"�iI�a[�k��*S�p�/�"�P��61P;�mM+��WN�j�#���T6t�@�_\��n���yх�nC̍�XȔ$�E+��'H�ؾJwQ�VC�.k�0H�yy��,�))�\��8�m�$s�@��׏��V'�h�'�?�_�lGt�@�����ω̿�4���"�ʧ�y���'>�������ѿ��O�;?��Y3�B&�B��Z��D$�$1�c\�!���貗|�P{��F�e���E-F;ci1:��t ���������LtC�;r�F��A%)Y'%!�rT�D8G�J�/j�[Q2�-��wF�0��Rۼ,�=�a\z8*�C󢖬&�2E�I�.빚#�,[��|ڮ)�7ۊs`e�RI���h�8O)D���Z�c�Ԛ�m��w����7�x�|���\�z��G�B��c��c=~�G�X�[�,{���dy�ɬ�����q}v]_GR�0�
�Ԗi/9���{�bPs�� ���S����ّ��C�g���f9 / ����Zݱ���l������^]+� @�P�;Cy�"<��L8>�N��x�:�]����Э;oD�/]}T��r�7��2���4r`��ѕ���k����dJq4�[�"1A�C�n�����T�e4��z�)%� ��9q.ī����������M�d �i�x�=�r�K��E3:��ͧm�T�ʣϵ=��>~��I02e��%�&Uf�����C;��^�wLc��ZY|8*� W� (�/��R�T^i ;������LQ1������f�)bO<�������������Ջ����?6�.�����V1x,�X�jڼ�$mW�dBc�1E=[i �R�C֤!e�[k)dZ����}p���gg�m����oS/��gss �L�4�]P��F�nJY��)pQ+=��^uY
t�2�<F�t�z4��>K�"��R�{��<�U,+]��r�Js�Y.F2]��DK�eR��F� ���ﲆO �m������}C&TJ;��c
�_�)뗼�W�l+�'�s{��_9>>��}�ʕ��c5֠i=���lh��i�;������y^�����u]Kﴺ���]��� �,�Uf(-r��w@���N��t*޽�=�� ��
�Q*� W�⿗d�f��Mゎ�R�ۗ,��A��$���;����LXO�Q�@�b<'�A��+�Rg�կ}����i2�����47���KY���K�	ݼyH�A�.����Ɛ*���"B���%�n��h.当�3j�;v6y]u;]�B�R�t�y��6 �7�Y��Ԅ�� �Z����B���-������v��I"Jf#�|
'3��9�|O<�(�8�2���?����^+�qױ�C���,��0��C���(I�Bm}�ߢr�����)%��w-M*�z]��N���r��eV�	��tͲ4��9�����u������-˼� ��71��s��-�.��mm�R]e4ŢG�N��A)r㳅 �>��Y����)Ut�,� =ؤ�z�p���S4�����'1���ލ�4M%n)�ָG�YӎDn@q�D��PM�����)`T�*��:�����J礥�p�`�T���VA�֜/��U�)R{�*~�ڟF�ʺ�P�V�̓��st�j?E���f���l6�����~�5Z��X���X���T'�0)����'˦��<ϟ� �[����@M����k��(��Sy/is��$8�� V���� ?�Zr�DVf�{MG�"O$@�Z*j%M�����V�r C*Ӱ&�=��I�S��QRD�]c���E/��:�|�6ݽw��T���\Э��ʵk����G~Х��-�3�s��iH׮^�aw��jJ|�-
�W"u1�08Ki|1�����u7z4��S����*x�"	> v}�|��Ŕ.�܎C��Q� k>̈́7x��ۢ�~��[�(ة)'OǴ�C)u"0��qG�l1�@)�;��FqiJU:���h�2��S�6&%�F���"1?�8>�Hda�<�-��	���J�CL�.ZD����͈Jz���/�����x��oy��W>-�K�je�`�8l�ÐLݽ�Y��C��w��`.����JQ@�%p��u�3^V&��dN�c^@������R����(�{�g���m�E�E"�H��E�@!7R�o�|�ꖓ�{��tYn�^��=)�iФ�ג�-�#T��<�c�7��K#�K5=l$��A��`��'>�_�t��4� �i�� �z�����j�����m�����`�o��Bk��c��c=~�����YZ>]��O�e�3M]��2����V�����@	C�4�%��;�s	#t�moo+{���2 ��})�aT�C ��UFc���?Bs��I�9�!seh�@�2Vw�(����Q� &�4��l,m�A�O=��v�n�;�4�i��M�4./�A�ɺ����ms��nH�#�Ft��}2����9A�u<��ڦ��!���#�N�i��t����<�=<):S�9Ǫ����az丁��' ������8��ӳoy��vv���"��&���X$��~����[|%��W2O�~�v�����Z��;o�k�ߢ+���7��V�a�PXe�Pb��H��	X"�f�IJ'�g��ܤK��ҡ� �e{4�F�W���G���k�|����`L�C�,G�W@�ֶ�30F��!
��ʤE���}�O8U��)� �:�� ��sS񱘈�2�ܖ�&K���EE�����)��9�ZyJqN���ry�SRzJ��
T���c�s��PJl.�KJ<�X�$�,=�[��h�����6�qLd�%�����P-Dyk%�i�ˑA*q�$�Ehj�:��4*ɍ��$�
Uj��Iʞ8�x�{��;���5hZ���|�sӔ��I��*����٦���h�E�T|K�hS}#��'Zh���Lf�nw�ҥ�j�a8g������޾�mP��0�m*%܈� �t�i�7Z���Z�`"�##��(�k�o�l�@�g�| M��6��.��J���������{@�i"�dh���b���{{gG��x@�F&)���_0��J� T�om�iw�2���%��5��4]:�)�����}��gGdy>=��3��SOR;���|�R��}H��:��tNaV�9p^���e0�h4Lx����w6ɫڢ�=�i�e�)�6��@��4�2W����[��ֆ�ᨬj�\q��4��/Dgj�צ.��JE ���4hݷ�X��2F�J��,�`��<��hN�`� ����v�|�����<��>�u&�H�4e!`�@�!�d@�xb��ve8v�y��D�@��o�.�JR-��Er8��|���bXߌ.�CDiSʈ��\&rހ���ڍ"f�[mQo���2M��L�Y{(�I+[CK2-��K� �0h�_�xQ
�[+%V5+2y��'�0���O�<�p%��g�`&2ê0��o�" 
��*��:��,�Sz�M�m�̶��B�O��>��AJE�׃֠i=��Gjh�Rk��7�Y�<+>YT�;�"�)�]沼`�];�%;Q��dHj	2]�z] .�GGG�uAyhwwWu�Y����\|�N��fE.�\���Z^KT�і_خj}��]�+�H������J%\��Ca;��*M�e�sߵ��[������ |��W�)�;e�-�/��M�iɭ��UF��ǂFt6�h<9c0ԦA�-v�d��]��.��֞d-F�s�^��@�[���E�i��?ා��/�D_�uz����]�>K7�N3������&�}��9�x��M��6v�������F�D���ag r��Ѡ�M������	�����S�� O�TU@8ViQ˜�k������w=CW.�r Y<�5#2*�O��%��i�"�	�X�돿��ؐm��C#d(��YIM��rq�Y��Ǫ���� ������varG��a�U$��w�����M*+ShEIK1�	�^>:[�A�l,�"&�w���*^n �w�XdP,j����d�@�0M�7�}��\y*.��0����ѭ�S�n�jP�&+�|��\=M��~Q`H_��N��2�8w!GU��xJ6g�V�g��"�լ���玲�����+ ����q&Zy:��9�~S;��kд��#2���Z���>Z����]�iʪ��J��;MC�j� lP�XZ��{�O;��4���޽{©���5�J�j�
�ԢS	��J_�C$C%1�*aG�oK�@�|I#�Z�@�(�*S��fs����/������������[�^���3�/�}��[Ee��05`+�Lo��c�^����SC�ݦ�����Kc)7���@q�Ӣ0�I�v�ƍG���78��)�G&[b����;���v�św��n��߾C��\=y��q倮��
8���n@��%��˛���|:���5��K�W)0�?�@$LT	
Z?(�L�v:����h2%�?I��/��1Z,�1�C������������m�J���UY	�8D|���ƹdk��� &[�����B���>9;g0�(����Mϖ�#1ܜ��?x7�[�?�)�'���w�m�=BI��c>u�RzqBn�'s������|�ng���ߡ��8�<g��Tۑq�6@��lJU�"M��e(^OA�HV	��DY����&R �T�f�F4���|'S���]RUg^�Y��u$m<�U�G��0ߦ��Л����4�[55��O
�J�A�˙Z�
LA�R�� A%4��\��N��e��J��C8�DYJ�x����;�4��z��l�(9���U�?ǁ�)�l!�(m�|1��A%�8������tFA�-U�>�c76(�z��4,�tv��5��R AǪ"6 ����,"�����uby(M��JHe�\K�eۉV.��dWH�et��Ѽ�׏�������������y{��ml����8�Eѻ��c��q5g O�\�N��� h2Wv$U�
��}x���L�����I"��U��g�y��^�D��\.�<���s��zt����Kn������c���})e~�k��F�MO0�zǳo����L�9^݂�
�����!����-�YE�Oj�KC�� ��	r���),,*���z�!��&��1�{"ƽR.��(�%E���5��'��[��H�Q�E����tO�k���H���\���Kbɂ��Q�1�����b��V�&-�����X����6�C������+d�~�|\����	/�JR����fz��`���P�;���1ų	�"1P*�t�$�t���.�%j�]Y��@M�t�MpO-�%f�� �eYNI���)S-uUL3�s� �!'����.3Q���w�t��k
8���E~+���ZDJJ|zY��C[>��U�.�C�.+�
4�T��#̛5��]}���7����?�����M�?�@)&������q�eQ�/�7˱M�6$�	�Ȣ$��������5a\0��i���<2I����K�"=ׯ^�I�Ӓ@�Í^�T[{G*���x���Z-(=+P���MQ�W�j-Xʃ�bԝ|�.�p>�����N����^�3W���𶆆��[���>�b��apv6�/�k�I��y����gn�hS-H:וm(�y��LA�FKt�
��jd<
U�ʒ��Y!��}�t����=�N!��Ŕ?3���ѣ���p���\Ы���K/�B����X`p�����;򝚼*(h
5C_�Xϩi5��\X<:CV�fDC�ݒV�ۧS:<�0�h���Snk�ܠ$�^�!M)G4�b"��%f%j�5/��fdUl^�������<�)f��j�i����i�1Vv4�h!�)����D�*Q)�����?&�������_�L�����c	�8&�ш�](!'�,q��@��o	��AS��9���	��k,x��^��F��K�5��*�S�m[�4�e/ Sվ4����2�54q�)eq :��hK���]q��R�m�C]'M|o����;z(V�h �z��g�ȘQ�=�����Wz�4	�b8�����w�5hZ���!(��E�$#���y���2�4�}�7=�V����Vk�>jG	�IJ.�\�`{p&�yD/���9P��|�����=y����� 8�۔��)"/��.�@�,P`0Rw��,�T�ZҀ�O�����f�I���7�������<�v�ҥ�/37O��)_m����s�n�a�3iQ>W��yݗ�� �]��OE�ρ����L]+�_���@���;(U&4������OD��O���|�q::>���#�9yA�.ic�GW����|���?�����v����.��إ�]3p����5	���!W O�b��{TC�!WV#��a�T����Ӄ�1�;qf`f*�Q�Xb�m��|�s����� ��C�c23��"���-�R8�7^� e�Jt�x�	��������"��"a�T(˜��Q���T���פ�@���&�;;�>M�N��%���X�q(�����9'���KU�0�И�ʪ��@�ȃ��� IcC-�O��=�.9C�LE��"9��YZ��lM�6�#�$�h�nU�,�J��r�$.�5�	XZ�P������UU:��������K��2�	3���U/}���h���ZL� D4M͟������T/=������׋�v�EZ��kд��C0,������_L��|�{�i:��6C7K�FHԨ�[TU�P�K8h�w!;��C��
����{|�~.�ɏ߸!\&d�p���7���r!p(a��mskK��L�p����mX�a-��D2�Ix���ȑI�r���<��X�r�w��o}���{d��R�9��F��899yi��N�O������s�z*��P�pW��� �I�RjMFw����;���헾�5z���裏��m����g��tz��s��y�[���-��'���:&e��8�E��{#zp��l�M��xB�̀[2�JJ��t���)�qB3+�g����lJ��!���vO�B��L� P.Ϋ���̍��<�Ɍ�n��D��s���q(�����(\�bs�.��0d+J��Z��sNt~~N:�e�b	R����@>�Sv8�~�a�s7b�)�,T�z�yХXe� -GD�R*��,�}�D��Bi�!�yh7c*�$�TE9K �)2 ���l������[%Ė��2
̐�Tٟ�����7�����]y�4�h	zޔ2i)M`�J� ɲ��"�+5�FI ��M�����J�A��N	xB�]֥E/�:M������^�wD��]c��c=~@_��(���ҷ�O��;׏���	�e���=��OQ�V6���LYT(o��]�|�v66�<�wH��ߧi������Xٝ���7:�@�Ev
��w\jw:��iJ�,�L'��d��m���T	+�7HE��y��ir����u���}�`��ׯ��s���{{{~���y�w��E1�gYY�-J��0z��^QT~U��0������.��(�"�����Q�L��y�&Ә6��t�����;w��k3���'{@�����碷�@g	���Ǫ3�0*�_I�Ѷ\��2��m�A�%d�2�RCi�o��q�">��~@����9�����q����&]�&b����ȳ�D��^ۧ)3!�;>��lR�L�t�5��iy���%�D�>��mupWtz~�.����ʊ�X�|�m���|MF��|<��g��.bj1�3x� ���� S���3����X�m�*�IK D�CN�F�R7��&6*X�k:�d*`�2P��Y퐩�������+N��̇\&�)U
8�T���[>4fZ�Z�2V��Ւ(nh.���X5M(B{%��ekř�A�i���z�9���e���k>Ư2`����Ƃ���4��z��� ;RfQ�</?������d���ҙR�& 6�Q�)xJ��0z(��#h,����ݾu��޽+ZJ�N��y��eB0�8��Ñ��kf��h��� F�M�g�t+Lh�ƽ �+ۆR��vP&,H�I�& ��qKz����uۿݿ��ŧwv���yխ�H����8��l��-7�g�������x�Y�]ե��S�����4�$��ymɞa�5:;�(ߦ��]z���"�y~vʟ��B s��I��<�yBM��	d��%��g��?:�y8�;��4m:���z乖O P� \��AݞOO>���t���'3�Y 3��x��=�6z6��Y@�r�ز���p�L�t���$u0v̊�]٧-�^�U�|4��w�2�󩷵ǯ1д4�b;��R1~	��agH�ǔ�@����<H l�����y]C2@�>����L�*(�#ŋ	�"�*6,]TǗ�"5���Y�	ZR����Zi�`�ʢg�}��)�c���,ս��Z�nh%p��j�߫�ऩ��V�.aX5Ɗ{�VU?�$-��d��&���Y)Ry�&QJKn|���C'd���^�-�%I����_�t:�ZZ~�M�? K���$�H�V�V���86�9��QA��p��Ѥ֔v�w�P��m$�8B�zc{K�	IR�k�ޣ��I�h��������C�a�@i)! 0��u�&�%.��
�e�jCȦ�pL[9�M�|���L���[O�
���wf��g[������}鱃�㿍��~����s������~g�&�K��eU}�"s�����ײ���d�0o O��`c4���@�i�;�����:�t��lSN(	U�&L���xdT�t4[М��-5�MAG�3��S�����6��q��B��g`���r7ڻ�G�߸F�E�`w.%�����Aۓ�T<=a \P'����G�_��4�H-`��K�#o�"�8�2h2]� @���v�30c ���Kվ���~��%������_��K����W��	&���$���^�o�Df �s
\8�r�<�tb2�i��V���P��.��I��Qm���3R檵�0��,�"�k��1�%��-����gjr�)����)+�y��|�{
/��1�Y����L����3�k��(t�z:��<�\(�K�ْ�v	�0ޜ�#Zv�*ҺL��nM�����,�_0֠i=��oq4�y�c,�`�zO�U����M��u�~�� �!���%�Ɋk`F�����ם�=	��b���1����6xGמxD���]���h�Z8I $�(��}!��"MK��r��lh��4:�JOF�N��0���E<�����4{�/�������p��k׶�yY����/�O�p�����b�{�8|fL��\�ʻv��K��!�h#�Se�k�ՕC��->qw��la�?v��PHң������R�M�4j��K�ܼw�^:�O��ct�t2�}ڤ!��C��/^�ݍ��x�v������ZR��M|ܪ�.�W�(D��I�dU	�?�ݮ��֢�kS����1HC˾����6d�c����E������Oi�Q�$��� ���~����x�Э����F s##��g2�D��n�hE�xPGw(@�F�2�KIK���Q@¥ g�%��J�T�q�b�	8[�,��}��d�j�b��W��*�d>�@��W��! Q���y�$w��C�M�=bՕ��X+�&)Ñ.c6�.e�n:Sk-i&�Bt�ꚃ���Kam]�]����l���W����@$�x+�qx��΅_��Ϻ=�Onݺ��}���=֠i=��oa�m�����eE��u]=m�n��AP�����)e���`$�n%��nJ���41��bN|�b.�ؐ�|���,]W[�t�!K��~���o ,�%܄��q�E�_I���+��҆A�)K�&�a8���E۰?�����-��#�<���0T��	||�8�RoM�fi�EY}$/�g�޲˕�
aA���;pc��<��;�"�9=>>����v���{�����wНh�)����SF|\�пj(�K
����lS�͏�&�|Ҝ2 ���{T�?��J����
�� �����v�����^b�}r*��*`Д0()��=)<7xm{�I��7t�ԠA�K�(U׼�M�o�&�]�p�rp� "Z�d�B]B&�K�T�4�LQS�M%zS��+�a"\��#���m�$ :�p��`��,����(�n)���ܲ�O-;�V�p�k�U��JS�=�����a�U2�\�Z�c	��`�P
�KIR.t��7/S�ҷ���'�]%�m�W���A+�ehF�����0`/�d)��m9/�ւ�%X���oY�N:C��+U���.c�N��}0����1�y<����֟����:9�?�c��c=��~p���,��}>��Oږ��8v�i8�ėZ�?� eOB"Ĉ�Qw�ˇ����GE�Xh�`�Ν;��@�C���!]HI�[^��6E�΄/�g�# d<O����0%XaP
�JR�ڈ�(.9M��)��&˒���7�.�S�n���ݍWߡ�?C�aO�8l���Q�o�,oVc��uU_�*ӫ9z���c��,.�ޛ�6-�##t��5~ޢ��c��#r:�65��E�vh�צE�0��(��(a`z�2Z4�G�6�ҰO��/&��)�1	��^O�'�(d8�A��
L�S>.�6�\ؕ@$˦��)dPj�Pv��ܢ��6Og�&�����]~���@2F�^w@;�5�n��a"v�B}��{C����Φ�5A����J��U��/�M�dɞx��IUF��T
�  �R~#%<�˒�t�YƊn�┥_pP�[fP�t��-0)9�Ze}T��P��z�0�U�V��<��\f�c	�H�%�'e鲟��Q��G!����`Q�蠊.�»�E�a� |��9��f�CY����J��BVM���K �/,|p\+��R}=K�xvt��h:�������}x�P�?�c��c=�`i�eW�q�q����;��u�/���b��G�I��
��c%��r#G�Y�V���V�x4����,Ố X����}�U>� �1(��:
��pq���L�8�=AZ��R%��4�UY���R�X��*���ο	����׽�����0ߩ^1$W^幼}~����,�^$�GҼ�9>�O�U#�2˖s'Xyx<_��x��w{G��F����
3&�ա��z���9Ⱥt�lB��B��t�Β)m�-��ե�����,;����Uϛ�~L��� � ��\qAi�؍U�ǆB
��P�~J?���J���K'h`	C; ̸���i�^?_�n]��2ϹU�u	B 8Ө�Q�^ի�u��9y�������< ���>� I,�R�1-�Yqc�Dr�����}��j�>�ha�`)�4���.ωƔ�ѐ��F�E��"�C�tӉS���yt���Zh�\�^o*��΄��M6�0�)u��e���T�:���#��l���{�c�zSݰ��.�$�q( pݢ�͒���^pڠ�'-XR��Mz��*[�������;�p�_L�|�"��X-�C������P�_O_xj��T�"���b~٠�$y��L�,��:$'Xr �p�z��@����*J*�(���5�|�w�D�����ht�ƍ�������k�>v�z��h����>�8��?�D?��?�f�O���2
/7p�jH���"P���p0�F��1��Py^YX>���7�Нۛ�7Fzii���V��n��ض%`���a4�-S	W��3Ў���X��x����W]Օ�L��h��F�ǗƼ�1��u�<}�=��^l6��g�zЪo��m�w�������㽻?��h8~�w�S��W2'���#"0����ں ���]�}kC@���"�[st{w�ڽ����ש���tz�^�v���G��b�_յ�o.�( �H҃��9�ሿ�|DA�L�jE�����t$���t�z��OՒG�|�+�&1z'�����|��&�8���Ҭ��hQ2Ӡ;d���y?�t+��l�P�G�馔A�g�6y�l�&o���3��c~>�R"�@�h6z���(3�k�^���k��AmS�j�8�!���V�[��Z�5�|]��[ �"�sd�RNU�^��E�.+*��I>�qrT�I��r�d��BXR�)K�M�S�G�D�#'`�	rm�$���GC�e���� �п�^�_oq���� FD�EG���Fa�b���J�E^��?�~G�����|�����3_Y__�u~HSv3�4��=l<�6Q���3�x6
�?�z�s���,����(����D6�$3D�H4����f����Ҋ94��ظ-������IV��9��9C��J ��3X�
��[t��Z�@BZd Ug~O�[�\%�/���8�%U'�y�	i�AR����P���j��bsn���5z���Y�^��~d��|�R)?���{�$}2��'�4?�l�T��^�+��yـѴ���J���3gh��O[�{4��m�ܢ�4ߨӍ�z���hgwWJ�窲�D����j5*A�Tcp��
��T=:���=dD1�nӁ+b�ؤ�nFs%�:�N�;C�N��hD%Υ,)�N�GWoܥ�7�js��0��N�H�DA�)N9o�

\�.����`F%����G�n�P"��y��{HO��T��*3h�S̷�S�
F�[���[|	b�F��r�&Um�����rI M �c���2 �2�S�  ��IDAT�61�5�H(�6���Q47�E�A����@��i�-��|r�BMS ������Ka��Zͧi?��3���"N��PEIoBB��x$��Z��lɑ��}�)GT�A �:�/��p��T_��U)�}$���?��u��N��ѝ��o�g{����c�@�l���`��I?����s*�%�;�"����Ɇ��fc���Ӣ�D��x��eqqY�J�1:&�����v��E�<iu�'%�RN*�p̅�yi[��o>eW�� ����j)���JUIǁ�$=���ABgO4�Ǯ�.��V���f�������[=���v��a��Y;\�t��Ϗ��^��.󆸎�Yf*�L�?1P%ˋԨ5D�`g�CI�Z�F�s�i�n��K�|�^[*Ӑ2��M
�s�����(����7"���^e`>�erk��yԫ5
ynlm�ҝ�;4��o��S�t��9:ub��5�3��2:HU��0b��[��� a�n�9� 02�������$C
�|i�25�� |���HáʫnXI���ѐ�"�l Q� ��Ӧ��mp+��L9H�I׹F^ "���Ij��c(�ɤjM��m�"1�-���qJm5M�3��3��6��Zv/�|�r5�E*�)��i���`��RVD�\m�kJRP�$��;F����1�T�q��P��se�Y矁��/8�oPYt;��ߗHe�^��/Z	1�B���_�ć�q�?ܽ}󱃽����/~��G��a�����٘��b���4�q|���3���8����؀�\��2[Qx� $��*a���DAR���x��&,,I?8�
Y�3Pڤ�w6%冈�@�k 1c��h=�V@�T˝9sF��liO84]���I�7D�@<���J���1���|����q4�ǣ��6��_h��Z���?�<pfeɖ8��΀�˛��U���]
.���|��N��<e^�gF��`�z]%��T8εFt��6��})���t�v�FnB��K�2�ڃ9�����n�r>fka��\��v���W=`@�	���l�:|:�v�I��.���٥�ׯ��ez��y:�4�*�L�t��:mm��5����!K��$���clHLt$v�5����P樤��Am��Z�	�;�5�T�U���)r�X�ؒ�R`&�)I��F'��d�P�+i<�_�$���^����d&��Jے<�\#���$�=�B�T>���gSq
�rIIZo�p�|#y���+j��K5�gR�r#� �)I�=y�F��^�F!"NU���)_CV�(A\�7�nȁ,�5E�m��j��/���� ;e��V#�\.��|f��?�=���^o���n��4ϩ���>�<M�1��@��ض�§����I�#ͳ���&8 ���褩�q�e���.!���0H��)�\|nN�.�:�q"���b���)c_YZ���ia" ,���le�,1�D �@�V�n̆U50|8lؔ�@7*��'ܪ82b���mk����+A�������ZǗ_}+U����������F�����?7���F���q��+M��$͂f�7;T;�GTc���@�-�s�.ݾ�I�.���.g��SwM$MY��G1ϵ�~H�x���l�7�j�'Q�F	@t8���F�Q�z���'�``� �d^�Ji�L��<�;4��Q��֍�i��u�[��y�����I��+�ߦ[��?d��|�$y�i�x�%�a�#���-2!���c���0l�;@���Fe�Fo\���r@I������ #��Eh��<*�䄯d��4��4
�H4�'�֥�= ��L�+K
���L�pl [����H�':i���r��dU�S[�GJ�N�P����Ǥ����H�U�.Z�@���ߑw��=9��xn r��F��
�����$:��K���Pbp�4*r�.�LH����,������6��b)L�s�'ůW	�s��
V���v{��n������?|��W�����4��l�=�a�m��N�Dӻ�<{*K���4]�\��чA�ީp���0�
�0�wmW�K?��ǎ��*���/`���qN�>�`��= #Tb�� K�d,�&��ɥ�5�@fe�K��(Jk\��p�
^�s0�H�y��%~/M�/V*���>s|�t����q~8	���8�8(W|���W�;�?��OD���a��#K���97q �Ftwk�j�����&X�ׯ^���'���i�A�-�h���s����^�C��X���n�*�!�,�xC�ȥS�.�J�D���F�,|HE �2D�:Ҫ��7�,� ����I��wQ1�����mz���頟Pꖩ>7OK�+�m�>�3��=O�T����� \H��#�
�#(���=�A@�v5N��x��m:��/ q�F2�u���h��DHؒ����4I�4UG�' 	 �����+3=�r��d��-���39��af�JP/�?��R�1���J"H�MoZݧLw���d���F���7��k_�P���H��R���`�|�%��#q� �U@�^� M�L'��;�߄j^Ñ�b���;i������e�O�t:������/<���h���82LD���ג~���~����>g�Y6K-7���Tr}x���|T�i~*)��%�r��f���@�+�m/���!����.�"��#=������+ؤYD��--�X�T�Y�vC9� �pk�&�{%�nA@��=I� ���g� � �o5�������t�v�ǜ�f�����ѧ�x^�����l���#�_�яg�/׫e/�Rg8�R�T��O>�0�I�q�z�]i-r��1��Ѝ�Eu�o3���ߔ��e�U��\[Z�G���q/q�C��m�}�GhyS_���>��I��JE4}B��������ep��+�hs�GC����%�uJ��� �]����BR�A����	-*��E >�{	}�x�cN
��
���=�T�e��\�!����(��I4W�,s�8S:P��p��5t��4�ᵙ�kq�C��R�Qb��8��Z�N}^Ҕ\f��<b��rI��#�r��h:��� 
�*|�����g�����K�nU"I��3Af �	|, "U W�x���;i+��c�Z{U.��Є>�@.�<C��}m����O��D����h�t����׾����Mz�ҥKcz��4��l�����S����(~[�%�,��l�]�s����R���dR����DJ�$R���Ʒ�p�F#����� (�%��9sJRu���L@��L�ʺ�H T�7����R�l���g�Q��#@��' &�a�t�9G�&�����F��0J�M���0ר|b}e�/z���,���F�`����ߺn��x��(���{�RP+߻;�ԨT�����X�ݸI��6���.�1X�ѿ;��-��3 R�)��U����������/|�ϜFv���|�L�:�I������G1 `���q�V�8�QZm��W^�k�7��c��o�ޠ�cǄ���+)'<�DIة�%�(�nS�L�LBWR� +���h:��7���=�-*���^!��avB�Ht�2%h{F0�C�6?=GU��QpL+�T���4��r\���%�2�*�ޚD�&�:/�P�p��p�l�9R�q���zO��W�R�Q�� �&�(t5:��ExL%i��`*/�gBjN$@���X���8���7���R�ZU'
�TԎ%�g�-�* ���� >�G��o�ݩT�
�����ϋ���^��˗/�xP�1g�i6~h���թ7>���}v��O�g���G|ǟ�M�츁(���[��UA��� *�,�����<#�~	��í���jg{OH�0H��:uB���B1ư��p Q%�%�5@���Tš�eh �*muR�Ԥ'<KM�<*������A����ˁ���|���Ź�W/_>���� �4������p�Q�O��S୒Wu���l�h�{ᡳT�ۣ�{��#jU�Щ&�/�P���t��]��Qq�*����Eä�}��';��ʵ���N��ǻ��S��ߙ��üٵ�ܲ�s��A�7�:��2��cz��jy�Tk4��9q��V���6�F�� .��k2Z8�d�b -��4U�����ͿW�-�<���>Uy����X֟��A��SU�F�1�-�hR�/Q!�4j�*���Q:���H���<�)��$d%����T�)�	���ܢ!�hS	�܂���8�4��ɤ}�l�l�h')p˥�N�ˡ]R���P��
�w�M5��^�F� ���v���U~ ���W����]�A�����F�F�C0��iI�v���0�Y-������e���^��Fq��n���_y��?��û�3�4?������l���8������<n�y������g4��M�#|����e����f0��s��e��*���~,�F���z7��KPߝkhwv�$��{�Mm)���s��qL�΃*r4����(�����$ewlM��+]��ew��%�P4�*�*yF�O��r���ɷ�Mb��y�"��G��?qj��'O�:� �[a�z����[��S����y���J��Z�����A��j�&�<}�����m@���Be�['$�0L��]!?�����|�J�@[+����y��v�1&�{��_J��Cn��������F�NPe��_m�+W^��w6)��!��z�) _t�r��Ry�ȋ4�CS[)��=	�X�n�k���U��F��ġ�ӽ4! �4�bI�K#Z�4�- S���"%F
�<+Di�؎�r����oZД)Iܳ	9��"�*>+p�9�HSn��FR�R��j<��Y>���{g�2%�$⤔!=_����@��u!9!B�&R��H��f���9J�W�mOHصz�!<�W�^��6��#���LlN8F�6�8�4��U�V������D+]���ϓomm�moo��_��_����o�?���g7M��]^(�?pzR����zni8�?����@�M��Q�Y��7���	3V��E�yQ?�?0��wF�Q���
Ȩ�i�xY)�I
d��Ԁ�0�h���!�anR�\��m��2e.��������,-//H$�ΓcZ4@�R��@~����gΞ���5CZ��+��w����_�K%�{»�z�<6�|��ᨿ��ٗ�����O���7g�o�a8O�q��|zp�k���T�^b7�2`�����|��iZ\^�+�� Tl�?�L�sK���ݧ�Wc�N�ܝo�kKT!��##H��z��\�ƫ7���x0|�0�B�%`���я�B۽!}�ŗ送yZj�À�ܥ�Ԝkэ�Mu   I��#(6H�4M89�F��iW$�n�	�;3t�0��рR����*� Τ��iQ�>s&FdSpEg�e�ܦ�(�'�=��kn&" �B���gC�\��cA�Myn��Q��1�$�]�� �:�f��F~���3�r�4�)�2�����[��L?��(��%�t����3����#c�ܽ���Ҟ�� 	r6햰�*�2�ch<-|%ߑ"O"ě�&m�-M߹d��K�u�c�b�8���_f�w�_s�����p�;s���+���C=��V�?3�4��������h4z�����������+��(R��2�����>�"?���U6�!�7�~��p�.������c�x�N6
?�:�S^���`)���V!�:$6dm�'���Ί��J��wV�T�Σkġд�Dy?���T�.}�T�{,�3^�>���7���j-�ӱc�h
�9Q�����}4�-U�}+rL�"�Ȓ
RJK�Q?���_iի�k�}�\>�9#w�y��J}c/��������8��,I�w��,��a7�y��l�S�^���ߤ~gHK�%�-7h���p��G��buo��3��O����|������Y���zcc�����T�ϤN�7��x�5�z�.��޸Ѣ�ĩ��;o�H��.�c�#�o_�$*�LFfD!�a�Z2�UR��S�&v�^W"�v���N�
O��,��t�E��0D -�xd{�9L�hXjT��9|h�8��h+)p�
Pf{�I�M�SZ-8���iqNB���y8��2aOLW9=�̨�J�a�)?�T�A�I��V�a���3�. �D�[$<�A8�Ƙ�N.�o�r�:�||�*M��g�ʥ��>f������ʈ��m�{�J%���E�ͳ|�\��q�D��,M����֏�k��c��{�n��֩S�~���v�@�l|���!ѱ�0��h�b�ď�I�����g����i߼��\��W���!)M/˝��A�kl������J������ΏGßq]�ggJA���%OR�rƱ&-#�M�[Xp� |0��H�`�.�	)8�JIE��e�\��ۥ^�/�o�--�(�hF��1�F�G�:�/��+�Tk6d��:t|z}t�'Kc��}�ꍈ��(ٻ?�R�����z����\�?/,־<W��<�C���AK���9��������q���y�v�`��cg�ߣj�I�9I=�F��ģ�\��Z�F���9��������z����vs��߸���.-ݞ~/ �;{�[��V4�ɩԨ����/\#��%^ \�'~���i�?���Qrh��Z%����T���ƉhIƵ(I9?��&���YT��F\���I�kyD�B��o���݀�ȡ�_Ab\[��Fy=���_�������f�����H�DAlS��5b�gqT5�2�e=%�Cm[$��ƺ���T ��x}�`� (���S!�KO:��s��h6���g�9iz?Ri�:SW�w^ɗh�Y�a<Rޙ_��^zI�jq\� 0�4��8!v��r4�$6�M��� ����/dp�7�k�F�`�@R��]�D�y�x����`�� �E�����N�ѳ�A��_y�?|��f�i6����?��a��~{��,�~���Ӽ�^Pvj�������/� ,w:�m�ʯو�y}���y�@��Z����,��Cy*���i8���(�&��~>Vr��y#U�x�5���nn��,����=�h.�̸q�9H%�v��t0�!�8�0�6Q$@FH�HH���S�/i%����C�ǉp�z�`7 $��{��ӕt�-i�\8��j4�=q���5�u
J�)�ˡ�%���Ȩ�Ԙ�]����U_��?C���2LC�M_��*Q+W�|���?~nǙ���räҶx~�O����0��W�!?�n+t�j�A'VQPb $=�k/�Ɇժ��Q�qb4�}�ƭ�������|�k=��G�3K�c��U^��/����|����/\{�n�uɫ�$���ﱴ�,�A�Kc�gDBȓ�%m�MJf���]F�I9Q��R���:� �o��u{{����^�28J�(������r�{
Z��6�N3c��ݟp�H�����c�c�}�-w9����4]F�j8�wLY�g�8#!VB`��4��!���x_	颢�ȅ0���<�ҁ��ԋ%RTչ�ݼ~S�L±ʋ~����jHQ�KT���BG���~���Ku~�ܲ~*�p Xq�V�N줡*�܂Ǒx������������O}�������/?���ofn�4��}��-�:z$I���i��Y�>����t�O@8/�ZG?�kds4rB~��Q+�O��ü��1Prlx7���e@�޼������`��Ȟ����\��z/5�7�mα���w:����DQ�>��.A����h�T&/p�5�6	a��`t"��X��L4I �m��Q-�|1.��j��|��y�(��4�Z�&��űV�)@��Uꣁ+�o
k��iqq���Bmw��C�r%bs}6|%�a���(3�}
�#���q4�˒��%?����§�Ǿ}���������D<�t�_���	�PP�a@�죃���e0�y�$����Q���eT�A�����B޵q�Γwn�|߱�����Jn�Y��ί�k��,/�V?�_�.`));�8��Ej�\%�s
y��T�CD1�VHye��-9ZI�K��+J�e�V'xR%DKT������^wepjR�C�*�ݐJ=M����!ۨ�;�6��PQJW�G�
���nґ�C>}����)�6��+Ҁ�iS��&:LFr�4�_�PwUS
Q�R����f��>W��
���D���W_}U��h��Pt�R�+=�ՈSC�\?_�e���2�bI�rM�s�E�F��� 4�ةF�]W���1���Y2��n��h�?��/~��ի_�x�b��h�f�i6�h>�s��$�~����gy��搓�F�Vc�Z-S���~5��j�����8N���q^0��-Kͳ	���0�x��s����$�����F_�)�� ��S�j�	O,��d�1�G�F���(�6������@hR�I��)U�Uq� �R��l�:��ϩ\q$k��k�(*���Oh�T�@�C��Lw�=�n�����=��V�-�!X�kȹ�Q.܃H�:BB��Rue�O��#�P��k*��p�I0m�f�j���ǎ�~e��t�ᇗ��,=pÀ��y���n��~�˥���ل�R3X!7/�7(�E�}J�W��A������`����͍'�_<y�tu����{��E�2=��U���C5�����r���p�B=�!��+����'��5W��L��x����(���&섇A��]uj��jrj�{�/�"�,^w�1���5�0� �n�ߟ)?;���!@u/p��xob̐�s�$��2�F�R��,R�� 4��I&��@����z-��w@3d�Ԩ��֭;t�fe�uT>�f�sGid�HH��\Iy��?�z%S��.�r&��p6�}��:�|�0&N~�!Ք����>'�������x�G�N��<�t�ҥ.���4͆�)�:y4��M���i�=
���n2�����Z���T�����/��G��=����}?3�(�����3�59�x�{�J�4K�؀<��n�/��>1ת~*���A�No���s�G<?8JF�Q���?!���b�u���p6�W�02�5ՎI(�\���+H��0&D�Tb@��b�PVO-)	 �#�U�	�%�%is��R��EBD�رc�����L��*�42������;�`8ql�[gڥ�ᐆ�^����>ù��5뿵�Z}����g��֜���@kH4w%�>6G�̋�C�[9��$Oĳ��� k�]�8��r$��18�O���>��h�Tu<��!=�5���g�V��Og/��j�F�;���d^�n&Z��NM9��rH*�R>���'"�*+DMp�9��zkA��f�78���h��B�	�'R��d�m2M~�n���� �SK"�O`�ht)���I��`�N�~^~���"���fR��L�*|��W�}e[�h��W��E���t���;�$�np(/��m��ÎX�X�O���64joRD��D�I"���9L�-��m�[�v�T�_��bJ��	�_����������^�m�Y�\�����n��/��K�������ӧ;o��4����ߟO�������<�����m�Ɣ��t�XX)Ru>/R�1�a��,�&^���M�m���~n�fޥr4N�i��j��,�k<m�q�����J�������o	�m)ח
��#*�(iTj�{�b׼�~$ ��G���6S��{�eKT(Q�_�%p�؃W� ��rJ���W����P�� �j���4�4b�(gNs�>$�;�7`���Σ� L��V���u�Q�����y�����l���Qu�����o�y�s�A�?Fi��㕚�����;�yO��*�:Uk�
��|m6�䗫n�6G�ܧ��o��r�U+���ҙsg���S��E��`�}���r�l�V��R�l���c����McZ�[��tR	�S��YW�����c�7�R��٩Q�� ���6����Pș<6*�~���*��'=�9޽���0M��!~Ք-����i8�D����sE^�dZ�8�r.�,��hZm�JF�5�ը5��������>	����;�2�بO&p�^����J$˶Ù��G��I�Q��
��z�)ϣ��W�W<dͅ`/�I���zOD��#{�?1?�n�}�֭[��]i7M?�b�QD�i��$M��3���,wr�c�&Z+�a�HLE���F�zLG�����k�1ZDڊ�L�%-���၂G9'Av� ���k���\���ܨz'�B� �'�ƞ
�rY��������C�i#; ����rvSف�Ύ����I�u���!@���B�\[[��h��Q�^�>Qx�p��sc>�0��KLsM"�[��� %{��Iǟ/��� ���<'��j������{�>��v%
���XYqz�v���۽9
�����Y�>��N�^SM0�Q���DU˵*��Z]\%�:O#���Ô^��C#�D	�rJ�h�hw{[9N2G�Уc��,`�%�S쏺��x�Q�6,$��y���ṁ��'1�l���J�*���0���l��H-��K��p� �G۪���F��L�-��Q����Dn&���t�����Ñ�>vʶ t T�A<R���;
哵-сC�mS�eJ.`���x�WHu��ͥ�i?ح�_�¶�#@
�-v�ES���l��kt��u����T��G�d˽A_�ڈ��0h��B�L[\(}	��;�B��6Ha��X�P%5p]2�A���N�{r0����|������w����3��C8�2�1�Ic�	^(�'��i��xz��03%��k{e�2��LtI\�)�Dd�̴��kx�N�<�˛�yA>��ˑ|:�i��:䛪��z���p)�KF�3"mF2m�ೡ��Z+	�!'��F���Z���KV���W>7Rh���D��9��%�Ʀ��_4��^���@#�*���l�m�,�Ch��<m�(bC�NaC¼�����.?�B�����b�/揭_}��c�L�{6������>������:��?�y���(��K�Z��2�@5���
s�AJ�����{��1�ʩ�s�©����J�i���؜�B`���3M��D<L�G�\Y���ng�J��T�<�GH�����Z�����/�@��M)p��G���4!{����4�۔����M�}'Q%����@���?aOF�!;V��@�T-Q��(��P6�����@�[�GF�a{{�^{�u�M�\;��lk��@�P�lf�	�9ov��h7Iɰ�Y0׶R�AN�l6ҕAO��Ԫ?��u�+���ֳM�UӮ*q^q?��c=s�n�o�~�}�~�w<}������0M?$#W����璈~���eI�O�*OrG�=!7��I��<�Z�,"���}�9�h�B�-���JCI�0��+�B����L���&�BrI��?�")3~��X��"���8�R=�R�]�&��j0�	ʁ�` `�%?�J�dUq� �&�>'Q�� D��U�hi�I���FAɤ��:�>uB�NLڍ�oB�#-P��7����?N�h���/T+�G�Z��?���(���7�⬨}����߃n����뗃ˮ���&8�"�k3�o����E��1��e�5ʴq�'k �_����DCYQU"���T�툏] I��!��
�bCw�\2�@n��y�3�ߚ�c����]{E��.�ƒ�˄(-G7i$)AD&O�7$t��Qs
�m�i�r�Z��8:�K��p��#��T�e�DGJEq]�F�Әz�����l�H�B�����3����4�u�^�:�h$^c�/��}�W8m�vlk�ޤ~�g4�ܢY��TR��ʱ���D�%��)�z�..��.:t�����HQ� ӶZ�^�ı��Qi��A��p��,��&�O��d�������~���|n0���իW�z���[��띁�|@�,�Zy�A�{x���'�|k�M����Φ�	�b2��.&��1��T������Ns,GJ_;Cy.�^��0 ���B�R���}����;%�.�J�2�fY"=�FE�ss[bݩx�r�oGy��`s�H��V©rw�`F�� �p��M6
UZY��r`�C��@�\�V��(T��V��e��#��f(g)�i<������皟�.����o��,��w3̼y�֭��ӻ/���_R���g����W*3����:����^��������������h�i�x :�N1�y���HH�Q�O���C1��f���&V!H����s�IJ;D0�<�?P�XHu�:���3�=��H����_��L~�~��c��~�M�ɰi�7��cyV*{ �3�Hwzpۗ������-*�FJ��*���#��m]G(�7��ܾ}������a$@GԿ�D����!�d*��|��Ơ<+��Z�b[3������v��}�[�	�qp� ��8*�z)C������	�UO�����R�k�7��,�3��v���t~������۷?q�ĉ���^�@�<xr�x�~�'�0�t�f'y��P�6J�zD���dJd�"N�WJT8dKjm'l*�:|�(��J�k񔗄�a͜	�Qº�S�h�u/$I�@,,̓z&��.�j��曒k4+Ԛ�j���STnD�-��E�T�y
�r¿2e��|�X�C* $o)��[j��Ғi�R�L4)p [�r�eÛ Ԍ�~��L�R���4�MyC
���;A�������_{�폟�sf|����S����Om���w��_���.��K^UERSק�~J��ݦQ�k�\���s��kk��O& k�Tg��w��M��I�$�.W���ة3R����ǆ�Y��*%���d�}��D�Zp�T�^"��er�<�
�h�q��S5VD,4�-TE27Oh7���
I�@9Z��J?�� "u�R�}:l��uou�ܷ'bFv��I���DE� �h⑈�TJ$��Kq�#D�5���'��u2U9ܓw�i��^{�6��i4[��F� ̬�+ZW�[�ȩf�i����4�?tPX\���{�Ν;C_����Kj����(���7�K�T9�<����8*C^|��<�c<���8��8=�������k׮}��>�hz O�*O�wFQ���"�ǋ�Է�,s���FS9��ҡǌ:,���(�I�8V��4`K֜���߄;��(:r���a�E*ᤴ@��K�����JH{um��T6W"EZ�QJ�8��g��8�esp�����BW"�U�j4��q�8�<(P�����G��$�+V!7��X���p0�T�u�p�����r5����<���}����{6޼���)/����n'��?��8M/�^�b'���]��t�G�8������/H$��FՆs$���=�@Ã}�=�Pw���z�~�8�J>U��Tơ?���j�1#��q��DX�J[8�pt�^���j6h��)%TiI�%��8	��1��{n4!o�]��7M~}�4!�H�!�OA-�=7egs�RוA�8�4&A��T�t���p�҂ɑ*:_����/
;��.�8T'Q���-��ʫ���A+���9��٘�0���W��[(`��&Dx�1�x񼜋��蟉���$+�?T�@���:S��3Ԇ�p�12���3�u6b��\����Ź�`���z�����K/}�߯�������\ s����v�'�y���,K��ZV�A	zf%O�R2mD�R3�1i'�4��>O�J��OE̟�Ǥ/H�Nf���M&%�9p�q$��s�N�R��Sċ��� ��Bx��Հ�֗�g�m�%�!��:K�ؒTXXH�p'��$%k��\q�4~���"B9�0G�V]�.�;2׈�T��k+��D	��@3��L����&��$I�f��j��zq��G��/_�<S��XZr����qg�[��.8岳�7��v�������S'��G�2L�a�e�E�F��G�~��8D�'5�5J���ͻ�[T���c��qO��)3<��Ylz�)�S��T�]�MZb�UB��	Ua�?-��4�8�*=���]r��������7�t�?"b�
�q�8Ӏ)+^bS�Fk	���	��P~�U��zƼ����B���JH%��q�b"�]i�h�v畗����]v2+4)�B�Lq�Yf�s{���'����V���&r�Ϟ=K�Ν��h(Zt��j���L9o2�י|�i*�c�T�bB��T^TIN�w��%uK������[[����^XX�����2e7MЀ� {��	���Bz�o۵��z����L�$�<�7ٛ����V_�E'� 6�ގg*��"R�g�[qܚ���+�Hl��+�h��t�2~��)c��j<O�w8�g����ñAZ%�y�]B�[��iI6.��{M*�1 O	a�J�< t)�k�H$z�G>��]SQ�m� �����C�8�ܱ[�Kߨ�+_\Y��|����O�����l� G����بG<�olo�ޠG���;����	:��@ݾ:51O��h���R(p���?�ߠ �UZ�u�^w��>u6z�ټC��c4��H��U���T�P���kI�w��c/�3���Ǯ��y-��[�To��O ҙk-I�Lx2�[����qߠj�h�i:zt�q�?�F���0R�i:j��I3\�M�H�v+`��Ƞ���@�'-*M$�6Q��8M�t�2�%-ѝ�mi�b�J2}�/dJ��Lա�L"v��\�Z���y��O�#�<$ i�
P��p�;;;r��Vъ8O�W8�ga��H ���S�S�}��<���F��|n�9��Sb���p88��t��v��իW��{�,>M���O�ƿ^&��������c�M���B�p�X&l���Ֆ��1z(����BڴUna]p�)�E��f�J�q=�/�qu�D<�7�'v���0�h�B���@Bеj]�F�@���i�D�9}!@��3�c��7�h.�Z� ���e<5p�,b_�:���l0.�� � M��dc>�<�^�}�����O�-�^��v._����l����^o����e�o'����i�ۥ�Xu����9yJ���Ӑ��0I�(�<�=�Ǣ>��2�Q'��ۧx�����nnPwo����ed�h�7R���^�F��q�U��w,�=jU�-�ww�~��d����#�V�����k�7�s����f�S���k1���W�M���y��$ϛ"���h�R��n|�y�H��_a;<Dx�Iy��C!sb"���GW��Dk)O����WK5I�0��홨��r�/��	�"�Js����lZm�rZ�U�0��`�D�$��i�}kkW^ W )�D-����5�8�2���*H�=�p��	UD����DZ|G���_��k����p���ǿ��/�����7.\����ZY|�����O��x��q�4����&��q��Aƴ�@&�}�h���7N��)�F"Od#V��zSB" n~��yM�9�z�=,^��`���J��G�9�i8��� �\�nP3�v;�1��Xh)���Q�&�U\x+å}I��G���5���x�E��P �i��4����g�Z��l���?q.�٘������V��$�W�,��6���60��j9y���q��N@�QgR�A��-��O-v0��ޥp0�N�K)�HM�&~Ҹ�G;�6��h��qZXZ��F�F�G}^;�MI�=(Sk2��vh}�I�Qn���W �x��36t�>�s��4��j6rE�'�0F��;�s�TO�3:�%uLj1ub�x��z2�v�D�.K�fA��B`�Gtű��$)ν�}�~��8oZ~h��~ 0S�(��$3�#�j������8��g�IjN�eiQ��y�^o ��}k� &p9�bc5�
�[T]�D8+$"�+q�"fS`�F�˦"Xj���"J<V�vw@�`��Q��K�Y�0���c���z����k���;�x���h�D��^�($FJ�	�fEXӢw۽Z�Li!ffD��\�Uf�v]�`Ѐ3��׫u�3�i��P�ʑ���ch�i�Ա������ 8A�?��R�2�4��kt^����M�VU�4�T
j�?�r�ڹC�0Ѷ(^&�ڠ(�~[uG���i��>H�� P~V4NU*ɴ�V���(V}(M%*�<
cQ�����a����7[��-,,�ҥ�W����1��wwO����[=�5�݋�v7�a^�Hm�R�gO	/i���Qq�l�"H��7�us�	��-Z>S��mC��Ow�(�ߕ�Y�ETS1h�y}��cui�z��[5j--Qku��Z-j��{�.��Ր��ս}�u*���:kUj�C\(�w��1G#�e%S���t���C��1Π��F&�gۑؠ������"6��F�1�m����mD����RB��i��p��q���R	�'5=9'��L^Mb+�9 qPX��5p#D�p}<u4�f�z�����!�p�b�*Cc	�����3�T�Y~�o"w�"�w!����qZ^Zg��N)�|��2����8(�c�[�vo��ن6�8!�_1��,5Q9i������
�dN�o!��h 0� ��`�WC�ЫJR�A%�z�x�9�D�/���m�}�ƍ;�����Ǐ�!�h�������Em���+8����)R��CUS�����DX��l�(6 �hŜ�݆z����w3����ȑ�(�~nAbO�x�����І ��r���t ��cЄ��h��j5��[�5�9U��3�|�g�B�l��#1qTh7Y7��d̾X�f(��x��R)p��ı����+��#�Rp��f��+7n�w��%
j~g������.�MkiyU�!����+��(�(�6)��%j��
o�A�Es+����穳}���4��o���#p ��wnR����
-����ʲb��B��[����lP�-9Л�ת��d�,��h�ܽ�����t��!�8�Na;-��A�բ�I�i>�T_KW[6e
��|Q��>��J��o��mi",͉
�Rj�!"L������d���;w6��͛�*J�������=z�i�Op��C�$����qQ/WY�T
i�b���!�j%�F<\S���0 �[���jG"�+K�"�����a��V�xu�a�s:R�i�IH&��������'��@����_��*��=̏�a��}�~��_��<�p��%g����hz�z��S�A���}��!�d
%�@{��P�QY��������p��>�/� �e�㹓���l:�>�/�)�fIj+�����sE�����ќ)�*�s��
�I�	"GR�3!�� À��@>f���$�S.������ㅅ��y�����gc6�ǫ���3�W	�S������}Iu�H�)����lMuh���um�(�F��-�U�$�R�jyYz�Ux-﷚���&l3�\��6Ү00���Q�\��i�ӡ�ݦ���,/P��g0S���X��7ɃF�L�Ј bN%����h*~NU_M��Q����=�Tz9لem@�u�cN[�ؓ�Ҫ5_�J؎":�F�+�F�ȁ$��RqV ��fqT�/8�g2.�cD"Kb��\�Bw��5�jT�l�~N l���v-0��^'�P�_���`á3g�����4k��A�����&|������*�&}��ն�a�)��d`Sa��}ר����vs=�KO�BL������
2N�	�q���F�PE-߅�[�Ǭ�g}��m?��W����K����Gο��=�x3��`C�z�>dE+��H���i�4]A��W̥E*n8�P�~��9��9�U�ߖ�b�j:��C��+M.v�p�x8>x������Be�����"{3�^!n�T���C6�b�4}h>�%8�~��K%x��<%�h�x�l�>����O�}�m��"?>S7�x��Y��lo�{��81�!Ⱥ�9-�4B#i��e]&W�6��lĢN홊\�"�.����K�Z�Z'֩��H[w�4�i��JJ�1DJ�ܣ9������)a�%1�A��9�I!�
�*٨�NP�=0e�4Dp��J�9��+���!��M�d�f8�����([KT.��M�K�n��)�E�2J��7��j=4��0X��P�f*�+&�o?/l�����%�L�"SI'v,s�Rp�+��D�S[y�8�}�[�$��/б�U�1�=�a��U�������rmʒ�Φ7Q'��a�+�G�ە4!�_�>ͺI��L�|E?=[i�N�Z&�cn���0�l��쉤Au/�ߜJ�D�t�������h���^xዏ=���d���h����$�{S&��O<+��7�#�7Z4q�S�9����r:�g�=�;��z�_�	��F�S��2M{@� �{�3`�ƻ���쭜:.B��O��j�mD��?
G�IC�ͦԤr%�#u j�����$N����}��}fu���ե�痗+�._�<�E�f��>.��x������p�;���b��Q*kmeu]��퐽t��qTЂ��C�B֑�D�t�>�n�p~|�"~n���5Kt�y����vh��Oi��.��ϩQ��Ƞ\��<���@6P���H4�J�#pU�;C�=��NG4Q��E��p�,h:J��������d�t���e�)�YAFO"��?gڡ�3n���X�V�(W})|��+ [���V��riث�k�����6mܹ[Dɥ�g�kd���T��Dg|�V��˵�Н���^|.Ǐ�S�՘j®�*�����?�- �T��<�Ia��GQ)�掶xI�$���ߠetz]vR���)4� ����s���c�%
'�H��ܱ@��I�.��=�|����~����ۇ�����ׯ�ٹs�/ܙ��h`Ww=�v"EN3I̤��F�E�E�r��{��V)�*o�o�ݷ��QGA�4p��sVY) �(��i~_�i��Y*߈�����	��@{�i'm]ԩ4�U��|w"�=��"����Qf��]7�S���znn�Z'Z���Oϴ�f�62�V��w�qF=v�F����ؕ=���E���8�I�;�*�\6�̔sX���pN�a��}Ԡ��k��B��E�U�-.Q��vve]��D؊��}�*TO�)SŅP-6h�M�@Ⱦh��4��s�l�� �0��v��PLE$��Fzݑ�<;l�����jJ���Cj���P�#\�>ۛ��B���j�Z��%��KE��5�&�/V�I���lJ"37nܒ(�*}��1h?�2M��G�4i��"���6���=�`���u��Cߺ�T�9*v��x�D���v�2�����Y�b!����Sn�ʩ�Mw��Go�r-��4�k6$j����ك"U�箙����!2M��z1S�m��騜�3}�k�\1~�Q�ރ�������~��S�輘��h�DH-g� c��:���ׅ�y���\�im��|gۧ��}�L�mX�w����0"�ލQУ`I{�9*l�L��:���h�E��H��C�@���[�q���m��tݲ�TF	E|�A�=�a,�K�sq�D!ʳ$F����T���O�<v��>���,�4o��Ǝ�4��F/N���j���$��퇒f��8��.Z����8�
�"��M�m;Y� K�ĕt�x0���S�7х�uZ[\���>�ܼC{wo3�H��1KD"��:LnY�2����Z	�=�q��UR�l��iǁ2i��q ���ؚ~���
OFZpgr�H�^S����h�}�ܠ���PU�n��Ғ��[����h���L6yW�PB�vD�YoB/�t��nn3�(�ޓ��o��YGמ��8����F[���t,��'O��%Q��&T�	�q���!���m?*M�!3 ����(މ�ȍH���U��:�q��Tn��O#s����i�>r<Rw��W�k��Ş����i�߾`'i�S*D2��M��>�JZZ��2�Ng����	w�_��:ڂ�3��`��'R�po�6 v� �B(���)5
Ű:"Vc	���1�M�%Z�������hnӁ�yR6jD#�#a�۵��D�L�x$�	��0��P�B�F[T����¡�WꛈZ�J��V���f��ыg��g.���J��V[�Ć=�;��B�2:���њ��Po0�����(���xO"y�h���I,��$�8D �y�lSEN�Z�(z��>�%������1^���:�o�F��>��:�#>Io5�	
/҄�r@i5��$���r������'M����Q�Q�d��M�Y��]U���b��PI�4���J�o��xM�IhЦ)/�ڹ�QW�X6����h�R��S�v�-�"�4ј7W %���$�f��N�M[Z����V�	�Y[[ˈm�k;;d�!�&����%!t��;Ew6�
x���-�C@���c�Si9e���3N����!�<U<w���!�P� ��H�X�9����yM��V �,w��Є�٢t�0ٗ��^�g���?yc�����h�bHD�2A���N7���ÜIӬH�)j�M�>y����c�f����P����ˆ=��1l4ɦ�`νx��	�WU5�+�1PѴ�i:Yb��P��j,���K.`���Ry�B�Kkt��5��آJ�.�ݠב4\8�a8L�q�w��:�/[_��O����g�p��`�QD�6�ﹳ�mluz�4ʴ�vL*��:}i��t�D*��A�.����(�h�M������&olȔ �d���K�l��'��P*�$* G�wc����'hy�B.oƛ7n�h8�*��H"&R�oj��`E�� ��4p�apCE�pJ.��7��cJ���M�X�Qg�znҌ��$5���Uu���p�@��3��=Cz��ר�2M۾��ՓrE������9W�Dv��F�'�/�x������&��߶�}�D�wB��d\Ӈ��%)���M���-���U��J'h��z�粼!m�N���(gN�����pz���8fz���V<pd�Wiu�m�^�9��]��蔆����9�[C�BDZ���
ތ,�;��V41�=�>�oܝDI�m��qYg�?k���S���E�}s��1M��%��&���XOC�֓p줄_�4�{��t4�tT� c:be�%�n�<�n�hfHe��<�'d�{Z_C�R��*�X��I���A9/�V*0��p-Ξ=O�nݢ��=	�2 ˓t<��p��gߜk�}�ĉ���t��k�.-}Oz��l��/�[!�c�7�|�3��j�+��&�PT�t��f}w�u�]:}��[�6&�J@)o�A_4�*����!���|̪T��i(�ၧ�Ө~��D	�A�or�,.�S�T���["��8�;5 `[j�^��mt��5g����4���6*S׃Ȉ'�3!JO��i�v�Z���y�6NISn�� �ˑ��Mq=)tɋ��t�^�?���!M����U�`xHZ<6��{��}� Oi��J�D�N���'�@�D���U_��JcM��"7Σ
>������&;����"��e�H�����j#]H�J��3��q�B��#�/�%�IMT�D��%O�����Ѥ�I��S��ψt�������;y�-%I����0M��/�/��@E_�m5�k<77�����d:L�p�9.M��^�StG��d�tɆ��HЄ;��C���H�V'G�����A��ɤ�����K��Rr�+w��q鋴����wci����K˟_\^��r��y�ҥ�H�l6f�4���9H~��Vwa{� )s�G���"��S�ߓ�����_�n瀮��*����U�$R�WOE���x-��ze-�M�H�}4{x��M�%��ؑ6����*���`�'r�;�v���t�����! ��.
\)�r��DS6'��ܛ���! XXqK�~l�?��[��i9ی%��j88�B*�K)�$��F�lt߾?�	0`�Dx�hD~Y�Z�cQ�Hz��+*�哤&bF��&��g�d�u&x�{�}e�jW��@h4,AzB$Ei�T�fVk"6F����6�o#����~�je'fF
qDO�I��-��}Wu���}�{o�w�MR�$6�6U��|�����P7����H�&F��S�������UW<�P$�uzM梫�"�x����"W�mr�G��,}+U�
-
Y��(���8�u_��ct��[u���\L�h�M�)�S,��L2%\8[��n��T�AaBu�[$�.��T��.��7��t�I[�����	7�nto�iS�waU7�M�xϳ�����2��f��M�nD������R/*�MǙϘ��#�i��d�8�c��X�� �����XTE�ظ�����j�]yr�ğ~�ȑ��4���yc�h��k�����N�SA^B��{�x��X��Qh�4j�M$(��#�6���m�>L��85y궫U��C2_[P�o�W�#� ��ޓ�$��/` ��n���WdfǅZ�xc�^�CS[A�"�Kq�jh��8Ib�^�4I�3WD�nQʍw�ޔ��-���Г������Y�M���c����ʱ
�g�IN�ͭ�D���|�V��Vollѹs�Ե{gRM*�nu{d���Q�V�դ�H�'@���!��)G��L8�0��d1I��
8��vP8F�`�K�ٌ��]���5Z\XR9��H|����F�)�)_\A=���>�V(R)Q<�d%)�i\��(U�~��>!�߯��TU�Z{L}O|Y�?�7��t�����h���^�E�S7 �� y�#��QM�Zm�F�&���Q�� )S���%ʃ^þqcK�x~/��OW�8��{�3��;>�jL�r� }�0�%d-m�CuH�TD$SM���4�-����3�4���D4<�w?1�Q/�W�5x�ȎɜA��N�?�����%*�s�B����4�I�ܭ�<��@���a�T���G�P�ZH�1 (�T� I�0�'��}���T-�)�Rz�~���v��P�����uJ�����"bkRx����3ևmn4���C��_ۘ�+�u$F�fߴ2n�$0�Ň�^sJD�b���'&lxY�&�[%�l �7٬w�����cBS���e�4]G��N���y�����P/�&j�dIE���86Y'�_�¤X,KU��ݎh2)�H�����2�����(<9N�D\�Wwm����K�J�"�P��i4k�����`L+������굦�\1��	e����U��g*ǭ�C}�������^����M�h���M��4��!jLX�of��m�8��L�T/����� ��32�7�Q���n��[���z�~Һ�2F���UK�o��_��3nw|�`8.D�rE���[aј)���X*���. �`���s�Aw_ZZ��Z�h���+mR,����Ij2��H��hC-Dh�Q.)� I��H�<h&uxA
�h�T���%�G؎d(�)�b���k��B��+���Ii+�b
��>����c�.7�S4�(N�h0�y7�N�Rp��YzZgΐ��X}zMd8M*�'q�T�]��Z�o@\}��ֳ`��r��SwU���4�,�J4�58~�JM��qN�O\R΍�k�t)��=@��}��y�+졐��I�u�z�6c��*��5e�%�,@ ��
�� b�;J���\�)2�[P�;ѐ��h4����@w�Cm+g�S��4���o���ۦhum]��n�
R�Єk%�,����-T�=�G���p����Io�fZ@*��HH<�.ߔT(:�4 ֑H+������hݤ�7 M������7@���� P3�Ѷ(*����	29�~��_n�qsE�V^W����9�݈�$�cT�|׵���0u�X���������2��&:������	g�2���-� ��Q2����ձ.��~���`ƭ4f��͏,��ݨ���mv8�!͖
y5��W[�T%��������i
�B�/�)��?R�@�K5j1�qy��%�h8��-v���,>a��3�p�H��`��ףl'�˴��J�h�K>Fڤ�4��)b[�O�".,��!z��9��5�ql����ϧMkB?�c]7:e"��)�l� C�Hq3��&[�Y�
��(�k{���-yδ���   3����Ҳ"�{�n�ͤ�_�7���Zɹx�i��L���A���Ӝ*|�Q.��<$| ��͈W�H �Ч��-��,qNm��5	irr\�W`�E�k�󴾙�5wf�']ܡ�}�P�� �kB��
׫�Q� ��SUvѐ r���k ��R��*�IT�5�,�R�w�oߞ��;��[h�R�v�\��n����8��/�`6����54V�]O{OШ(�%a������~��(`ڧʝwnș�J��,}�~EqW�7-�	�ػu�5r�pU:V�U���������vC��a�Ѩ�d��"��^�t��@�{0n�.ӱ}��z��\�K�y��M31J&�T�թ�N�M2���.��T+�(�H:A#�ϱ�,U�_��(�L�s�\ߠXfH���!JF#�V��µ�R��S�z�H&Os+=^���4�1 �{$���$R��K��G��t�b�v�LU��[�t	�:�g+��BZ^T	��7|"�?�TL�=U	g��M�#���H�]�&2��TTL�7]�LAZ ��2eB�c���/����K�>��8�J�	t�s(�����yj1P��DbP�bT�U#tG�`rN�!�d�b�`�H� N�Ғ�� \X�G*J���C��@E*���v��#B��'��(����+��ٲ�i묅#z\NH���*���7ic+G[[y}���j���$�=�;=ǿa��C�=_K�!�Ui%[� u��Cv״�$���J������[|�����x�r�Rm�ؓ�����s[d��B��Z�m�A��<�#Z�KT/�G�-��������IU3�H����S�ZɎ� ��lٽa�s����H�V �n4J�W��[T��U�_AP<3۳�!�ɎO����GA��R-_��عH�1���X����7[,M�	��P�nP��/k��.�ݠT���bT�M!�g1
�k�{ǄZ��
�B(�a�)��[���*�6"[�"ex��6r�֔da��>�b��Z^0�D��P)���*���d ����U�޲(l�U��V\!��E��	��8�qDʞ ��Z��	�4��/!�[�O���������@��8ԯ��R�|���>mt�T�I�S����:/Ъ�p��a2��CY���;x���C4��@> �*�l�?�����H\E�I����Pl��T��|�Z�N�k�6�;ZM��ay�w;l��(�LP�R�����u"�@o��<*�J$��"��ڡ�_`��fԛhoG7�ŋU8W**m[k6����X�He�)�;t��KU�(XZZ��ׯK�s!�.⨔@�I*
l{m[^�����	��C� "P�z�2�����;#�)߻��Z����?in@�-6���n�HW��U��T��>�u��OR�ҡZ�ݍ��EB�N�����s���L4p{�q��޻��?���T� �^o��ӁQh�[:��58R�.�G(��+X"⤚@z�aR���G�x�`O�<11��={��i0�3�Z+4>�\�?Qí�K��"'c	��;T��=�<������J%��<�.4�I�0d[u=$M��
m.�u�����¼ g��w�RRs\&+��P�E6H*m�H��HX�����Ш�������XT�"�`֑�sF�������m��
�� ��(U,�a�l7V��]bu��Ȓm�(����-EYp��e�C
H��s�F(	�@�V�����,�HY��Z�'txx�fg���sy��H��G ��]�uv�xn��F�ʆC��B�\�s�����	�iD�%b����:#r,8/����*�~�*��:̱���u+���G�n��ڈ�(�{�%OG��]��aRdl�2C)�(�<�����A��M
D�z�A�mpU�]��V����)����z�;�11'p��5�F��s���/�4	�h��F��h��6�@	F�l�V��;`/ �7V��T\�۲���EC�È�Q���
��N�Iʌ��R��~��6�mהi����\(��G��mmp�D�FÒF�t��]%ۦ�zk.V�K]&�"�5̉g@ԭ�3��10y@|��(|�->B-ڷR�}~-_�4:j�}v�\J�G(�HS�^�2���TI:"��v�J����ũl��OV��q+��;`�V������.Rs�LRT����@�I�&}E�H�6��hcm���1M��d���3�*�Ɠ�&-�4�|A�j4K�!K;r�.Y=I��{��3���R��7!�]Uq���f��H���p=�`�@	\&  I�y=[��  "�%��ӭ�3|&��<s��YJ$�J�R��#R%`#�R!��Z��iAq
�h��>x�j�� B 8^E\�`Cp)�n����ۜ����;^ǹ�3�nQӖ�'c�U7@Ň�n��\,�r��m�$Ⅸ���
������"�j�}�jC\OD쐝h�S�5��vRݖ)���D�d���_�o�w5���� 4�"ß���KKo�n<�FF2�j[9������	����xr������fO�oNq��&F\x�mnLj]iP:I���ݰ�i����-M;�T�0¸�f$�$5WoT�d�S��A$�ժ�>�ƒ>�O�o�7�������A�i0n���ы[�'r�{�j�]e�Өwx1��*�:ϝ|�IUp>,���u�B��ҋn(�����*�%]�t�H`aG���^ݭ	Wgdd�� �\((R0r�S�,NH����Wfy�KU�+�.���(�KF`1��W���3��֍hX�����|�q2$�~�ӫ�_z;��9)��(J���~����<��H{)��Te���lEPj�$d���ש?P�MA��4F�	�"�@��st����K��������vz�Sp��!U�>=�tB�K��Т����<�2����
@]�o�ke8����*2����G]2�A��;=����� yБ�x�2�I�)G�zEҢ �H]�<�S���u�����i��	�U�����}~6��<?==�S�����|���N�����GW����ٳ���:p����Q�omѵK�hzl��vK�t-G�;A���� �a2���j�}{�d?����tm#Лh7�QZ��m����"��B �o�=�����j&��3��oQ�5:R�ԩ<�M�$\[o6�|>L�1���jҎ���G�͡��ѻ��E�	�K��9��BQj������hR9W�/j��C�t�� ���D�yN�sT*���|�|B�*/v ���J�b�"�T;a���p8a��Y_�R���ﯢ�� ������� Ѥ{�d��
��l�'�V�9m�.͗��X�?%���.�p�tt�Z��dw �]�K����l�6�:}�5���V��"-��>QH�\J8R�ѵ�BZ���ЄW�:���3C�	Q!67�������Cĩ�5ՙ��C��*j%\*��Dq��BX�[��QO����� T@1dt��o�\��i�n"O��xi>�t��Ig�5�F����8nw�5�d�����om���<]�_�J��"iB�w�{@/R��0�㕵��  ��k�t��L&~�+��_���CW��;o-^����O_|z������f�x}�����O�d*)�B�L6���󴴲B���i<�j�1�8#��ʪ(OE#���b�z'9!%��+�{����㕟���s=L&|kLB��Z$F�g$��q��P�������0�odc�����[t�����B�q_�I���j�N!,q�?�V���*�n ��Kk�n`���<�<5��8
@��R���}��NDt� �&�o�X*N+�9�4P��Pq%�����m6��R-ʄ���Ds\Ӏ6���X�-���$�����5I�h�n���
h	6K2Z���y[G���d��|	�������V��=��޴�L0vmRQ�z˖�=G��:�J��TXq5%�e	�x�xs;��Jst�_[�E�x��3��τ|�9p��Z݈�i%�*H��ȶ(G����D|�%gn�Й�`stj�B1׍2��:>��/��k���Le5���>)�ڲ@R����c4�P O�����ޱ��-���Tޡ�}�F��)�,�38R8�z��]/��\�����?�{t �~������!:{�f�x��̹ǭ���r�f�]~��ݨ�)O���ym��&'Fi����$�I:��/�����`�O+��ϑR�,�bB�D�*���vwA18�X���!���B��xd��P&���C���-Dt>n��B�X��ۖL$��dTah
H��� �tc�FOaܕ��k�Nǝ�N�`�-8�Vit!W��zg�OU(sw|��e�kl[
,Tȣ^e�?�I�}P8dK��oe�?,�>�T��w�vE?��hS�ޢ�����S�١j�A-��)�U�r'.��f�syl�Z����v�P�	�/�����_mj�T�L8���PS*l�lɮ�O���k�C%�t�L�����5H��ĀD���*�48��#i��wf��j�@���,꼸��?�n��D�Dh�A�h�=�`����F��:uJI ��&�;
�
���	�sR��dpp�A�[�7@�G�۰�r�>��P���2���~��2�	2F��P'��5�z$���\C��EE� �Q[']������8:Zf��"m3�%<�k��>�@KK+�e���Q���f#F#�C�b�Z��i;�nپV:�~��q��@ӯ���t������B'W��X,5�y��Ѕ�^w�[9
T;E)�����L���+�f�㰑����Y��w/aZk|�A�' �C�K�E�_�}�7*���p����(1�gT�&�ږ� �h%�Y�=x�"l�	��[�p;~Os��O����nV��(���t����5�4�-;6
t�J�|��t��E�ZSJ�'F���/�X�}h�Y��#���d{T�|����P���꫐l�x��B,��6>>I�
,�Ut���A�C.�����*@��g�vD�1��$݆h�Ĉ|Uq��ҵ��tKW�	�et�#�|�AJR�4�)�#h0utk��j�t�Nu�U6�*9"-�k�7r$g�L5p�8$Q�#��z�*��� ���0_[�TY2鏢�b[����J2��Q ���eB��Pו�B8����*���#�c?6ڐ������8�4�"��h7�cJ�E�����_�g��>�����Ŷq�X'&''��86�p8� B8n92����� �����:p � �Te[D���(��bs�Ѣr�'=D�E	{�hmmC�M���5��ojۄ�ךh>)�z���^I&��a�T���� 4������^|������v+�����4�K%�۔
���Q����kz/wL�f�DǾ�v�{Tz�@X��ۢiF���,W�[Ti�e+���u�Ŵ2��c�m<WU8@Y�QojO�?��醫m�v�Iǩ	��8����X+ˋr�0#�a5��P����s����$%2
��_�5�<����X��~_�T��ܐ���������-?����G6J��k3H�Ey��1�F�ꭶDeÎO)^�ꍶ�y!89:J�L�BV��+�teu���Qr����luh����T(Fl/2#��s紤���6��Q�.@���.0�&��t�Ǣ��Z*�T�O8O
�X� ��Quu�	B��~�� �j0�[� �-��B�Tj0�a��bK��D.��>��"N��N�ϳ{NY�.@!*֚m����p��HP"1�tBiIi�H��Գg"O��	H�v�0D�N�8A++k���(J�Ī�>�\_E�Ħ�NW{H��:y�)C2����#C�H��#����O^�mƣ���?c{�f��;l��]�Q�(��(o�Q�Q��7)�� P���k�s���D��2������K �n�T�~�\œ�mTC�x��Eh(��{z���nڶmR�;w��#�TjG
���d������>���CRq������������co�YZ\�#1jV�t�{�@|�i��?B��sh��Ѥ���/]���Ti�U��!��_ZY��V���C"]�r��yZ�ڤ����N!��I�wJ�g���#DJI�r�%��{C՜���Lx9&�dn�~����Cu��-�oH��MU0����=��4����t&�_��w� uJ��K��T,��l�&'$n%O.?���-7�<�rt�Px����2��jå0"��!�� ��ۄ����;�օ\]�T5ihb�2�6Vi�^��;H�5y{�D�HT�\�FG�y[�nU$��&��P�4�/JHav�@�^)�J/�t���64sY	��^r��R��HE�=�T���\'W �j�k��=�%����0���Q��v��{����zwgN�T�=��R~4�6SUi��������j\���!9x�~`���f�ҥK�+��p$�W *�Y2U�D?q�T�N�I�&� ���IW���r��tzvxx�k���k�p^�|��iD���g���نO�qE�<l?���chB�?���8P��
�V7Rf�.t�u?�L�B�|���ӫ���B�������� ��EE#h!������˙L�簾�j��������ܸ����ϣ�ǎ7���ݫ����^�bc���=ɤ
&�V����f��˯��g?F��0-]�����	���F��=����О]����4ϓ�����W����S4}�~��7Ov(���'�8{I���H��Y$xFe;i�ߔ��"���E�tŝɪ����w��S���@)��'�aRn*,���g����?+�H�S�'�*�I��w�t[�����T�P��V�3�hx�*o�c0n�q�L�����V��=U
S��zӣ��a��ttH�G�HȦIs=M�j�����;OPC�qvp<O�5
��գD��-����6*��Eg���$D5<R���'	8`łD�ca�"Dy��u�ȡ��5�ܤI���3pw�����׏NZ��N� �b�J�&|,��N9Z�IRr���������5TsŜ�\I�����%�	��
�w�!`I����X�V�v{{����_���tLg�Z�@5W�����
C��B�rչy�exU&b�cB@e(���LF@����(�-���畑��S��c���%��K�����֖�c�����>�	d��N��"Z��� �!�������
`��U[���H<J��Z�*
� c<	�PnG���|@{b �$`4`��~�5u�� ��yK����x����|��Ɓ���œ����w�����|�8������O��}trsw,�����;��?Z\��d�>����ѵM�"mň��_x�Q�ً�鍿ڠ��8Y�嶶(;>A{���;i�ѻ�R	:�7��c'���葻h��5�
EcQ�:M����-��Pi���wH��8ި�Ǣt.:���A:�L=���p�M�'M�'������n��j[���=���Ç�ǯ��u������O�fs����>�"��k<�/�`�-4 9��z�޵Z��O�/�58H� 2�f����� PЊ���T]hu��[�Ս���Ȑ�P�_[/7h)��Cu�qM^]��S��i%�g'�R�$�D�]��ja��Y��%�4�vFǡkNʍ:n"g"�\q�|_a�@v�T�&[K��#
�*߷���g���-�2D���7`z�i�*�	)?�Z���F��� e�0CT'ʈ���tq;�n7�3���*�#f���իW�a���y�]K� �cH���y�Os\*Z�hhLY���y�����*b`rexx��۷o_��h�>��~��ӱ\nm��V�AE���j������tF�	@G��� (#�ixQ���yS����Y�0!}>�R�tZ�FW�kk��n�yS���3��Tᡁ;��o�d2��?��t������ynyy۷���gN�<�����<����+�mb[������,O:Aw�X�W7����*�S�U+3��Q$�� ��	��3S;������oӅ��41���w�ɷoV�oAo�'���9z��O~��cq�\X��~�}J%�tρۨ^�R=�%�:���|���H��D&� +F�r�=�\�q�G�R������I�À'��C������;����n�nc�T������4�9<�:���|�ľƟ��s�f���4G���ʮ]��h0�Ǌ���f�[kt���]�!*��5^Pxn�-*�������Lcm��#:ލZ�3�Y
�#�^	�B+��K!F�P��2��Rjt�����u-�T�Y-V*��+�HQz>�2eSIi��Fd�略dQ��R��t�N�Y�6�K��R`g^�*;��	��L��!�� ���vT;��%����J9�&�_����t�.U���<W˩�*��z�F8�'�a�١$�f��2A�*O�w<x� ��l@4M=��h[��L�����})f�������Q�*��z6������kZ����!�������Od�#_��6,�˿��?��bP��8�`D��^�����T��E����G1��q�:���8!u����2C�x��N8Q�B���M� ���[|��w��E�gh�> M�c���۟�����_�S �@e|�'辣�Ы��AC�L��I�ͱ��7����T=}Z5��Ì��<��~�*~�6��<|;=v�m���]a��p:C�S'h�\���8�9	���{���m;h��hv�b|�W���]�hs~��l� ���{ǎQ�j�>��g	أm���
���h}}sM�1w���g��F���(����.�I�&����Ͽ�.���Q���Lx���,MNN� ��6u^?c0n��sW���Y,4>��t�?�`�AM(";aj��@
�P��'G<I�#Ҡ*��ò ���b��cֈS���8;Hh��U���>���잦0;P�J�� 5#��rq��4�d��� 89׮S]�A<.��Y��8�OD���`����{�%��kR�.-��n���!;ZtWyV����+�����3x�u�*hYQ�'�~��\�0��b�};$��F���q(i�ž��xʾ�#*����tV���M�8�|�x`�y2���(�lQ��}�
0��Į��7�Z�(��UqP��%�%���k*3$���f����`�j���'O�|kss�K�F�c��{��;� �6�t�l�(D�����0�r:^CT
 	�I�p�y�&���( ^n�g�E��}����ջ�h5
��G�^�Y � 4��G.�K�ş�?�ӫ����S����;����<9�t��h��6�r�
-��ж�1:�s����y*׷(�o�jWf��`��r��7�ȡ���:t��U
�����e_"@��=F�m�O�?����k4|�"�v�mgø#>DNۢ��}�f�;C�>LN�Bw����_�A��K�W��l�H��vc����1�56�%�s�D%M���f�ly
�(O�#���k"LtCZN*?<O�+Ł0K	(8H%P/�z3�Q��\��`��~0�V�������g7��L��C��AB��@�\���.U �A[@�D%�65��ҍ��1A�g��%+�Q+^�/PU?Ot�OfhxbB�y��ج1��@Z����(�6!��!@irx��FKRtx ��T �!i�����;'s�n��DF-�(H��;K�8�6�V�0�c[�+� �W�>DO	�j��j0��.E#�6��ʌn��y���B�T�IDʩGM�%��QN	�I�	�iw�$l &Tz�f��!�J�t]�w4����K�e&�٧z.�r>&DUD̖�� W�);"\�D�j��2}�_���܏:�������.//?����h�����w���e
)B�nsk]@"O8V�FA��8\< � �� K�G�h�C��*P$����;��%����y8a(�N�~4��������i@ӯp�o��K/=z���g�N0�1�.���ӏ=&�o.̜�|.G+��4{�=���������L�]z�ғ�T/��S���Ca�������P<9�e 4:6�6�V�)�}��ҥ�c�C�M~����s|!V���s��t�_����N���0���;�m�J�[N&��-��m�Ѥ���@�S�T�I��Yr��m�)Q�uM�^�]���Y]��{=]�,8�e��)��)���Ws~�b���J�uw�cS���	A�'N��~��h�NL�
��&~C�S���jS�g\$UP�["I�H�F���5۔N�8�(����u���VC�SB<i� �/�
[A�M���d����Sh�fӨ�����~�\_Y����PZ�9p�L*&�"y@4k�H��gd`R-S�H�+�����l���R�n�8	���#�f��(����� 8V鯎'<q����OxH�]1p�FcB�O&�4�2�/-R ��@��q�A���)���l�~�]^���C?u���1@�ޢ��zB�G5BWAz-@�C�3�L�;�w�n�"����(�w��+Wf�����r�B��[^������6d�ёq��P�Z�M*܏������ڴ�����#%�8�SCv��VW�	�@^��	jb���=����顿9r����s~��+�11J>���������a�Ȳ������ر������!�u��7h$��Z��&Ŭ�=t��g.��^�t|�VK�-6���O!�J�7_����&vOS|8C6l�����r�J��q�Ӂ�u�D!��FF��t��өQ���thz7U6slx[t��$5�"a��yJ��R�'_&;�'f��*�k5���9!�G�V�)����XK*dD�N̉�)Ik>� >�V���C�ׅg0�ݎ� �P��.D*�r㱘T%� �4�acӢ��ړ?���T��9b���ҿ�Qd�6�&���9�|�@�n�C����(��s��
��h�E�QJ����uc�N�j�*����!�K$��b�g��y��kUjWk�I�E|1�1���,�&�l#"AK�)���n�<2/���Ǥ%��~�# ��ԝ�V�:�D}�W LCe� �Bd�S��� ���hxm(~��+�C�S)=%��)&	?W�*�A��Wi�vhn���I М�@��&�ۡ��P��hJ���]a�7�zK��x2%�2��d��&�����A��U=!��|,U�9�T���Z&5D�-���C����T+�d�A���㺅ɑ�g2��_���S^����t���������7���m��)~>�Te,�ǒۑ�R�  )����H�g0��pskK�x^����Q�� !>g��x�h3�K$Rs�����1��?6��W0�f���w�
}q|r��Z�J�)e��$��;oE��8�q�������]����Wh���M,;�	������	�J���*m~���+�k��#/��:ѡ4��*�<�Ii6�W�ΐ_(ҝ;w���-3h
3̨�7������|��v���9MK�-���4��� ȭ|�.��@iY�<�����KͦSd�d�RwW$N"��D���&]-΃H�+��H7O�4�NP>�����4 H�%� 
kk�����ɱ7xS�+�>�q+�˾��X{`��>P�CNŃ�%{֮*�wMs[��5q��G��!�.P��VD����ݭ*�`��A���աvS�U�^��Wb�E�
-���s�ݠ2/zဪZ3E�o��U��t�7�-s��mO�
޶�Ru��sT
�ᮎn[F��p�<E&'��aԱT� 0�B���Wr��BJD1��p�Z�����\}�-E�(���WE�l#x�"U�&�bIP�F�2��1�Ѳ �D�T�ϗ��̹K���.Տ�z�qb���ܐ>�@,	��D��@7R�E����S��x�H}!R`fR�:-�%���ȫ۷o�Ud�whpr�����2p����C�r��`0<�j5B�"  ����1�x-�{qqQ�G��+���j��4_� ��95���	���M%��
��[����l�����KH��4�7�'j~���t�]G�$߻�nZ�2�^B�N^� ݯ����С�hv��hr���{z?�w��8~���M��&Ȍv,Z��HŅe�L9���R1O��E�|��R����q'm..�^y�jw�A�Ω�Q�<���wӶ<H�Vh�P����$�T<�v��Cwn�W¥>O����aZ^]��c�侙��6��s���/BĮo��F�*�.2&p�T$[B�mxm�]��.w�-]�C<����!6���_�s��%�^狫[�333_��;Z4��0xڏ/n��(׆�-�ʼ�Wء����C}Q]��tM@�0$ऍ�b&XP[.��xApDE���#�$L_	����X���b��Ëv-��Td�Q+�)n�M�_R`�0��~K�5O%�6#��V:NMj�mG� G�y�� ��U�uK�M+(R~�i�����^j��'Ŗ���I�.��^KdԱ8�"^K���vG"�ғS/��B��I
e�(ʶJ��+.SG C�T�o�K��4�.��KfҔT�]&#�����h�׫���ڵK 	�Vȱ�N^�D#�N��cǎ��Tߵ_d��;�������ɇ���>� �î�Ce�B��W@��C����yI5�SJ<3U��b�!ׇ�]ALD�Lc`u�����þ}��~V�w���_��K����v-�KN4�v2h�8=���������[�~���=�S1���F�r�ξw���$��
R�X�ͭ2}�')�����>kU���SG����屮�� �7Q��4O���<�9�.����g?C�j���9K���R9O�/�#��NC<�]�!w��G�}��d��E3�kt�G/S���#O~�^}�u���ȦT(J��$5
%
"�S�AW ��*��;z�ފ�B����)��7_8J���⯴���`ŅjC����u�?e ���>K��ҹ�3�m��zy���gO�������M�\����_�������ʭG�
�ZUٷ@o��B8�oG\�V�趥TE��y�+�+M}y��:Ү����C�A!�۶Ւ-�CR<Dj��,ΒKA��Z�|s}���2�6ݖ%�N���T��%	���$~X
H�]��MG� |`� Rs��e*�\h���+EqE�V�:G��	6@D���KO R�T	 ���2º���YJ� \�&��d�����F�_���"7�ƸҸ���3`u����}��e
��k5�n�S�i4�~�^�lڭ�DY ��B�	�FH�"��%ctt�vFHP;u��f���4:�}�U�~ţ/m��_�z�G�|��\n�ߕ˕:^k$���Y8 ��FKKK���*�D"%�	����@s�[U�A����Ġ��>z���_@�/8��
ҕ+;���/��ֻ�����}��@Ȋe�P,H��0#�O|���V���_�r��-@l+����2}��ߥZ˓�?��lf�~���4}�Rl�^8?C��Q�~�]t�/�U����8]y�M����ɏ>M�7_�W^|������ΣGha���49T';�r�F��&�)�h<��;����3�ۼJ;'��x��|�Y�&��	F� ��r�"l����A1�#&6{D�F?�j�*E���TZJ;Ť樂N#_�Лm�������[+V(`Dۥ�����|����@�kkb�OV0�@���ѩr�:�)7���X*�?�ٲG����6c^�ynJe�
6Q�V�Њ����mI4B��l�ZRJ�Ȍ�m(\��	��k�tUnWG~:P����PʎHL��v*D�B��2��R����5����miAE2J�*�b��ѭy��
��4=���K��}ΙTP4��A�f�"��iQ�	p�ԝ�%���m)rA0:#��s��:4:������f�*�,}�_�T�!�����:bs:2�:D�ਢb�P|������h������7�F�.?�5�͈-EZ���o�m���#[M��{1��FF�_N&��~����;���[�k��.̔��GJ���Z�íVs;O 	�Q3ط6�uBꮿ�
�+"PR�jE[]WQ].1 �S�~��h���r8���>q���w��cO/,.f����^1,v4H�|_87#_��?�)!�];�2���v��t�^b0��hdlECQ��T
Eڹ� �F���ŭu���i��շO�z�Hé]{�$��1��S���-��W�Ny�㴰�IM�����S�ȡ�(R�ӵ�3���Bo��
=9>I�=���ht��/������V);9F���f�P]._������v��C@������`�@8�JS��S�U�M��W!v�
�����u�x���[oѥ��hmqI�PFUF���b�`�h�������iߏ_��>�R�=�ղ�eס
/�`@�sN��Dxj~�7d�Z}�RoG��G��J�����R��L� ��^��ߑ��ۛؒ.j*�+s�gO?Qnk��P����b_PB 4i[@��� �Rl�N�!�e)�o"�2����X�>]=��$uv��!�{ ~Җ�4�\.G��C"�I^K�,��ٲ����8�x��D�V5j����
�z��J��ƃ�$"L ��KH��9zf.����
��qKzI=ف��@�;��HHq�t�8��m�}m����ᑬ�(�%l[��_L����s��1^�.�������_X�X��b��v��h�^r�F��H$�ȑ#"���@�xO�2)Y��U�����_NLL���
4c �~���ǂ翿9��׿������Z�:,��+�`��_C��;'�&�^}�ua�q��F���{m����)�_zbh�.^��3oS�T��}�3t���T�(�hk�:�&�Q�ޤ��B�|�7Z�N��������|�S<i_��~��裟�$��~
�!,��tey�V�W(ēe��5z��FG>�ii�	Ӊ�,�U
��MM�`Еo��aCSa�t��i�vZO6(�z�]K��Z��&�b-�_h6 �=s|U-#�qW*8�B^B�;'��U����i��iZ���D8JIT���h����N'�Z���i�����4�q��^]���+��J�=��8��ty�T�9��'=)uT�6* �տ�-����q":b7�s@��V�#�MҨ�Ӗ�;��&S{2��j	�.��P����NԿ�����(ن{$`��b�:U�Sx��� �I��v�Q��^�+ ]I�RlF�H��+-%�ۄ�j���E�@jqlLZ�R�����s��z���3p�yH��ᲅ�JI=��:t��r�E�@˱�Iq��;|�� �;�֥�E~yu�ff�H�S[x8��:u��ܤe�3mW �y��-\@�i�6v��[�.E�|���ɤ��`�䯒��~��������Ͽ��Q�����g'� c��f��TjN$�IZ���8!%B�zh���f5���9���}��_Z�q ���@߸|~6U����/_����o=�x�ħF���)+D1�ۥ"�#�s��,��[���w�C{�w���*��hkc�<)�0��q���~��i�{����ŋ�Z���~�s��R9'��ŕej3@zi������C��S֭0�85;��`#���＋����!.\�LY�Aw�v��&��7���u�_rb��J:T.V�O�w^{M�W##���=)����o�<�i�
�R�u�PR,i�^�x_d�j���l\B��d,)<��O�닋B,�61A�ZC�Q�n�Rh�MI5�1�Z�=/�����u��������[�O�W�Gr��W� !x��9�xF�Igip"|���%</�/K�MB̆����>av�:~��v�j�6U�m޾+�a Kpz@����V����-
x�x)�4���iy]��:����z������J�	C��|�1M߿�L�Uކ�a;�qm\m���'ùT��Dyf��� %!U#*�\Ǔ�Cihn+�f����J%�Z*��,Sb���2 i��itU���w�|GPm �D%�����ҢD�|-u �h��0���VT_�I��`'Z�ۄ��gS<�G�FF�466"�7�) 0a��X�u|tt�+��������H&��W�֮���Y|ps-�@��:��e04�� ��H�)u{�T3���������855����~��7 M�c��s����cǟY�t���?����Xx����p��9
�*���)_ܢ��u��1Mw~�T)�)5��{��/��W^��_z�b�ϭ-S�]�-����k��m׶)��g�������Ju�6�H�e�	�ع�vO���z��SD�x�N��M&t��ߡ�����K�TA�i @O=����C�	��W����C�G�mr�F�Fs/��m����YZ+l�"�	R�]��kWic=O=�Z����!
���u�T���G>�(	TX�<zA���Yɱךti�4?~��IEJ�=��~S�=��Ĉ��Y!�J톻U,�;��Ñ���|�O�{�}��\z�1��R
��3��Om��T�Q��	_�\&�����j��r�����,/�-Q�P0 )+�^D��C�1n0�R�ڠzCj�<��,�oS���x&A��e�fa#\G>�HP//:]�����"u�H�dwE)�t����n�^TIHJ�b�KŜ�.3"�D|  �Ok-y�J��M�;OE��9W�z�5��F���t���1`b.Ɏ%����8'b!���u�󹹶��Gij|T"S��J�3�P�Y�E~e}��|�mIɅB*���ͮ 0��Z�WI!�� @���֨(C�X4���wK�z�{�n�&�H�ڠ�/J�+�w���###g�%�L�gh��u>��l�o����8Q(�����C��Z����+[�?/�Jnbb�9L+������2YZYY�.]�9��~�g��n%����υJ��:���S��_���,5[*-�)؄@Y��\�{?|?���܅d/�������}�������O���]�|�
[��0�X(D#�'�l��t���HU*e�Xk<��lȢ�T�:�⩳T���|�ԙ�Ny���Vi�'^u�2�(�Ӿ��'?6D�/�Q�\�k��х3�(�����F���+���BV�%�����o}��h���4��D�Klm*J4:2EN8LB�5��(%��B��I�i�%��8�NS�R�^V�y9�	�sk�Uz��W���Y5�&�ɔ�|�}`��J	ǼR�y����F������|��|�����a���_Հ�P�;W+��ߨ��Z�������t<,D��p|T����#* gۊ��Y�V�$iu�$oG�>�>��`5DY��Ϡ����D,vv�l��E>`�s(�� QK)�"��8���_�$<s�����*���T�=bDJ�Zq�,����j<$�]��3�,�SD���B�71([���}��3�<�cÅ��O�B�C���u�}m
��d�#�R:2>����_�D{�5�<sf�Jl-' �/*,N@s�z�Ǟ�]�V��P�Rx�ۃڣ������a�8!���~�iG����#߃ �+���8�333�0�����p�Z}��ҝ|M2|<^/VS��+���?�ݱc�/��t�����Tyeexce��co���[/�������ߎNM��Ah�믽H�<A=Lg�"�I	+�g��W)���2�@���.����t��2=��34����L��7M=�05�ഋ%�
�]�NW�����Y�
�<�:�2�d q�#�Q���s��N�9O��E���3{���F��z�lb����V���-�K���Y����7���V�'t��l�V̍<x��N�X^��J�HW���(�a�d%"t��#T���^.��;���
�����f�$�6,� �M[4�ІF7��!|�8�{iMZ]\���O�����~	v����3[���?�Uu�W�Us�E���c_������Y����~���c0n����Z����R�����=�j��6ݶ������Y�/���l��-��C�cxK�,!�T�%�嫴��B�ʍ�5�٦Z�!�n7:d�Q��K��i�e;N(Hq�I�J�� Q�_��V�-]%�n��P]�Q�����);���<vSs"]�I�DE��Q�����T�\-�)�ej`"E*6i�I���ۋ���
�V��p�Q��93Na9�h8��U�|�B�kN�i���{4!m�T"���Q�}����s���F28�i"}�Г�A�����'�,	�Q='Ⱦ�unth�o������ȿ��z|s|��;w�{�Je�뺻�����0��G�W=�&= �hm-v�;?�=����;�<��h&�(�;��C�:w�&&�B�{��i�Q����I����R9_�R�@5��^��w�c������h$�F�Z��/^��];�P�R�ĞAD���Kt��wi��y����<؛C%G~i�B�����Nљ�����<�s*��c6���[����yz�/���U���t�W(6<F���2�&O���v�ݔ:��
<1�{�*2�*-m��ǈ�I��(oTh�=$g�^&��K���\a����ŦtЮ�-��M>�������0f�����ڕYK����iB�$OG������mU�^�٬��gC�ȷ8��Ǐ�p��0��߈�t*O�k��7��P�Z��I7%j�.��e�x���;��~j�dm+����Srx�}��h��T��ꀚ?���΍���h�5^��A�R�:��@�;�?�*��D�Vw��i�utSU�Ŕ�"|�_-�Ҭ'��E��DJ뉴¶�+}���u���%N!����Ĺ"���SſJ/�Ow��(���'M;�䄅F��-֠?e���u[J���%iq
k�l+����"����qp@TeA G�0`���ynӍ�Mh�#�H_]�a�"&''��T)�$	��M����z6��\�ܡ_ˡ�O9<���v���:�ƃ&K���[�}~���'��?}����#��d����=��>O��ʌ���"��._�J>{^�Z��]�h���2�V��^����Q���#�����t����������8C���gi۾�TY���k�t��%�,�R��,%+m��P}c�
�˪+y�N.O�
�.���GSd�$��o|�R����ie~����;�#B4ϳ.���nP~y��U�@$��0D��sM>�0E����"��7�I��Uj�K��(�m;v3����+���;(62L3r^}�%r�=p���y��z
�!��H�F��PūI�;G֠�Uz3g�Ѕ3g���ձ8%�"3 �j|r���v�/�k^�^�5ͳ�d������'~����P�_k�}0�W1V���*ݛo��ŶM5�K-%mK�Dz�Kы�ߍ()1I�lW��mK�8 p^�^�rWs�H��h���1�+H�A. ��l��C �V�B��!B��)i��Q�X�}�ƨSoj*�R�$*;��I�%1���Mɿ-�o M���3�9�O�ǙO�*@.�i^lA��t�:�c��NxX$ �tDSE�aH�!��)��]�&@���ݡ��u�H )��i�勗�Pj�Ѹ|7��̯�VG�����z�kEpB�ώ�X�
���Q\NMM	)ZRz|ܞ&�7�Mlhhk�6q����}�Z��v����Ƃ&#JY���.���3+�����;*n+�mǸ�Ǯ]�H�wl�>� ]<y�6��7^���y	C{����^X��3�c�`rhH�U��$]�I����Oi�����d�R���A{o�GHVx{���|^4��w�4�@v�(�mǜd@��SOS�٢/�����>F�~�sTg���k�Љӧ���{�Wi��Շ�x���3?�!ͽ{���������O=�a���菿�_�����|�m�z�J��,,Ҿ�m�x}�N�{��|�q|�D�?D�J��ַ���1��ݔa����
���I�C����fЬ�� �M����3��mI���P&��󛘚�[;��jg�XX+7�ϻ��7?����G�e��`���&#�V��6%ˮM^�_*�@Nh�]տL�O��%�f���mR_���,�J� �$·4� pp��6
�;�&��!k�x�cΡ�� �ޠ���$j������+�_kB��Oh�]�(u�3*��u���tjJ	R�5
�jѢ�U%��+�m[���G�2 �$KiY����Z� ���\.W��	Aݖ4�y<�d<&�,�Ѐ��i5���2w�V�X$.doQw����Ɏ*"E�"����m�j�j�%Z�U��e�,m��=<�m�FS������H�\����[Y]�㍭�׷��O��͝���^A������ɿp!��Ʊg��9��/���Ό'
'�D���{���{'���E*��5�T��I䦺�'�6�����(ݾ�vz�A���,-^�Hݯ��7kvx����MNѿ}�)ٵ��ltV7�x҅�΃i��d?�����Qr\י����Y��o�*� A $@p)�Z!Q�%K���˧{|N���Ϝ�i��i�m�ۋ,��(���/"	� ��(��Bm��r�������*�ힶǲLI��TU!3##^�x�{�~���Gz|c������X����OKX&w�ٍ��t�-�������=� �C�"�I!�;`��:z���#oX�����q��	t@:����0��pBX�]�����^�ͱq��`lx�R;wo���u��p���:��׮������ ��>�vF>�]�󘞙����1zcD"Kv��f�UD�����l��/_)Ւ�x2�I]����oܽ�Ǜ��Yd������a���_����2]��u(_ѬE�6)4]�tU��Q�z���uhؒXL9�L1�q*-��E`���Q,=`�fZ�f�K���ɶ�X�Z��b� I� ��7�CG�6fn:����t����D:L`��o�L��tb�*����)f��X�i[ÔNh +%bPdi�&�k�S#��Q��7��!g��HPm�sDR�������Z�(�����)�[��M���>�bY�v`�=��8�T)+�4�j�o�btt���K�m�J��IngN��\Q�^i��!�e�d�*��9��/�~m|��tu�٭Ve����<��p&��{�8K&S'�ѥ7<�G���jq��w��M4���}�;���7o|�֙S���)ۀ݁�����	���=@O;��I��$�f�Id|�&��%��l���S�ٹe�hmڴ	�����!�֊�u���A4������"�8
��.�抦 �'�&|MA���C����c�0|�,&�n"���3琥;���A�Y��7�ɹy|�˿���.�ǯ�,��<i=��kb���qb����:v��PL����ſ��%2�Ə~��>���A�ij�]���><��C���¥��Q.��G0I;�N_��C���`O�p��4�G��M2A$�1|�|��܌���n�J]9�[��=.�~���T.S��D�J�nܵ��{yd��'��c���զ�s��|�h.�t]Վ����]RL�TX�L=5�?�8Z�h��%�&�����)*� *�)
�-ۏ(}$%`c�"�( @Tbq�ZE>�Ap�O�(Ȅgp6Ð�Gn�f�Đ�5�r�P�'$@��bx#�`g5��Y�fz�z��jԖ�Dܤ�M3L�3^����f���5�Ĕh���D�[t�Y��P��,ጉ*8��^��F�������?W����W��E�%���*��k��Y&����Ͽr�b��Q1�)��b��:=�&Nkr�!�[[�
8IJ**����DT�K�wq����Y�rd��MQ�ӻ��d�3�N�%�G���_NOO����)`����4��.�l{���#�/]��k���y��}�G=�]?�R���*����u�W���X�׋�o�ͳ�����^)��`��u�?�+���e	g����w�>�uy0�i����yq;�@zzy�M�Ϋ�9L7��BUv@�,�3c2ɴ��p� ?��Oc��8~�(�_8�g�2l~>�姱q�f��p�c��jnƓ�>L��".\��D:%�Wo��3�<�/�)�"�	�,��F1�����<�E�������x�������q߯}��} �[�X��s5�����A�hcO:��"'0��	���abd��7ŕ����ʶ��
фP�[��n��>���*t�.fS�d*u�P�=�~�W��'o>|����a����&ͨj�j2�5{ z�-��"k�9m�2L3"6~5,B$���*����6"!YS�*;m���Z6�EUG����r�e%J]U�Jq[�(�
�G�PN�[�� �q���:��)�M���6n��R:/:I�"6�!o]��3i��/���uzp4M[�71 ��
8�f��*�q�Ԧ��GC�ID0-�Y�V��f}8���aC��j�D�/���9�4����6����4�]V�.�u�����RU�@m,�!�I��'����r˱o��bbj�����'�Q;z��ߺ	�T�͐H�T7�a=c1ł59O������yc��L	Q���L���_�.	���\.��V-��c�_ͦ���d�ڵK/��8�[Z6|�%	~���
4����k�\�P(�����,���h?��g�9y���F.]zx�������:��ڻ;�:t���F���rg�}z[+�=�)�/�;��-�c׮�x����\���(��O���f޳��vx7o����F.��T:Iࡄx>�X&���.Qoomg�$����͡R*���։8��KW���������*�ݻ���w��e�P����;�p0���W�# v��=�����K/#O�s8-�8>�[�(�؂�m�p��(B�k4����>���
�s�ix�m��D���^�Q��pKWo YDO[3��4֭[�N��hK��G��G��U��ϝEgWd�ȶԟp`��V[O
��)�6�@O,�cS�b��кM�宻�|�k_+�������V�j[i��{{<r�r1�ƪ{4�B�hN��I+��ҿq�)/�U��4�q��PA��f��PB��ZC=�& �yE�;��Y���b�$�2M��j���"�l¦�Lz洟f�й)�7'���
˘d�#Ujʬf��S�l�bQ�4(�g�*��x�im) ��$�4�<�5!K���UZ��]��umE��)B�1��2%����T'E��᣹���Wu�-A�J��W���l4����b���+�����##��<�3'�IT�Pm��Y�5���:����My����ȼx<�lv�����撩�D�J�7�;�<N��ex�Xi�k��]�䵡Hd��L�p2��ñ��g6͙�p�?'���crr���>��c�o���y����7^|q��'���<1`��QGt&�������+�-k�^��'���#��(����ލ]�1�&P����P��������̩O�x��G��,.�|'O�FK�sKl?���&����c�n ���m,�cԳ6��������W�ͦ��8��awz��x��]Z�l{O',/��Զ���K�]Z@o{;��܎����;ￋ���we'�~�f�l]�t�� ��������ν���hi	�����׍d|�Ǯc*���͉�@t��z�e�����w	8]I.���8N\����<غ�7ĩ��G��m�}�1}�*N��왂%�maؼl�s��uЎ�ׯ!G@�B��70�L�d�f�O��s��;���o=q�]����ϯ��W�j��@п�ZJ�VS��u��V4+��ۺH}0��ʾsU���REDhq�J�����L���Z���4.@����C��/`KS�w*��=�a1��8�bK�*���Mn+��X^T���y$)�Dpe��@M�H�eY���O�������͒*�g�V$�R���F�`C�0�r::M��&T�Q1�4��dr��N�|��ʕ��n�lu�mb�ˠ��mL��j��I,k'-�� s����-��aW6Cg�b�WEI�,2�n+bf?�W�>�Uw
2���;��@�#\QњT�0��Z��*�-W��uW��|��!�x��.}L���2��R���F�����|��ׯ�޸q�OՎ��}lA�H`�57W����o�7>9���Ց�G�}'�ϗ4B��D$���us���oss����oNv��o����aw�5:r��l!�{�^��}�H�wii	���!�V��ݍ�z�7q��Ab1���߆�{��Lh=r�Z����`jqk6�c��e�׮���'N�ƍ�1lٶ]]hnk����͛�N�nuX�+��Lwv��IJ�Ɠ���ց�KE��~k��SG��N;�g�y��w�O}
�g�%���dC}=�§�����0�aH$���^�����ٿk��1��<y�SS8��s�U.aln�{����r��t6c��C>�F=W�*4Zҕ�oس��N�эy����-�L���>X�Nj���h$_���pz1nz����G?����D������ն��ǭ-�HkG�;s���D���`��ּ.���u8���i��!_��ȕ����aQj�5Qv�����V�Vv�t@�U٫�X"���3þf4G0�a�Tc~�����:M,\2_1�����QU$�wM#�rZ�f�tT��&���K��f��B���k�f�@C����2�P?�\Uuy������HM]��bS�|��x��E�I���4�ȴ	G�&�+b��>0L��gqЌ���W'31�տ�>�ў���P���0���s���qm+�Fc�
mTْ���#M̧b�e&�O��c~aV8m�K��^Ü7>J�ǋ�,���~�^���5#�I�\*�t$|p��3==����c�̑��%h�Ab�u�����ا_�#�ht��x�OB�я^@<GOW�7:3����~<���j���Kg�l=s�l���w�>����j��_E��M��C$��?܄<�Cܾ5����`qۃ-h�VQ˔�}Ro[�޽ގ.\[�F� ��}{qs��:q�9�h��}�Ql�{ cW�a|fV�Q�t�B�%t�����%�C�}1��	�f���i���E�i�ew���y��݁���x9q��a�W���p��p�,�����qt�C�|�$B'���Ž;v��ED�b���D�Ӆ��O���"_�Ѝ��Y�������w�h�9h3Q̏�`mK��9��
[7�rp?��z�#����3��G�&AS|"�Yb��J�X�]�V�u�C�>�+O_?r�H�O��m`,����j=�Vx;o\j���rKm"rHK���R�dZjX�v����&�,@��A�t^ח�78�� �&���hAg�r����vژ9E��L����jt�#X��N��4;�d��,�L�L6�kb ŉҍ�Jj�a�R}Y՚�\Uը�&A�nZ�@E��K=��:V,~���!�-S�a�~6��Q!�(B@G�bO�ƀNU�).%'];W:�E��4>fpX3+�L9�U�$j��L�C>srj���&A�T�6#S�@h�w�g���޸F]u(o�-�o�,̎1��9�43=�ťyML��Ƒ�L�$�%�/ �/��-����9;WЋªp��h��8	ܭ�V�k"����l������GGG�]�v��/#x�؁��Ȉ��?w���6:>~�X.5u���lׯ�@0����8s�b�<4Do�����?�o�:�ա��E+j%�oM'��a<��� ���.��t�Z1�|<��=�,�N"�xm4P]�Z�[1��xs�7oD3�K7n�܅$�(�-����cp�l p�#I`���w��̹�RE&do�1�(�EȠ�Z�"�oC� \��\3W������#�L)��`� I3Ξ;/�ן���)|����f|�W>�x�o�����C�v��BVn���ߏ��چr:#�Ʈ�FgO'�.�`���Gi�K�/BWsq�g�� L7T�z1O�p�j���t���4���!�;ɀ_��E�=�H0�*���NZ�p�}��o|#����6V�j[m����aX3	4Ӽ�Tʊ��+�%�Mb�v�L�BN�6x�8mu�U��5�RUEw�ae�)~���)�	/��f�MWN�1h*��Kq:�N,Ҽ�W�Qhu�Q�*�5��8"͈���rL
�M+�L2K�Ub�&K?��m�`�p�L�)`Ń�U��@<�,&ZZIT1)�P��:LB��j\Vf\��� ��P��W��`�5�D]��ƞzV����a̺���S�&�� ��Y�);I��].W���P(g���Q�(&�)>��r<�G�S[I;��0?�A�W�1�ilbR<<'��8����EGʤ��f
�I/�NE��h���v!�Ӧ�%%�*���)��hQ����^Z�ڣ�轹\��x<򃩩�ӽ���_&���4q:�ƅ�����#7o|�\��۸n�}~)�-.."�/`zf�DRU����X�V�[�ѱ[�dd[7�O��]�)��n
��G��o����z�D]A/օ���ʈ�����������pR6�_*c�΍�=�e��+�P-���#��]{����l��Fjj�0:��'`��=4��Q��V�i��,Ӡ�݌���Dv�V�6֒t=|�4	z��R)!$z��C_�xmm-ho��ȵl�=;�ƹ7���f9G�Í>?�7�.nݞ���߇��|9BD5��tC�N�y�BW�!�K�-a��i�Ȏܠ~�A3���N�Y&��ca�6����={
��I�t�"���dJ��?HǶ#U*�i��%�雺��������ݓC�?�*���V����� pyv�H2�Z��`q���0/F��uUFϤb�r��d�4�B\1��R���{�n ͌�T�_+�V��B(���Ų��!���ZJ���P
z��v ��M�U��]U�����/#S.��(�r�]��ҍ#M��ĥ�j5E�B�E�����0�c��?���Q����|�a�"������,ZC=\��X��ܟLeW�&&`2)3}������ƒMҙ�����8į����3�3iƚ�j�e}%fVG�פ����xӪU��]4��XX�"�QA<ڊ�Wߕ��	xK^U	
x=N!�3�e3a>����RMҾ���.G�V����_��r{���[�t����t��W�411|���:��o�����������������։�+>P�W�;`5�ź�.e117�/|]����9P��D}{mgZ;h���V��'P�HC��f��6Q�oZ�,�iB��0\vR��o�
;�,=� �K� Z��K�9/lJ �e�ۛ[`�cdh���C4�}H����`��	�W�c.��<����Q�dq���u�^8B~��p��]\+9��V�����@�?���><z�Ah�f�&�F�q����y�@8��ͫX�%�~�:�ٶ���t�}��q������y�D`M��
�w&���l%��h
\����a>���5��6�T��n/�����������|��?����J�^m���x��Bq[$��D"��2��E�ֶ0�b)虼R�:Uj˨	)�v/
Lq��j�$GE!�RUM���/�����FM-R��Dp�Y%�ĩ=o0�Z����\�L�� �Z�t����g\�g(�]��r�f�6��aF�t�X���w��QJ��K�S�R�΅?dh�*���k�E��6�#�!�j�*r:���&ӈ����+M;X�H���07�Q!�L-* #�s��dH�ԧ� ��ׄwT,U��Z1���=��
 ���A��6S	\�M��������R&��Y���jU�Uv�%���:��{�s�$���ŀ�v�(2�M�Y��KѪ`q��m���
�ң�X��/_~�
��E�x�M�~���/�/×�~���mnoi�ǣ\�~��3J@�������P3Fo�bnn!��lm-a�����S�(���gѺnk6�@y6�׾���8,t�hǖ�� O "�
��'�χBwg6nۈAڵ�,��`
�8ָ|hjn���+8G�6[�aǃ��tts��ʖi2I�����dK�TF�_@_G'�t�{��"1��d'oc~~�t�#���0�{5G��Btf� P�6nĽ��Q�t.+侹�E޻N��lV$��$n\�?��z@�oǦ&�A�*U�"I���"_(bdr
��<�;�}x~���iU��*A�>�� fT��Ү���_��*�T�j5��Ē�썺�ub��?����{�|2�;����V�j���7fҡ�X�D�4X�,zŨ`M[���&h��seQ�-�?�J�7buZD9���áˢ�zF6�E�n,r��BD慑�M��%*ũ:��XT�L� y�6
�p��BM�z�b*�C�@@gS m4��e�K��3<lnk��ǝ&�HR*'����
5�>8&"bKC�.�KM�)~������R&�3���4&hZ~V�k1��%�X�P�	�X�����W:O��fe�	h���.�T�	�c�;]��攍����Gr{<tL�T8[�XM%�>3�Z_v��(`Z��i����S�X���� ���qT���R���ة. �� �������<������K�*���yUqW��<����XbPh���w�O&7��
�����iӦ�/����hbͥW_}���W_�J:����jmvx<��[�0>z�x�&+�^���Z�;#~�29"R*�%^��ժ�r�ۆ�5!���z���������[o�p{AB��l~��ᛳF��঍ho�Aw�v�J}�lv'h4���>>�>m��G1_�!
!�Wx&��c>R�&�b��VK�nv���|���FD����� �P�N�fE8�Gdz[7@���S�ٝ۷�M;�a��ܜ�ن�m����s��/g�}�7|�<�_|�w���O}�,&3q��ݴ3���I��۶�N�*�/�=kp{|���\Nd�,0�׭(Z�(:�0­t�����t��GR�d�o��Ł��O<�؃3[�x"�]Zm��ӆ�~e"�`,W�tI�yS4y�a�y/��	�����.�"c� `"�Λ�.$o=�X��[��B��D��J�[�Y�t��t��7�ͺ"J��(�,�4�Yh>0�gmhK���n-D1´��fmD34������ص0h�*51�5� DӉ���3Z(c]CE~T�А(�$�4�8�'����T�fOꦚ��
��;Sv�^32ea�N�&�,1��I��S��˺PJ}�R,);�˚�Nq�&�	�����F��y�!�Yʆe�_M"{�J�G��Ua�uwF�Q��A#����IU߭T≾~}��Uȳ�J%z��y��z�0΀���e�t؅�V.�?�d-�s$<l4��H$���{�FGG/���~栉�r/��`��������ժ���vKssZ��N��!ܚ�ً�D�w)�F%��`af!.B��jV�J���6�GH��(t������Nh?[>��G�M֦0�a4��{h\�&�.,�R���8~�8��2IX��(^�wSV���4��>�0z�m Bn��A�.�G�¼�A���E�r�~� S$���<t����t���Mcvi�&�t�ɩ	�c�M�w�O�\%�I�[�aQ^I\i�7���-�ܺ�:�ݞ�[�5�S�p�7#��N_qO �d"=�G��WX�f���(�s�("���ٗ����� �\�j��L)��N[,�g6l����'�qQ���?Xm�m��t[=[��^J��m�X*�v�T��3�ƹ�hC(�l�0�nC�P��%)����I����R�j��5K*j��Ԓ�����9{e5�RBd��,��Ej�{$
�і�����ݢ*��:�;�J���h��.�1Oa�����6���s�Av��͉J�" G�LC�T�V�)�S���j(�/�ME������;�Lu���[���A��DgD�AW�%N��ue�lz�5�LԹ)�b�kcK*&Ls?��;���S�������qT�A�9�	�+�
h�L{�e}&�q��!� �@T�@EQ�4,�кy�ֆ�KE�^uu�{�Z�p��W���uIֳy�����@���`��ž�]��">{�LF��S�\i� Te/�����oG"���fS�Ξ=���������(���)hJNM�^y�{��=}����3�;�Π��У�˸{�.<x�~�ŏONɎ���򥤓qz$��ފ��
�ˊ�M��Ê���}�S�K�T��W��6�����^�x(�Srs�:1�{l�a��g�41%f��x���\Ӆ��[��,��h`�Ϗ|,I���{��ݟ��]��7�R�Fo�
��n�%]��v����iS$��Yl߶�>�
Y�LOa>��~�N��|�ߵ�K]����;�&@u��)l�D@��c-XK�'?~���;��^��s'Z��-[r���&�pu���x��ױs�:��wN��}�n���A7����	oktw B7O�R)G�b�zE���u�����{�l>r�����Xm�m��t�d2�'�'�-eâ��ht_��^�BܪT�A�xҐ+WբO_��r=g��@��)(6�5jv������b�j:^Q���aF.d��	8�Yb�����E����E��J�3��^PA��F��%��Gya�m�)��\�S#`U��@�3ȩ+�hK	��)�m�n�hfe�nV�A"@���+�9I�	Ph�~VRsⵧ4jfƞd�ˠ�+��pV��
�)� NJ"�A�R�~�>�����d�2�3��� T����]s:��M�u2�Ԩ:/3�WkD�ѥ�2}�4���eZ�Jj�e~]MK������`������[��r񨣱R(Va' ���N�A(�,�X���EW��]EU���q��iwh�@�V��ה˕�����x�8���n�::88�yO���@����;�x�_;���/gәu-����������s7�sf�'q��	�ݷ_���Ȗr�2rC��W.� �����Foo'-�	B~�g��������ٳ�����������Aj	J�լ���(�� \k{��A�?,R g/�̍k�lEyj[�zq��I!�ݵ�7������/�lj�3a��h�D��z֯G'�15%�h]����]�~,��A��DT�I?-�%D3i�!�<�%5��96*���@#��OON �8/�0ݘA�7�����A9����a�>71E%�����>}��{�v��2�����������iӂ8M�s٬+��b���7o��������O�5m�{�����( ����J5WEw!�����X����%]��&Ds�6��`a���Q��\A��G��G����灝�>;-к�D�T�5)��٤�q���&Zò���hJ���e��`��2#l�]aaGO6otG�MW�6��r�\�~m�����m���^-J:�ʕhX�38�`�C�H ���c����J��/]��RXtj,˚Lwڐ���e�#%��8O8M��(����uS��nڥ��P���L�����;L��`.�W��U��~�M���� ��~�(�ӐhD�Xˊ����L�um��N�����M�U7�t�a5���w�P��3W	5��3�I)EhB�O���|�@ #��,|�v=�|I:�#q5إ���K���A��s���z�֝��>S.vr��
�̳���+���?���v�t��Y���������I���)K�=]z��Z�:�]Ѻ50hwr}�*������p����/���!&gf��ڎ��v�<<p���\�Å`s��b�I1,��q��'�	0N �<�زm�f\�=BH�}�ܵZ���/�^E_g���.|�����/��܃�c'�4�����?8�k6���^�y3@*�J( �����>�sta��{���	�eG)����%������:���l���!�߃*��|��[7.a��n�W�_DO{'6�ۀ����qn�!�M��]��͊�6l��N\~���y�+���T�A�,_*�ĉ��,n�=�ӎ4Ewe<��,&�����\?�������%ʆ����V�j��kU�^/�k�rMbsz���6���m4g�	4)`ĕW�.�hѬ6Z�8�/B>A�6`�!ڔ���%a���W��R��7<��|��mM  ��u�<_1t��m0�P]]��M�4��E*��]>�h�Ȥ�Y�!Fsd8�A����奅9ϙD�q���V��D�t�2)��&�a�g+3��H�i
\-�EbE,���Q!IC�K�ʢd����r����)P���M H@� ":E�Ү	Ȉ҆�� 8�~�OKD� G����B�cY@����k�[���r���2.ՍM2=�����S������hZ�D��D�8�ȟ%ZTJ7����<�E�̜�������ȸ����k/���%>ӬX-��߯�J%'��B��;??�`�f}7��<O����#x�gM�]�z�j�o�y`x��b6�nz��u��nBOg��`��J0��(�޷� ff0|�*��b릍x��G�އ'j
#���@k��L fl~c7���"�)��oB��rmfiG��J�ji�Rv�]��%�nw?p����.�������a���������_�����qt�ۈ�Lq��X6��T;>�t�w +������>���,f&�16:�'�x�k�e��hR��0B�i��ņ/�$+�84���]p���yc��|ML!R8�v���{�c���&H}�M;N��;0��i�/�L!��cpYh��P�����EA�"�ւ��4�-��V[}.�'2�y������^_�q��G~�k����m����MsX*q��y̰�����r�H��r����~�׫Jǋ�X�ʕYF���U�dv�� @*W�ŻH��"��B^�"V� �R�H�f�e��(��.�e�z�(���X�M@���5��ӣ[L�JM@�n0���B�.�ª�}t]vŜ���b�d�@��^rzM��6M�YD��*�H6s�_�0���&F��cj�6xNfuL��FL�aD|'�jX�(�mM"Y6S�@3+��O�7S��N�&�$�^x҅�L&�o�QAv}�~b���>�>H�5�_�Ћ�Z �i����&�kX�U��A�.�G"S�O� ������ �C%�D���N���ȓ�M1hn���L��aA._���mx	4����4�X���r�ř�&��K�$ _6͕��.;���kؒ�凪�ǲY�w:��ˑH�&m�3�9i?u���"�h����_~���w���=��鰶����tw���A��ᴜ�v>�C�RY�nEx0��K/��L.�f��vmۊ�d�t
}�=�[0r�&������]�N��̏���I�ba�i4�H�s�^�΍��Y���?�ɋWhnqa���x�Q�Ȣ%) ��`G�<�ۻq�ӟ����P�GY�w� ���qt����M��.\f�*>�駰}�v�5-�ϊ+y����b���v��O>��Aj�I-/7���Y4�5��-������0qus��ܲs+�{;q��Q���˰�N�M��儫T�%��Y�r~vS�м^ĳ)d]yB�����7H���H�V^�s�t�V*_z+��yl�Ν�~uǎ�Ƒ�ն�V�ϴmoo�=;<�_�S��o�+�.XH�Fs����h�����׊l� ��2-XVN٭�f��H��Q��{�d�y��\��`犺�&�t�Z�^q��pz��>��U�
�\�_Q�il��!5�l���B�b.'�:!���h޳���P�;Q�� ���T�+�%:��vX��i���΀�mo�
pNSѡ�>L���a��e���
����T~�u�"��0f����$�YT�E��P\&�T��E�0�t:+&�4c��rŌ@9U�-�/�����.b�6$�#��)B��8*Ť�J��ꬸn�#zV[�����+�k3#V�2��t��O�����@�R)�Kt�O�yO�2u:�r�TZ�3�=��X����\e�x7m�+̳�摡��U�,c@�I@ ]��^��-�fdd�P(gbb�e��;�?����*h�/�z���M�N�����'�*���Ͷ�뇴��N�8Z�����.�9Ku���nF���L�	 |�n����>z333p��ްfH�EN�=��O���]c�7��s �~��{���km�k*�����-�J��o��##ױu�N,޸�o^�}��[Kϧp��	L�̃F �3Kx�՟�������?�������L��_��f�B�M��i�&��ਪ�ѩ'�o�^t��Cnc��3't5q��`�������; 11;���i\��}�a͆5�z��~�Eu�Hu�{z�n�!~�2a���+݀�B���[Z�jn���q�s�:,F1��,�SSI#�c{���=p�+��I�ȑگa�����/Վl�_xu4���Xbr|)��d��ͭ�|2�k����%�!
����.G38�S���H�9��9
Pg�i����ePq����N�V)�ar8W�U��*��|�ќ�H"��I��F �mW���� Ut�d����(S+Un:&[�� ��V��N�~O��%:�r��.%�p�|h3��s H��RΣV�Ӻ]�c�uy��CpǑ�f��T�N3|I�Aٶp[6!i��+�9!��̀�0RY/E���L��̍Z!����N	bҚļ ��2�Gn��D��,����d���&�KT'_Ns�ػO|�LqQ�e����3m�M�N��[��4^ը�q�{f��b�w� �rS�T�Iʏ��@�c�i1Hͼ�1�c�t{��%����� B?�n�d�JE���H`pb��A�]���V�F}��������O�X;�N�_M�Rp&>����Xsiz�F�����ϝ=�㋑=v����=���A�1G�����>�ѥ#	�r�U}{��ηJ��s�ׯaz|
;��"�����0�]F:����资~+4�^�HΘ-Kr4�rsq�X*�E?��֡��#cSط};ʅ2ݘUlش�Ο���qLǢ�d��>�=�V,D"x�'o���/����]*4ḽ�x;X���:]\z{��	�D���&�,���"��LB�effi�p�wM/lN��f|�+i'`�a���LO�F2����Q�������_�%�3�q��ͰCHM�l��;K���4ir�]�p�!�@7���� �9�H�t-,F�����p��������,���*V�j[m���Ps�]�x�y���b��L�3�f���|.���b�m*�м)�7��su6�t2)�$nZ�d��4��;�����6�p���׎��+"¢,��%��+��/�a��J�����b���L�� ��Via�L�i ��4��H�D��%��Ud��;�ؖ,��+� r�<2�"�\vt�y6Y	<�_+
X2j� �	i�I�b��)�r��N��WD(��R��Yr	����Gx@u��R�J�D������0(0�sD'�@�fS�9.d��d���V�Q�WDB�/��4�,���^<�(VBt��H�f�}4zT��EhZ�S�@ �� r� +�R�(�<�仯�/�y)�D2��1���$�$��pԉ?�Z�
Y��Q���μ.�S��阾j�zw<��I��H*�~�����.�����1k�d�4::�x�wv_:w��cccOԪ�5�����[�l�Ĩ;�֊��f�]nB�E�r9���îm�y������g��܉����m�lp��5�hw¡�MC롍�a>�J2�Ն��I4��hi�T.IL唙d]��ä�p|�1���0�0��ÆŅThgK�Q��K������I҆�����;�`ȇO<�8�{�a�:�90��r�Ϝ@�� >q�q�~��ב����$`g���\4��)�n8�)�i�c@p�D�J�2n���)�������'��\}�=|�O��?8�YחR��rh��2���䖫�P���G{s�m�	�:	���#�\=^ȧӥ�Bo�l?p���O|�֞={*Xm�m�}��aM��3�B�?u{��X4�ɥt�~��X�t6g݊T<�۴`9�>[Ze���8m:��xq$����i��în��Y$"���BqQ^�"������م㒠9�-:Z�����J�Z����ܡsZЮ�S��ݨ����_���������P�%H"QU�2�,�P�%׮x�l����М=9���E�Z�fz��tK��m�r2�Dˎ��T�ES�9%P���M��e�H�h7��@�rzo9�dQ!�R[M�9c�����V!pS�Y%����Z�%����Ze��ҙ,4)�#�J\���zN|j*�(�GS)��;%A�\ig���w���Z�@d#�|+��[}%���I+�����`�&ѱ�X��"9s��;*Һ�qL�Pd�晼���~�@/s�A�ƙR�gS�^[�T��_&�����}������1j�$�ĞqN�̥˗~=Y��t8}��� ����N��v�����@H1�sv�d�y7c�)>S�����(�;��������V��/^��/"[(��G��D
���B�n��c�P�g������a2�����]���^|�MLG#8s���q��*1>&�%�|�q�u`�p��uDg��F��^{G��;�d�9��D����Nn�@�F�P&�F=~�!�[�;u�&?��֢nA(�yz'��<�;�$��Kg��G�bd�l���Y��+����G���S�����y�L��`�����6enK�P��Qq{P$���<�J��[(���[^�������WԴ����ն�~ٚy�&��k�3�s7�^ZJ澜�򇼆֚�y-�B�D�L��Vh��xݢ��dp�h���x!������ps<.JY3I��^4s/m8��M�Z>�Bl)�b./�a;m>�;-�J*.���j9��\I��!��4���!�Б�	⅗ � ��Ȅ��hTJ���5Z�+*�
��.Qz�O��O]�J�����N�N���q`R�z#�gF�TDJ �ֈN5�Q���'e6EE�Ֆ��|�
�h���S�)=#Z+lL|'�Q!��)=��&���J�Gc�T,���;@��H)�XZE�(h�B��;=���cs%��b��R���E��ajQ)��̗^�M�l�6T��l�|�\!��̝�u8_,���R�%�pz^p��Tv-�s
�{J�b�Q��.--�����,>&������}�FF6����_��,ud����z{{�f��O�l]]]��hw��넲��Q��ĵ8���qangN��ｇ��9�6�0���勗зv ;�����Q|�{�����O~
�H��Eė��"����u
�s��%q�l���%���_�]AU�|{�vI�2���/d1;��/�vcώ��������o��_��j	��;� �.�)!�L�ȯ|[i`�����:���>�ڱ����.`av�c��{�R�W�I�Y�b������:x�Vtu��q��N{�>�F'�M��O�kv���A۫T��	�J��F;{0[K4m9��b��f��l~�p9�شk�sO��?9���%����ն�V��Oۣi����S��K����Ǟ��-�6���d��e�Hg�)�\�m�|43O&[�#C��^*J�����^6�bEU��0�PsA''�h�4Ӽ�Ϧ�N�%z��E��7��`/;N��m�_T��K�ԗ����+,��K<Wfe���q�@�8�e�9;��u:C��J�Y��F�n�t��%��E7�ϖCHB�V����,G�V"Rf��?�a���i@�Fz��I��`C�VVM�h���Z�"i�Ȃ���nA�yd5+*���p�ք[ėUa�++�9Y$"ƕij�\�V_M���ؖ�G@Q�N.�Y�)p�,E Uz�'XQQo��[�[��1�W҂����_��cf��-V�>�3��`n\Ss�WlR�r�����E��?M�bk#�kV���h4�o�O�������Q��/�ҥKgO�����O,.��r�4w0��0�v-\/�Tu�;�Мҗ �j���DU�y�ϝ��3�p��Y��It�w`ӆuhooE�^O�7o�z���v��8��^�����X/��0�|�[6�C��x2?��]��z:�Wn㶭�i���/ ���O�w��O�FjOO/��g��o~Q%�����c}G���/⍓bx~	E�����t��54u�16>����0}���w��nEkg7Z�;��s�R[ \}W���]�/����&
�� d>�󯿎W��&F�!��O��d�����VMH�6���l낍���Q+����,�k�T&�,��u㕾-[>|��G�L��b�������>�L�\��3�Sg�#wO�s�rj����͕��$�J�<���dNfp���S�Q��)�<���W�P�N����J\��\�����O;�L��`[���Tq��C�ϥ�l��G��H�\-�|�F8h�������'Xt������� )�
������4Y6�e1N�k�*26/�z4zFUɩ����vS�)if��P-�h@��6�XI��!��9f� 7&x7lQ��P��Ջ2�����Y���@]E�8�e�JH]$t�j��E�G�EAk�e�T�;'m�k�6��)�;@�@�� �so��+Ud�ϯ��ldDuQ�����\7ySXN
��U�R,)��M���j�*�bE��u�h�*B�>��.�V�\,4�r�#�`�}�ُCv���)�D�����O糹0�L֖�;wl��u�}wtJ��N�˥�r��C��f��ݸ�S38�4��{�3�b3�c��%��D2_0���nttw�RLL��ޅ����+�z��� �����Y\DKs k�X<��t.���5غs6n�.Bk���p��rsKqq�LZ$�ݶ,�'j�
����p�/�������t
)�QY]	)�XI�&���O"�\�]�9��o��ͩy���!�mߎΡ~�	8�a�B��-봢J���j5��ܭ1\y�}�}�'��v\����A�'ʡ�
���@�L���	N�8t��X,dR�=;�I�-��l޽�խ[7����/���V�j�k�2�Y�xkm4�����fc_rT�G��MM�h6��4����p�8����fw��{�{����)�X�Ϋ�\W���b����$ZC!��t���\&�mL����h�(��>�nl���92b�T4�2XZT��R�eQ�nC�	�R�t
no��T%'K���u��A�P�"F��@�@�T�!G�Hɱf�Pi˶#w
]
��L`c:�:�bn��>-g���W2�r�I3	�ʤo0Y�7�,�����! �(�(���Y�f���sTmv*�$���J�UVD0�L��M1M��iD�Q�e��9��4�ˀf��ZYyL�h�ߐ4�K�XL�U��L3,��%�u��/I�����q��wus:T����h��4O?5����z�%z������AS>mkj
���͛��v�zStqI[;؏~)͡ !JZ�Z�m
��#��p��و��#�+S\�^��ӧN�ʕ+�S�4�����uĄC�߇ �5�]����E������h�1z�&6nٌ�P �����*_F���T�C�>����ctbv1���	����x����M�$�������c1��N(��Ս�p+�tgO�Ca~Ί!J��t��휣u��װ�@��ĵ�q��8�s7��iܤ�^�>�ĵ����=�S	K)��hwfJ�ߋ�(��(
�K�NO��4G>�^}�]F�d~�&�&e�� ���D�e�����Xl�n�}g���?ܻg���#G
Xm�m��B�#J�p���˽����M,�~e6]��[��rՒ-��O!N�)�Ԃ�p|Mʹ��1�I	y��,mrY��&�k���4r9����Rh����#��\*I�ɢ���<n�J�Ѓ%
%��8��gL�� �0�%^(�\�g�H�q�JP�ƶ/N�9e��0b^��À�9c+f��+�5Mj�Uonjf�N ���*�����3�x��a�~��^6�Z+.�,JRᎾ��R�(\}��ݤr�G��4u��72�(G�jֺD���A�nF2y����& �_�ڄ����� '�
^�H��F�K��r���?W�q��fJp�L9M7�4M/@���޵  5�IDAT|��<��u�m�e�Ò��B6v��&�1��{���Z�~y���(�.U�UN�itnzt@n?G��XԷ�j�Cjw�u�6M|GGZ��M �%^����7���k(��f���M�9uϝ��¢�w[�:��o@T��Bi�G�!��Cr���?����d�߸�=��% ��[o�pۑaB"��9jj����i�v��9>�ҏq��e�>�8y�,ff����isHP��t=N'r���Rp�8|4I��itx�[l�7�MDi��97�.+���-%�����k���-��fށ���7\G��38v��Ma��+JIskz[�q��Ugf���N�w�����_�*�]b[w<�7%��r4xc4IŲ�J*_����޵k�۳w���~�+��ն�V�?o3��»�����o�-<<I}v)ol���D�f�9%YD>���fڠ2���mEZ�8�g���E�9ę�:-�N���A�Ls�t$&��l��E�dws�Dcb���{YP��m�/ �^��]"-����VI\@���I�ge�\��u��a�5�����w�nn]7��p!���bd�s�Re���roHW%����l]7A����Q�
��l�r�@����ҭI�">k6�.p���j�(��:!� �hM�n���i�]�y石�}���]j�����18��8N�I���)�����|I2��j*U3UY<�L����`�l����6ZR�z������}�sn� Nr��H���K��v��s��?�����x�\o*Qh�5m��t,�XW�L����NEL�aG��;�5��zn��w�>�ڱ�S���O��{�5F����,P�X�Q7�ؒoW#nnT��6�������q�uD�n*N��nC�/g����Q9B���[�t&�s��ɽ�T��tA׿IU�}�F]-�ZMlCKK�l>�+
�@GG�888����jK����q�x���7�Z��T(¥���k����K\@u1��;0��롳�	�X���i�D\���O���D�yv��`��-p��Sp��Y�w���۶o����)��3�<O��Gp�����7���^�~M\�7,�䰝��u�t�V��:7�l�}�g����S�Lн86
�l"��"Ԍ:?P�d�	��ѣ��&��m��p |�)����C/��®u�`�a�{@̤ؕXܼ����W����AGٚ��?�pG�ض��Ud�Gg��JŚ+���m�������C_�ڬ���'�S	��/�^w��zko\�^88�+=0�-�-hN��~Bl�_Y\�v.ÑJ�D�a?�r^�͇���9zƙ���b@�)1\��W�P�T!C��c�6~^/�* T�	ƀX8v~��*FC�" w�f�U�gފ�Y�.|QO(Ll(V�rN��N���}�΄P`���Ũ"�_-�_��[��+��.��HVs��E���V�2��c�9[�x��m�����
��߫��<]��K�jĨV��^��J���r˥�W���0A%cy
�t�nzW5q���jw!vݹ�H�׽&�#SPHbǴ��1���ܿ������Go���Z�γ"nt��cnPH9�[���l��`��i�G|�~�y���z�N��x���E��5'��\;�+��2��:��ŀ����c6�b�x�t�]/%�Wcϛwz����i:���P$�@7����3�Ln�d��h�oҴL޵�i�3gށ�Ǐ;�O�b>�XB�� ���J$!�HA,��V�p�O�;7�o�?9~���+���zŀ���ض}���Fa?|����,� v�ٕU�X?��2]��!(�Ws�xx�B0��>��n����	7v��^�Fv �,.B�T��TJ�ͯ�Af<E�`���Q���G �R��K�L���]{�?g`�T�{��f����흐��Kg�0ŭB���� H�( ��L0��l��kf!�X������]?޹g���]�f��ҿ#kJ� \
v~;}T��)�lt6���b�������8����jl�]HV���]�i>�#��iXkԑLs�Sc�Qe�5��*�~LvQ��֡���+�2�gҐI� 	���g�l!��C<z���L|��9�i'0t�`�G�G'T4���;�KLT�L���hʄ�3���|&E|_^}f���c�R�҅�����+�ʝ�e���^`�m�G[/~����"ݨ�\�`$� P ����l���%xu6<M��#��e�Iy+O~{S����eMLL�X��_/r�^����>��.�D/����\�Y3�����Z�P�E.j$G��%��j
^�dbۿ���=���
*�pM��7
��HDdAP��R�ln��x"�q�:W�qK�l�paW����{�:��L
=I���$]�6�!u�����c�{>ñV;�4�͟#MnZқ�'�<�#�����FM^�ߋl#�ľ��n�?�6��nޤ�J��T߼�v���"���_�)d��J�"�R)߶-[��!�L1��D[w�m�W�Ou�0d+cӂ�rN�<	�z�g,��0;;:�=�vJ����D�=��2�BQ�l넥l�R �g��e���h4�r|���o�f/�h�;���R����Q$��f�{��~Hu��F&bT&���-�N(�
LD�~���j����_:�:�RD�8��%87r�����+��]���98��a����.�ɶE(*{�=��A����r��P�M6l8�ȴ=s���Ǿ����"4gA�O``m������'ҳ�ό�j_X����l3�Wem
.�!K��f�vd@�[Pf�;'�/�-l/r�5�GPx�A�R���9�T0��]!���&Z�����/�qQ�cG�䆛�Z	4K�QY	B�-�82E`뀪� `����ȑ��of���m|Ϟ��;����U��j��`����^i
k�ܚ ��� {~��-�6��R�g�a�C�"DM��Sdύ��&��~>E�.���\`�����Z\\�Ζ�k��� ��~�<֌(��!x>Q��z;�
(���y���c�Fg���.�p�x=���ډ�Fu�)�'>��Pt2m^���;q�Ղq�aZ-��q�Y�v�-Í�5�8��r���v{%iM0�Bpc��6��W�m��R����fa�Ɵ[���՚0Ӫ�����^2)ا�;X�썍�ː�%��6��Ƹ�Yiv�\�r�9|��t�»���`G#e˖��-�����*�qvu��������:~h� S哠v�31>���7�|.\8gE����{v��۽7�I$�ͺ&�>}��O����o��ه�����![��+#r��Vs���k�u�T�bb"�%�h��v`�	�E�������S�Q��������?��?��Ϗ@(�ev�,&�R�p��9ф�MC���\����<��a����\���N���������Ad��Uv��U{�T��x!�������|�w���y�_��? � �V�j�Fvٙ��-�zzj��ѕ�ϭ�澸��م^ey�WV �h�D�R8�	kv>�����*�-��(�
����E��K���+�vnG�l��s��(iy^��z]|l�F�0�_�c]��%���ė��.
��ƶ�K���K��{���Uc_F���'�"�������/���fò�A�)~U��?�'�q�V��i-9�~Sx�wǴ���&���b�����Owv�<<8����t���2c���/�������#�1�.��^G����-��`a5�×YW���Ļ��ʇ��0�[^��������;�����u%יհ�_�ݵ�����C��f|F��-<#M[�R��{�y�IU�׆o��3��s�x��Ov������?
&�ơ� 6�#7�xO$�)J��p4�Twww�>�#8*l��ٷoXv�߬Z��JM:r�U�ԩ�Av se���)lݺU����$o}Ţq���Á���歑x�����Q���G^�So�s��a��rv��Qڱs��=�}�@��WU�%�R7S�"F�N�<o�q>���w���7���C���Č�����Fy3%~@P�d�e����pU�^6��l��2(�a��.$���$��A;�bє-_��Pء	U�7�ª�xgaڋнqmi����¹s��믂�W`���ɩhkoc�"J�6v�Ǩ5j����,�W��oݶw�Oz�m�>x��{��@�a��������ً����׮,�~k�Qo�|�n
P\Y�*v��R�i�������T���cCw�	�F�leU�1�Q��)�-��{��o�Ck�:��`W���G@����T�{Nӹ_.�a�u������Z��bJ���t��ssso�+�G����՚���X���}�J*/�VC!^o�hh��,�$�.�M�l�e��Ic�d�;[�����ø�G�:8S�Վ�s�ߨ�K_b"f{\����Fq��=���^K��l�W��]�a1���<qg�6}w~��4ǥ����/�8�Es�2�q��#T9Zu����Ew�����մ��Ό��KZk�X�/ʮ�ێ(���ncX���۶A��ۼY7�Lc��U��O3�4r=eU~�1*�`̳��%G�K�B��ٳ�;�O�����9�;:�h����u@,�p[�8����l��q��\x^}�8�w	�G�έ��Zڴ���Jo���73��]��jß������9a�����q���}�����O��ǰT*���=�$�9J��7BgW��">	ۏ�H�
���NL)oض�}�Q�+�o���`��y�����qG��P���U?F���
L�h� ���O��y~l�|��a��`׶��}h�������V���P*��M[��q��gi>A%���rm8�Ĵ3җn�����o�JJ���;�\]�\nr�*/�M[ܤ�d&>p�C|~*�"/A��e\��6&���V5�+�b��oU���6/x��oK����,()n�)�؉�^w����M�Cߵ�c��}5k��������7�y�+�B��Z������Ý7��!Q2y�E������8<�%y�\��`rUZ�d���'��� B�}9���\�9}��|���z��e۲6Y��Cr�]w�9�d��<I�?��l��Nq���U�����cD�p�߱��[��Kq@�0m���c�{5�9�[4븚��%��>�@lqWL�gv\�E�l�,gm
���B!`"	��y&�m\L~O��ko֜�������L�	��#~遽��՗�έ���Y?�Pua~��u���͛����?
	�?Qt������b{+n�F�
2ۈX0�t�e���c#��<�;v��m[����Q&�^$��o��V�]X�[���Gc�i���	�2	g�yv���9p&����X� �h��ƙ�����^^1���-Q��U�n��c����͛�����ݝ0:7�ǫ���1�`*:K+ D��¼v	]wMv ᜺g_9�J�R��!���5��{Y&޲V�6��8J&�ܴg�w�q�Ϸ�qG��)	��V<�+ԱN��������-e??Y(��ֻ>�_�-W��<W�\v	bLe�:!��_�R����!�E?��Y&�t��h�XD��|�/�8�QT?D>^�\�W��[�
�1wXp 砙e#e�o��%���?^��ԙ��	��{����[����"X�XzL7�ƒ���L�f��Y��lnrl�6-g1}�����ݩ��
���e��}cny�B���Z�~�c�;I�I��:o���j�qĵ�\ow���]���u�"	h%��q�%r�#p/$�/�Ĕ�չ@�-W�� jF{�ƨI�K��0	�b���D&�����h��L�o_n!!+^����SD>OE��cT�7��p�)���:�M����gW4�������w�=���UlkkcZ&@?&�H\����9N� U���R ��N��C�_��'OB}���`�MNo_!�J������7�r��k�Y&�����¶��u��m���~��w�СC������[�O�@Gw8� >[���B-� s�'�<"�p�8Zp�[5v�.V��i05;�^��N �bbǛ�����F871	g��a����T����d�'���qȄ"|ho[2ů\p����/j:�kc�R����gn���3��r˅��{IpgMA\S����+�����#�잋K_^���)�eS�]���
h��3�'`��*���Ν��AO:��g+n������/���"_ ��[��)��f;�JX6!��7FSO�w�&?��������r�ʩ�B��B�xs��x�2����B?�hkM�#�w��&�6'�������~�+���e^
9�Z�}�T�?S\Y��Z����Yq"L�x�ܰz!��$�)7�L�n9��8�;�W�f���V��\�-L�`��-x�v&Zoq� �����	���F��*\pnM�W�.�%��s/ޖy$֐�|�s2Lnn�]s���u^����`�G�*tL�=wh���B�W���k�>v3���QD��R�'��}�ʕ����B:��vtvg�ѰK��<�;dW�ͼ17�m;59	'���CG^�+WF�N& �@�wyhh�d����A�"�gW�p��0��'*�ehxc����瞅���C�i�&���`~~�;�c-�!���^+�":S��DCn��cl��DL�]�PP� S�K��@Y�A�/1v0Fk5���!�#�� ��AM���&<��z�}L����]coMלR�a�Ɯ-^�tӶ﮿������E���8�!sl�z��x��pgv�����-��;W1S���(��xB�4����@�0� �j�����PҬ��*/x�} ���kUy7��r�!,Z��2�:;;U3��<������0-�]dѪ������0W��Q����l����qI�%���t�PVT�t<�������>����9�Ğ���6�bq�n&,��E{EA���������δ��:`�-n���=��#�\�'WX� \�	V>�ΫMr�:QpI\d��a�<��f͂튢��7 �Yk�*�`���������b1�}����ׄ��o�E�<5���f����P�G���:�#M^�+cccg�t��w����PUw�z�AGw{�m�VC�T(���#���G��ɷa9��[�w��۶m3����@8�g�������������w+�F���_ݰck�~Y���ކS�[n��vX���g4�f*��x�G�#�$~�ٕ��>��ׯgɂ���@2ؕV�/���K�����o����剉+Peq�ov����`�w4�W[����>!�p����-?ںs�K}t��A�^�	�3/� ��|i�x߻�K]ɗ�`�[��FJ�%�CО�A�P��b��)�D_� z�`�.M7@�� �Ӱ����ͅ�@�hU **�x�7uD����gQ.�����=z�l4>Wo��6c�e�~�fL�]���d{����m;-�ݽׂ������O�j֋�j�K�F�L��d�#�:�NX��4G���EY-o�/x�L�t����^���+b�I�@��BoY��^�h���3���f�� ��yMnṰ�z&�������뜣l�E�%�n�����G����_"5{-�HD�}Ж�nH��}�����r�Ϲ�jc�����Sp��7`r|��w��{��CO�F(|;������3����o=��sF�f�*7���u㑛��U-I�������f�ɀ
2�,5*c/�ʄ�Qg|I� ۑm��F�`y�ҷvtA[:�3SP���0!�
,��z�:�ݹ�	Xa'
�=I&�����	��0?���"����%[�w���Ԟ��v�����֭�]�� �[�'O8��=��#����\|t��o\�t��.͒	s�,�Kaعq��`��i��8�����ϼF�f���<��)!�� �@�'��yw*x�W���������R��L�\��FH�}�`8p�/IS7n��*.h���������ј?R.�V��v�N˲�f��=^HWl�'�ӌ85���!W�X^��Y�O�$���n�IB�s�u�F��ݹx����k�P<y��r֌;���ڼ=���(��B�@��p�{w7���^�R<{�z�x?�hz?���<�6�lk�eJr@�$�X���S���K/�;�΀Ķq:���;w��͛,��+$�����M���D�9M�0�V�R/#�m���ק�ܡ���!�o�����<�<�ه�M�d	�8@0���0��+U�?��(�J
���*>���Y����<h(�d���� �bap�)�h�0�>��sˋv�֨ɪzi`�����{֯�#� ��=�����:��lg��ř�GǗ���c�$�S��<LNNB@� �	�]��V�󺚐�x�%��X�v#�ڏ�B��#X�X&������G�kO���Ľݘ��q��o��V������������\�7�P��0�n&(dUT��#y�����kj�]�#�H�(�5��:�-K�f�4�`��O�Vá��,	;
��nM����4,�*� w���V���F�X���$�q�4�>Y�7P�{�z 8�ױq�5MuvY1ʶ�2���W.^��;v����l�7�|����[���ؓ�L��tz��*|��B�T����i*�sǶ-
�*PU�0}�m��sj�;L7$��ep5�5�:�����&���vb��=Jʹ,w�1���X,�vrHuwBM�!�nH�$���L��k�9��T�m{�k��s{o���m�w]���;:� n(nI	x
<���ɋ��g/Ng�4bUo�"��l�	�t� ��@�`_Da�0[�ׇ��N��ԝi���
[Ѭ��t"t��*U�^j�u���g�NM՗�{���o5��M�:�P	��Ќ6���_��iH�L��ܸ��[´�íP��� ����y����ټ����iF��h�5ŴPD��$n"�6������~��(��W)��^��
&[��+�P�Ɏ��Y���֢ɮ��:�6n���:q�8LOM1E�6l�`���7C�Ћ=}o��i�̯�'��iG�w�^Ku%�;�o��P.F�l�J��#��t�r�w�X���}�>AZeh�:T�� �C�V�S,4	K�x]V��D�}8���"C���e��˹�e��?<���}��2������eA��'A�ؠx��h2zj]��{dz�	�p���,��299sK����I�e�rbI[u}x�Ҙ`�2!�D�',W�۟��H�'ym٥K�������]�>�~�����"���Y�
��|��9 ��B�7='�)"5�E���.a����<��Ǩ �T�r�B	�SΧ���(����h8½���p�)w��P��O��RG����k-���_ZZ�*�L
���x'[0t��ۧ���f������֋�R�(�20��v�3#W�UC��D&K�
�{n�rRh�?�A�R���AE�Z��bEU��X�^�3�F��.5�9�Dw77{s~��$(05�/V��r�Q��K���o��y�O������M�"o� >Ax��hS�8���L셑�هgK��.ה�r�.`W����T
:�)DS FtvC�=�,��uNՆ��׆:���y��~�4�5[�~422�r���t�V��i��{;��h�)4�J�z%7}&5c�����r~7{t�Qx�aY`Ȧg�ď_uSg&��6�j.���-�4����ر��C/	��)L�9�ɍD1��[o`STB� ئ�_�,�'c��wٱr]v�]�5M����ېeF�Qg�Ν����T&�z2�=�i��ר3������l�xwBR~ۧ���_{�z�<�H��ހ(H����A  C�L<�
�5&�0����{v0�X*��OW$��5��Rɖʧ�m�ݴg�O���{����A�'Ϧ`�ݞx�X|qv�p��|�k��͋u3=_�)�SUX.W�=��t8�pD4@�eقZf���@G�:�+@��x�,��|dd�h�R��R*}�0����R�$q���A����s����i4g�6�wȹ���t=$��n�<���P�������%a)��l,"7�=��'r�C����sFBA�EB|�/F�|8��2��h�^H$������1�<�$��9@?����q|b�Z.�/������o��X!-7ZLOO���|qC:����Tn��}�4�0��!��*�6�2�� D�������z,��H�9��y�,��r�:,.�T�k��m����s��m�=z�m�}��"Ač��X���p(�83�T�k��xxd>w�L��5*07�CE�C=�t(I_�Pջb�c�Ɏ��o�M�6���y�ҥK#�j�X���Ѝ�m��@�'ITV�����fmS���闈�XXP�.�"F���p��ç�%Z �������`>r��Q��&���֬�*�>.�LC�F��7��2#�
�^��,�\4���a������?P���{6�L�����Ją��sְ���u}�r��M��}�C�]^��s�\5�WAg"��h���W�Sa")�����h-���!>-zba�)յ"��8���������A|���FCF�x�Z���џI<zq>����٢��8��<�@L�����Md���;rݶ�_�x�����'BWbo��+w�����4m�(XaUU��������[��=�u�q#t��/���v���m�,��v���qn w�=�p�+�G�@F{^�nD;���A�O�b���������4�;�,v���[9��Vt�O���/k��K��m�����wUX���aH|=��50 ��.�ba�1ȳ��n��n/O�4V�Y&��oٽ������2]!A����e�il �|��r������6���peyJZ,Z�~�PR�}U�&�Ͱ0����{��r���ժ��a��v�N��n��U@s�������Y8�����P�<�bI6X��ǲX|����7��d����TQe0�·w����TT���D:�s�v�ES�kQ��*1!��m���P�����~E��vՊ��SO�Y�@ww7�A0����@�l@I!o���r�8��񇢯���o���S;n�m�>�A�2�x:����}o�#|�����酅!�0�~�[����4�����Q��r��P�ڸ{�eY&v��Ap���ءX�
���<yf�6�Xs�~N�Syܛ���������U�S�H�>���LK�L�hZ�A>O�?��,�įL4}�t�"��L�/�`#Z��}qY���6z.r<�Xk�ܨAղ!�vr����l~T
��sϾ�n�s����K�A����ό;Υ��ؓS��6G3�m1������F�s����?�l��z�|G�T�����E���"�u�	n��'v�T�͛G���Fa2z4)�y5n��-�i:O�Z)��Y����z�G�$E�
�S�����g@���M(t��5_���Vm_�������� SL��*���j[P�4s&WX��_ߴ妿ޱ���~�Bi8� �Ϡ �H��F\C������ϟ��#/U*����=�D�>��%�M���	;�lὢ�G�l/�$xi<��d��<v��� r�w]��g���W�cb��6מ�=����D⇙L�7�ф�
B��8?�W��LQ��Eǉk�04l
�ӕ�S,K�Z��X�������G~g��Aq#Ҝk�8����#/�*�/��&�6��\�&7�W	����ݼ��Ȁ�sw	l�5��c]�Θő)�q/�W����e�����'��S%��@^mo�Ǣ��Z�-~�Bp�T�J�d,��S�d�n޽�[�;�M��W� � nd�4�����7s�ܩ|>�^�	�M�(�0���*�&	�5Ms�M���:�݂p}�$�5��>IígB�q�m��0&�� SdǱ�\0�a,�<|���|�D�7�w,	��(f�L\�c�P�����{^ؿ���]7��A���������J���b���Z��9˲�E	�\;Lۡk�{j���9��x�%����9���w���~���"�/$�����S'���m�u��é�����={n��G� ��0xk zc;q���p8��j�a]�a�m���,����\(�OSs�w_3
����H��?����y)���͛�n�f�O�hj�+�@A�B�`����������r��L��P�A�U�F��@�F���#K��rMP!���L��L4�F��o���h�r��S-�� �XM۽111q9�;R�׿j�=�g�fj�j�N���89kv������e�~����^����9$�� �hf_�0������r��j������d�'.���E��E��wW͹[K�i�^�ϴe�p o>�h"� b�fg����ߎF��r��=�Z��iބ�	��y���F�V�����M����������X��h"� �1<<�9�sNU��R�t���~?N��pJ[����6�׫m�"�(�gR����?��	�H4A��"Du&�N_�p�,�O����L<= ��s�:m�	I�$8��`�7���	'?������&� � �U<���x��Sf���-+���MNQ	)wo޽�I�.]�&� � >���8G�(��}s��)fO�� � ����Dz�[�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA����e!�3ۭ�    IEND�B`�PK
     �8�ZIRP4#  4#  /   images/2dd92824-eee5-446a-82e5-cb3be823b6e8.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  "�IDATx��|�\u��sڜ3}gf{�%��)	����Ԡ~p�ދ, �
��(!�BIB ��Mv�7�����v���=�w�z�+��_���7�)g������<�sfy�I� �dq�I� �dq�I� �dq�I� �dq�I� �dq�I� �dq�I�
˲�ҽB7�'�)4�z��8h���h`�^_^ �r�,�0�W� �a"��Q*�T�P�A ��`��`�j!������dt�'�	����˂�➃�<���iy|���ލ�gWc�`M-�J�� v�(�Y��@2o��!�	H(�V��PNT�� S.L��g|/�2N����</
�������Z��"<�`�	X���Ï=�=�gq���zOn��}�s9\~�%8i��3�Q$������
����q�T�)0�b*�%.Κ�}Xn1����7U���j"i)(@�\P��:4�@�L��*̠�T�E>�A6�ʦ�����[������o�E��p��	�5O��n�x�8uA&su@�LADi����4��>!���t�
*:�Z�O��yp��	$�
!��A�9$�#��b:�Д�F���w8�����dduJ:���X��-��=c�(������פ�n<�د���+.�d���E�1D�Ĳ�o���Z��
/�k��L�?��	�БS�&@WUDr*�s|DޭA/��2vGdԻ,ԺM�T��TT;,x�M�t��@�$ ����Օ������ˆ���`u�s� &su@\<��#c���/�S5��:2&G��@��"�f0��Q�`A\��HZ��kr���>����a�N�e蚰{"Ϲ*���%9:R�l�ˁ�X
�Ơ�D�̅�`�R}�]�Lo(G&/��r��9<���͙��_،�I�&>�w�ʣ�^G���L��v�霪���'&@Z1Q��L�����#N���)�M��`Zh�t�ԧch`��78�HIa��_wka�+ۥ�"�v�3C�HƛM�%3BR[�g	�� m�stKo��'�f4TW_��O����m�w=�����9���1�����H��R3�~��x��X�qx��b2,4"gZ#j_��!�SM�C`t*"鈋Ayu9
,�[x�<	�!FtB��s|�o��3�}z��@�N_����q'2��<�$�'%�XO�n^9ݷodtV2�]�f��-K����|Ak�5����è-�+����y/�We�?�?�3x,�:�}w����r}��f�\~[*��yp4�t��Dږ� 3�S��0�xe,��I�\r�pTE�Ü��Z	�w� g�H��i��Di!	�u����c�Xy�Ixe�zl��5C��Y�ֳ���m$�J.�]�;����%����;��{�e.��oܣz/H����F�A��[�ˈX�y+.��M�hy+.n��_�����m.����J��$G�'�;SV5�����,��2���@d��JK�0q��'U7�G�� K��{یR߇�|��U���t��с�_[���Q���De���%��3C#i���Y#����݌}�Xg��0�����_�5�W!P�dEOm�rݙ��74rʓU���W�B����x}�H���j��zu@�ne���[x��=?�ҖnI��j���"A����NF��'u��qh0��.It#L�]����.z���mI��S[:ֻ����toL��s�W4�'�s
�|������=�˃Ґ����=���7iKiX���7]��J�#�UeQ�4��:9��$<�/��ό��kI�u%���O�c�w<�Q+�؃�ּ�^r�{Z������9:�BBþ���馬Z�4����ȧN����\򎡉�	R@	��P���� F�)$��n���b �Dy��2�:���u�m�|��`�7���}��\��X���GM�)��SrL(���z�s���'�<��K��-��q� J�8�L�G��"%Գ�NddQu�/˰�K�5㒅�}M��3��{�:��u�>�������6��H�{+����������|�1�ۑ�Dc��qxKܨ(u! @��� �Y#	U/$�mpT�dt�\֓V�Er�����ܗ�-(�|k!�̧FmQ��{˛�~�m��Hj��X�����q�Ny�3ܭCޟ�A5L�/(�R��\c�Y��3�xh�����3t�0��F"�ҽ����8����V���O>K<��=��"��r�Y6���Þ��p4{k8�s�g��A"#y� rJ��t�$��Q�Yh�W�3��t���Z�EU�Q˄FvJ}�ƹ�PN.����2�����h(�:��8�͇�N>V���S�=�x���w��$J�v���N�<l�+��Հ.�C{!���$����9��>&�����(VM��Tjca1>2��s���_ǒw%��K�)�/�U1�~Z<� �:�����
7/�[�PB��n%�^#]1�L�
ޓ,0��?�3�ݤ^�s}kK���Ԟ�]��=��� J���h}�K��<�O�Y�q��^=�9\��U�������ɈFc�F�Ƕ�K��xY7������p@��Cդ4���.9ov��=�k��Y1�ǱD�ߒ��9�\����@�#���](���0K���˓�7p �G��%��!_�P�w�$���`�?�\%�ӳ�.�l���w���Xg���Ι��~p��5��B�읊�^�.����0�%�H��4�ϣ�g�B��m$4�s�����\9�EI�BW(++{�k1) �C��#�w|"_t�}x&���5��[u��?��j��浳Cw��"�#���A�� ��QU*$�d�wQˢ��<�亳$��Đ���z]5%�>��D�������������ފW�V�+�W�x��|&���r1�E�� ��VL�ƇgWsuᚐ��f:[�����76`�֭X�|��Z�I����U�� �*��짖�h[L[�j}����4t��*�%"�UB V��H��WX�i�&X,���#��Y��´�{ƒ��F._����gK��̂�,�ד�HO;X+�4:�%�y����r$'��Ff���T%��k��:k�bQp�'9ş�Tw.��9�9)1I�$�y$��*�E�1�уh2��tF����P��"��kO�f`4���(-�)�E�����22��,8�XT��4RY�%	�"�,�q	c���^3Q���^0��*O;6O���:`/�Eզ�~O�l�Vu��!���i��)�S<�_�I��w;�IH�L�f;wF!�v�&�Z"�©�G{ǒ7�Gs'f2���𸩅8���6Gn�-�o��9��hdA��uj7�en��E8�A()C�%E���G ϒ�� #�3�4���:���CEUr.z�����I>��W�AkѢ��4��DkH��;B��PrXN$�S^���ػ}��w��p@��\� �WB<�# X"g��JCW��]���Ss2�kr�����,�k4�\Nݕ˦���?}�Y��n�j%���w�f�j&�e��S�J����D�ֱ7�F)�;�`�[B2�����*��N� oW�YT�p��R���uH�D �N��%gR��`U;1�&���I�-T�����f�`7*ʚ�y�fTVV�������QDU�,�� `Y�O_J�$E2�*��`$I���(f�#�W9%��H$uA.���ȥ�$�<���렬4�D*�)�K���5�<�շ駝v5�!��Q��vɺ�����?��V0�+˼���
t����]��[�ǜ� ���ޅs���'�!9J$NN>-���J�*�[N�0 0�>78j�&U���0XXn���5���j��lЪ�{<�t9�����!�7��ׯ��o����f����������W5j�)��~��NR�d�h��@
e]�`���O��i^�F��sT]��i:���.����"B�ȅ|,_�N��?���[��qх�@"��W��ϛ���42��tg����F3�چr�����.[1�i��u{����?��vo� �V�x�ڈ�q�(Lx�����D����BK$�H*S��wr0L�EK��/]r	&�"�o_F��"%����y�I�4x���HtJߝ�</�Q��nہ��~���D���HV�yB��HN��������T�;�ύ��'?9�}�E�d�F��	�,�E�}� e�y{]U�\F���5�D꧳-8����oa�'.Y�p��Q[�����UL�>	��L�;�!������[���R+���������24�^��_��ZYxE���^|�Gm�%�ەBbB#�ch�e!7*�"�>��;�����()G]M�������v�$���/	=�iJN7L�����Ub��E�����m)������4͸زG&#�N�Vf�X���U�������Sr{�8�s(T���U4�h��@l�p��ң���/�M�V
2:ۉI�CA,���?����[�/�PI�G����o�꼏�Cwgө��*Zv��3b03��w�"�K3����)AXJ6����Ir���Ŗe��0z�2�}����<dy�x�xH�UcU���w=�$Iߩ�i|���S-�*6mڈ��{�?@lt��V�|��b�o�Q((G��e��������a����EI@6���
p88�d�9���D"���o=��U��> �ptˇښ fNm�{�?����h4��M�9<�'�8������vO�I=P���8: ���gK/�*�I�/��o,�{/A�14�2�co��@	�7B
�w����8q���c��hA,����>RQ�<Us{�ս�Ӣ����~�z�͟��{���[~Z�
�����I��k�3�4�i~��K--�d:��E��bb"�M�2�'��^uũo��~.Z�����!�y*��;/��b�~<��pAC�ґ3؊Ό�i$�,������a��J�%y��#���@!`�J�w���y���+]�m���u{Ƥ��1uZ+�|b�������1���(�uÚ�I��7^�,�ݹ|��m� V_d�����d%�1�*^6j�a�7�ۊ��ppzQzv����O(r�e���*!��ɗ��*hn��E矌�;$N���������9S"�`s��Ry%UJ7��D��A�k�h#�K���F	������8����c/b�q���1�9�g�=�h�\�����o�PW%���0}�]i�8-�KN�k�����C�܏�o�M_���h&[ .H�*qS��ϛ��*e�]Q5P���:R�e�1��I�U݉����*k����8Z�fW���b���Q}U��6ރ�� &��9	��\��)rwv�b�4�ve��a�������L�}�1�ކ���N�I@c]-j�1>6�*2�S�1:E��.���v������������W�<��C���|��|����I�߁�U���'����UEV!/��y���v���b�(ҩ�&�~�kxh�{�<'"��.]���58���� (aٯ��ҷz0/�����F!O-+����X>����c��){Nvu/R��Q]I��!_۹s�)�R���Ŵ�&H���*S4�\.���.�Ҍh,��D��mhn��[�or9��=buu����g���k�i�Ʋ��e�ʝq���q����"�H�Vg��*�`�"�T*I�)^�KyE��<D��~�ǘ�o첮��"|�}8�u�¸����z����~������&P�$=��1����3�	�aX��n���~�>�o���T��Okȓ��A�0�]A ��赲�����j^�L%�H&~[T�R��0�a�4�����߳y�]b
d�7���?��g�y��}���3O?�P�&��%ߑm�chB� "�&o�WZ�T&�8e����M�\,�5���n���mw;N:�C� b��47�iOL��J������^ WD�,���%��AJ%Ppo�Ҋ)��0�g
�D֚��z���#��y�f�I��J�M$�\_�Sz<�L�Vpp�����/P�5��\�GC�	�r����8����ûvw����ܐ���:�?�֜w.��&����ƢV��m�T��otIն��#Q�@Y3��^��
-�ݭ\��]��vC#ueQ%��зk7y���];�
<���7\�]�*� bg/	�g�<�]��'��L Q�g)��Iu��y"e�������mU��nLP����K8�U�<)32��)��!�&jAUU�Q�Y�ڟ������x���jj���{nJ�sW�bji�ڹs�.\�eK�% k�n���h�����}&b8c�|4�z2u����������,ǯ~��/}ܲ��%TUC�1c�sA�遻4�����8:^y]�Uy��w� ��gg֣��	T��x|������_��>��fh5J$�^Dɘ&bh!�[tA���N�*����8���ωN�����tw	B^����'x�{�`�^�p���Mo���j�,^���v�������>E)���ս#ڠ�."��G@��Y����m���ڴ����zOҹ~�w����_�r�cfE-�qsP�d!JB!,]~2�5�gb�.	�������Det=�xg<��E�9|?�	���j���v�e��[��7E�j�REˑ�fPᤊ�j���b�;ؿQ1��Ѐ`�6�;-R[��ji~VC�ZϞ�=�b�E��s��mI���h>_��z�q���~y�f��w_Q&��EX���	⦉!j�y�w��~�@���xq���J��B�dOZ��/~t�x�3�Q�9���ͯ"��Be�/]�����vuCaET� ��#��o�
ɧ�C��7��ڢ��'������G�~�.(��Vq�w���/�@�#��ЮT���������Lߝ��A>#��ؙ�0���%���6���#{�=bnuRV>7�2~������M	𺩂(����y�Uj�f�6�h=���߽��v�����Y�҇�����AJ̇��Z466��1�;wnǴ9�G
j�WK.\����>�١���D�$*��xW͝s�<ںsZ��ލ��W@W�v�Gcp���Y}ɴijX;"��=�'n��<3\q�Gp�'?�G׭��<�1g�N�\k\"��;G~2~v-p.?�'z��f�B�H#�tu�\���ܒ	��r&G�ɢ���L���y�xF����sC�qLki\��\����*9�o=��;6\��LD"1Fޖ�n�fa^x�g���C'�l��(�"a��x	�{}��r�͠i�4P9�M��8#PO���Ķ'֠�Z^���=?|kq_�Vy�l����*���e����'�<�T���4�񒥕��5��yf�:Q̔Q� ��v!CSD���Y|L���2��A���R�����ϙ�(���p��Y2Ɗ�OC�<��ر����1���憆�/��W�*�y�I��ς����<�<�3oj:���}�nhy��w!*����AW|O���THe�/�=8��7q��Ӑ�/�ߺ	��^����_[�q]�R���xx�9̝?��u��s�G�}��7����]��[��xZˎ���뎜�8e�Z�h6�ڠSJ��К�duk�Tn�Ù�5C����-0BQ�S���x���$�r�R����
GH�3HS��U��*�����v �0������dXz�b�9Іꪘ�:��������ի��k�6��݇��t���R޹Z�|�;֏�Sp�j�ǐ�1�8�o�,���?��ޏ�,=N���S�{�!�z�%~p�4L���x�s��[����;f�|��ύ��/�,��2ev���K*�Z`7u�=�`�m�D�~�`?��
�:X~�'��Lu���}T-�{$�R���UE���h4�D:_���B�c_2d�u��� �r���{�"�y������؏�T%���vm}j͓dJ�/0����s����N�l�|�8��VVP_V�)��%9ǽ�,-]s}_������@ޣn�\����b�ƍ��t��u| W�u �	<���W�?��/�	�;4���"#X���	F⦏.ǯ�o<`0�M���88&UP���g��_yy��X�s��#��բ�]\YV*�%H�d��I2�|��E_VJ8�[KC������[�N��P?,�Ħ76�-��}����k�{${�]w!��@v���]���x;�d���}����gל�ƀv�x����sq�>�O�n�[Q4��������Zi$5��;�ژ��Q�毞����m.�p8R�Q��̢�2C������Q�!c)J��M׮r0����p���.�P�0
j*Hk��n.��~�O�ɇ���*�޺�FD�Fq���c��wvka��b�����D���!~�ٗ�C��^52/�}HY�c�|��W�#'\��Eո�����H�wbv����t�BN��,w9�A\eq����'p�}}��_����2L�R���P����?&�%�}��*�M	�}���w�!�q4�e�UŌ�cޢ��Pd�߇�U�(����}���	�?���'u��cY�0;i���cI=���(�T9"�[��t���ݻ� ޾��v4�b�(��L�f�e=�:gR�3g�{�?��ZMmY%R瞏<I�����ǣ&T��S�ɻ���X�w��ٳ���iooG&���t���6���Q�����mW�q���eQ����^�_��|�1o޼���}��E᠊!��T<���F̟��O��ï\�W�Y�f���d��1@&Yd��1@&Yd��1@&Yd��1@&Yd��1@&Y�?�͕�UP��    IEND�B`�PK
     �8�Z�&�y`  y`  /   images/8c2f1315-cf23-4ba8-a920-becb97f13280.png�PNG

   IHDR  �  �   ��ߊ  NiCCPicc  (�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D�0գ ����d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c�%��V��h���ʢ��G`(�*x�%��(�30����s 8,�� Ě�30������n���~��@�\;b��'v$%�����)-����r�H�@=��i�F`yF'�{��Vc``����w�������w1P��y !e��?C    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs  %  %IR$�   tIME�WxG  �zTXtRaw profile type icc  8��S[n�0��)z^�8~$R��b;^eWݪ��HQb�0$|�>�� D�h`�dZ@�&F�Ąb�9��m��P=Eec������O8��`��Й�f�
�Q�A:���{�xt�k��7�����������-eP/���\!�����jS�u�mۃ��Qa;��B�["�,FدCl֤�	�����/�&�S�T�c��\���~�y�_���D6:J&�D�z����f5u�R�����Ye:�010�����?1:9�����{��5nH����^υZ�w�R��WU(5G�Ӫu2j�fo�-���)�:&c*+q�y&�"J��G��|/��d�c?&s&]����VG��^q���@����줁/0�   orNTϢw�  [5IDATx���w|e���3[�����!�XQ�	6�g׻��;�ӟ�SO�]�Slxީ��)6Գ��^C��m7����cӳ��؅|ޯ����y����S�y """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""�P �t뎇yX��s*�+��������L����>����<�r�ݵ/�ϯj>��ߌ�	�\51�;Z�w�e[�L�>��( ��R�	�NUo��W{��v��	댍
�_�f�|����Io[����7�9	s� W�>����&A����@��H��t@U���"^ n@U���^}z/[�j�[�*)9����n͚?VTV����� �*�, 4 ��{!��yLDDtX2�I�+�|���5]�dݸy����S�NMX�˯����^!"Z�SNDDDው�]8|�+LUU�S�
�n�u=&҉"""�����]bc�L������H'����ZND��fK�<�M��DDD p�ݚf���*(w��CDDD��%�$ϷX��'0���������p��a���ʓ<���#������	E��Qn������iӶ/[�lBaaAV�`�Դ48��vX�6�-fh�	�R�4J)(�L�O""":t��r�];���T�r:��'O�����z��:<7<O�����F�ۍ��*����v����"�_A��jf"��r�|��������Z�����=v�m����X5z4LZx�Ͱ�����QCrTAii)~[�+¹1k���e�E���;���^�&���� ""��:Z،m�tV��r�}^_��✕Nx�^�m�H�Q�6�5�_�6���At�z�^{�7].��#�WDDD������[u�ޤ�r9�q{"�F"""j����"b�-��t:]p{8�Q��JJK��x��.��o�\.x<,�E9�

�i*^=x@w��NDD��VPX �������}U�z<p�\�N'5C++)���r��~S�7}>*++#�F"""j� n��&"M����|��`@'""�f
�����D����>�,�E5AM	��������r��t:���(4��r� Ȉx>�N�3҉$""�������3ƌm��.�x��N%�������/ �y9�9Q���M������NDD�4 PJٍ�������(��@([�6t �z}0z������h 4��^�����(�i�ee����h�����(�iK�-W*D@�1�E=m����R�b� �Љ�����_�� t�"A��#""����+ �ϡ�ʝ��(�VZV��H�*w/D�H'����B�*�˕@LFx}>��NDD��VQY�D�Y�NDD����
��q@���;Q��*]N��!��%t�t""�h%М��J�u�h_u�8>�FDD��9�����_g/w""�h�UU���S�����G:�DDDdD��j5���~?K�DDDQK ��p�tݯCg�;Q4�b��b�W]t�)���(�i�����]��:QT�L���]ס�|
���(�i��LP�0��܉������2�fJ�r'""�j�)(���ua�;Q��bR
!:�܉���� �DD���ʝ��(�iգ�i0�OM�r'""�v͖�u]X�NDD��u*��^]B��܉����V=u��-�p`""��&uݸ�΁e������h~����*w""�����z���*w""��%���u%Ͷ���NDD�4�߯A� �+�C�)���(�i�߯��ϡE9i��5v�#""�~���J`\�.�NqDDD�N��	�)NNDD��l6[�����DDDQ�l65�`@oW�3[j^���&��Q ""#f��dX�~0�d������%سgv�؅��TTT������PJ�n�!11�������dt���D��@��!"�:��i!K�pr�V��"((,Ěu��ӏ?a�����ۊ����^�'��P�Q�4M�f��EJj*�w�#�c���5j��2a�4v":�(���fM�̡2N �ro!���b�ڵ���O���o�v�Z@��hI��� �z������ck�f,��������ӦM������b6��'�#�P\Z
�łX�#��9|Ĭ�BV�C�ϡ�I��x�d�R�=�m|�ɧض5��Q��V����TT�c�o��t����o�����_���{�]-��O7���������Wa�QG��f���x�� ��ZM�mݶ/�y�y��صk'�5�촭ܚ��-�7���Ǘ�č�wfL����/ 6j���m؀_|	�����xp�e�F:i�10�\�˄� ��n|��x�����Ͽ���"�U�&-��]��ۢ_񧫯��͛q�5� 1>�A����PXT�w�{���?�r�
��Gjj:T���d�B�*w�U����r�~�<��S((؏�L�Z���jVb��d�ɤA�4�������!�/�fK!��PX���gݏ��"�|�M蔖ƠNDQ������3�������rV�u!�a���|�8������x����sꝌ0�@n�� 33]�vEnn.�v���D���#&&�*������ �6m�m�6��
?Ȫ�ବ��g�����w/:��3�Q�Q �-[���x6oڈ��/��̀�B����F�}��nǿ��:�^�O�@�edfb�ر�:u
Ǝ���,$$$�j6n�p��(..ƪի��O�����c���5&������ks�"�S:��v8�vu"�:%�%ؿ?����p�Y X�6��҉G}���u��g��Ĥd�:}:���J�1	qq��6�|o�n�!+#Y�p�	���+0g��{�-��0�{=x���w�޸䒋�)~Y�(�(@)��ۋ �D��*wv������չs1�9�s��Q�����s�>��;	qquü����e�&3��G~�>�,r��G]{c
�Ņx���p�B��u ���B��.|l����7��ByY	�s�f2a���x��p��� !>�EA܈ ���p��31���2tx��jؼi#�{�y�UTD:눈�Q  ����]�*w���������];���t9M3��s��3�>��C��K ��f]O���z]�u�qI��g��o�e)�����.��8"�����ޚ��.@m$�q�L��Y�݋�99�3� �8�d���<1P(.*�K/����Bu"�#�D�5����EX�n^|�%���^��c�!�u�,������,7i.��bL�6-d������H��!!DBv3L�ڱK����[�0��<66�˵1l�!{LL $'&��+�D��0*�������?���9�te�:��}8��)R��ys$���~P`��f����+ ;v��']��(�O�<g�uVD��;f��8��S���/5M�����? /o+���m��������z�v���z f�6�V�f��v���G��4x?����|�=p{�����X,�Z��Y�0�L����zo��v��vCD`��`�X`�Xj�o��
��p������v�����������
Ku��6���������vC=��f��6��+_�Q�ן9p����z���`2�`�Xa�Ya�X`�~\���,=F�S�3: ������]�����f�ߚydMi��7"�^@��U�_�V�Z�S+1)_r1R����& 118k�x���QR\��H.5Kh8p� V�\�n�f��}{�b��X�n6oڄ�{������j�"..�ѣ����!''16[�>����rTVV6���dBJr2̍���/,Ě5k�d�lX��w�Fee%|>lV���е[W���#F�@�~����Т������k�d��[�{���鄈��p >>9�9:|��>�{#.6���T^Q�����u��vj����dX-���+*.����d�R�[�;w�Dee%�^o���ƢKv6r��b�0` R��[�6���k׮��ŋ�n�:�ڵ�������|��CVV6C�A߾}���|iN�M� (-+�֭[�v�Z�[�۷oGA~>\UU�z�0�͈�ۑ����]����4p z�쁄��v�ٯ��BIii��RHLH�#&&h^Wy<عs'V�\�իVa˖-�?�W�~�V�������Fnn.�����#==�6/Z���N���w�Ʉ��"��_]�QPX�������M�w8HHH`MBCR�C�r�ϡ+ e��OPU�Q�|���8��qM�Q�0t�|��(�!.>���ӷ/��!C�b�ر�r�]\R�_~]�O?�?��3�mۆ��2��kf�b��%;cǎ��iSq��ǣszzuN���:^y�U��ƛ��PA�Ν�ēO�wϞJ8�v��ǟ|�w�}�V�DaaQ��P0���ԩF�9
^x!N9eb��pj��{�|��gx�w�b�
VO��SV��;w±��/��=��9�Σw�}s^x���"���D<���Z�DFM��8����s���;X�t)
��k���43R��0b�\p��6m*R���-��������罍%K��� ��x;�iiiw�Ѹ���a' 1!�uU�G[�m���_�/���e�q����\}�j��l�Թ3����S�`ҤSЭk�6��*����#f�{����T�Z����o���hpL�UU���_���a���c�8++�)�dAJr2�)S�bƌ��ۧL��>��~̞�>��chZu�Q@iI	����$)�����nGBBB���u]�̙3q���T�� 6�M3�y)���7����DDV�Z%�{��~��i��Vy⩧#�?~]�9/�,g�s������g�Ɇ�����\��{Ӷ��p:�O>���8S��S덑�Ο��T����䤓O���������9�~�����������EV�ZU�Ϊ*y���O�-���XgBb�\vŕ�a㦠i�r{��O?�'�$�Vn'5-]���u�c��V��?�4_�R�����+���RN�<Ebbb[��������s�=_��\ix.y|>���2����kU�$&%˥�_!6mn���{��ǟ��#F��jk��^w�[m12�����?�)

DD�_�jm��x�z�.���9/6ȓ�k��5��t�Y/]-���"�ǞxR��燝��W.�����_8�9���Z<^o�cġ��������W�$&&�Đaß�L����y#�+R���_��ax�euɑ��GE���n�t��oi�t���߸Q�t�%%-�A<�">1I.��R� ~@��_��[��A�dw���V��H~a��q�ݒ�֩Z�~e�&�,�W�j��""%ee���K猬�������-r��dͺu�:���w�(ej���4��O?զ��G�̬�6c%���c�ʏ���$_*�Ny��$�k�6oGi&9a�I�h�v;�}~�|�ͷ2q�d�Z�m<v�C{L��v�Y���E��5�|s޼ꛮ���ify�ŗD�����s5zL�s�m�`���9�] �6l+�=^�\z��횏W]�'��}��|������?Q������UW�)DfBN>e�E]���b�����o����
���ߖ� �9J>��3���%��^�F��W]]�d�%��N�m;vH������n�#��n~�9���d߁�KG���Y�����n�Y���z��q�v���|)���{�%	���S&O����IgU��0�E�V�V.� ��<΁�,���x}�V�Y$t@����""��[�k���u��)S��漼f�π~hzBb��'���) ���X�|E��4�5
I���3\8�o+]�	���j����h�2�>�'PJ�j��j�C�����߭²%���k����~��#L{�R
%�������˯�����뽤�>5�9�K�����|�p&�y��g�tVɳ�o磏>ċ/�����������O<�gf?ge�i�k�O_Kҫ���O=�J�n��=�O<��#(+-#���?�v���k<��l���V���³�<�[n�۷�ե�����Vs�����f��>��Ar���5����Ǜo��nǲ�O?���|vl�Z�/�Ϥ���`�5T�����<���t����ԍe�7z�����c��
�Z.ս�Us1��d^}���طo���v���T����	۟17�p#�6oBM�4���cࠁ9r��� %%�����{����e˰r�J�߿��3X�sN��my����a��q�駵S/V�߇���:�x����n>�c��ХK6z��.�]�*W�����u�VT��:F*�~/��70}�t�\�
�̞�*���vLGl<r��W�^HOOG||<\.v�؉u��a���՝Ϥ�qW������8���o{GB����x�w�rU6�?&�YY��ݻr�� !!n�شi�l1�	@M�2����8��3P\\�G~�����=Ɓ��������HLH�����]��~�z�ܱ>��4źߋyo��̙31n�Q-��χ�^~�f݇Ғ"��:�q�ӧ/F��A�!5-q��p�\(,,D^^.\�u�֡���^fԧa��������O?��G�^�+��+V��9/4� p��!;�z�쉴�t$&&����@����!o�����=�7?�}�]L�>S&�2=�z���Q��i��z�oټ~_��ٌ�}� !>�i�8�ѣG�ꎀTK <d�ˡ�ܭ�yu�kQW�|�_""��J�R�� ��]��E�qy#"�l�
>rt3U=��N��?]#��^�
���Kc~]���b��_�o7��dee7S=	�?`����/-�[�*wM�[u�w���b���㏑'gϖ�+WIqI��=��|��z���R6m�,�ϙ#Æ�Y�e2Yd��iҳw�F���O��N?S�xk�lشY�+*l���T/]&��q���t�?&�U~��v�r�+P��0_Lf��5Z|�Y�t�KU��V�\��m�����2n�1�4S��*M�Lr�Ie����|Qu�㈓I������%kׯ�����RZ^.+V��Y�= �z�}�(��|�m���Z|ο�����_�?q����k�u��r�%��'���?�DN;��z�����������q��R&INN���uHjZ'9��d������������|�t�d�Ν��G˹�/�	I�^�:�).-5L�_MP����{���={e���7ߒ��� �TIrr�����o���g�����҈_'U��_­rOHZ��C��2�[��ʫs����楗_��fx"6\v��uD午HQq��w��m<�����O?�J���bj�""UOu��)�e����8M���v��
����j����Y��n�^�{<�>Էd�r9���͗���ӷ����\)*.iv;^�O���2h�Аy3ᤓ���(�1
���%1)E���FٴeK���˺d��[��$�kwyj�3�?���|��|���d̸�C�ˈQ�e���a狈���;��ԴN��{�!���m�\�����By��g�i�V2��0��)bЛSM4�E�?a�|��gRVQ��^RV&/��buڍ:�)霑)?���;��_~)���Azjj�|���I(��VFe@4x����^y��d`mF����;���I��������W_{Mb�/�J3ɔi�ʪ�k[��""�����s����Dd�G{\���N��E(K^z�U��x������V��s�ꐡ�F�7�~>��|�駒��E�j��v�!�W�{��z]�$����O>U{�nz��Xz����Ss���ǟ��脻��� =z�6؎�������~{��*�\w��B��Kv��2�5qU��[r�麼�����|�8y�ŗZ�
��,\��?ʖ�[�F���뺼��[ҩ�q����Ly��k�9�u>~u������8�����C-�˴��T]�;ŉ�����:nt��	�6�m��{�⥗^FeE�&��0�$<���n� �z����>���f���
��}6nl�����o���a�X��p���>}zXKgfu�=��N8����:e�D�v�ü)(����[�-W �l�⪫��UW���E�2b�p�}��P���>�)�����1c���Z0@� 8��8�����PRR�6��>�ſ�ݷ߁H��i�Ĥ�~���a�Z[tk�z1)�3�8<� :gd��5E���ܹs�s׮��Li�y�L�ݤQ�^����:�L\r�%PZ�c�������QYY����tPi����,p�W����LJr2,Cf����,]�zZ������v+���ݦ�5;��~+����k׮Ň~�E('�|.��RX�ՊI�&!>>�B���p�e�a�)���ՊSN����S�*T���eK{tcǍ��W�16[���I�p�ĉHMKCs=��=�\�}��V.��a�ē���t;^��7o�?���U�|�-�޽��wM3���/�%_sn<�	�g�v���
��֠��t�̟�em�ӑ��7�x:��55�%i�Z,8��sеk�n�桰��]RM��iF�]�H������^�Fb�#��eYE>��C��A߷Xm�����;���_#G��u�]�#�.c�ߋO>����k��� .>]t�SS[�@VV�/�:�v놙3ς�ln�vrs�"-=x��u?���ۜ#5�b����.@���V��O�>�޽[�|t��s�;���k �ٳ'��2�#(..��o�͛7�/�2X�����_	GLL���V��^z	�`�tw��~�	J��ڥ��4Κ9�n�q�>}0d�P��K��Q^V����@4MӚ-��,�+ >�����餶�>o޼K/1XBG߾}q�9g7���-���N��#G���5�VW����_�~?��6�%=-�YY!�9���ѿ�6m'%9ii��RQQVI4�|�ޣ;&L8�MkINJBN׮!�3f���)�@bB:w�l�LEE�z�!�����m��tn2Yp���!77�ݚ�@�=0��i�M���8�&��֩SgL�2fMk�Ͱ �����`�[e����+���n�t́et�������v�M�h�"�ݻ���5�<q"zT�õ�ѹ3N�~�aUdYY~���v	^�G�F�N��Plv;:g�يѣG���>�ݎ��$�������|�0�aÆ!��s`�X���a���0rԨ�Y�ZC!0�_rrJ�|q���1�� 2?��#��`������ĉk�@m/&MÄ	�����7������Ö�����>�+jJ�k׮0����|>����5���DS��b��9}��d��zz�`D�6�Jm�>�-[fp�$��`ʔɭjwn�0q����%���t,Y�eeem*i��V4���`2�[=�i��JHH@�v���b� 6�a����m��3�L8hP��6[B�4����h�a�Á�i�@����.��y�73���}��r�*���>}z�)�F��h���<X��o��xڼ�A�!11��n�SRS`���	H?����%���xU��HE�{ȥ������
@iY6n�h��]�tA�~�Z�w��}���m�6��o�1z����j�����$''#�Kv۷c���tٶ2��j��w�^mi�v�a����ѭ[ז��`;m팚��{��Q�����Ў��� �d�\ߴiS�o^�2�W�ۯ1..��fXD���F��@��r�4MCL��4�i��RXX��;w�߳WO����l����ܾF���cZ;w�j�V���;����iƗ۸��fn��N��:m�v:��m�-�)���X8���(_��~õ%/�e���f�w�.��c��{�n0��ٻg/���߆���vdfd�9��X���ۤ@��TbVJi!�H��J)$��#T�����6�5�G�����W��Ē����؃�̽�d�`2Yj'f���҉��m�F|\<�����q8���9 �)�@�MHH8��c�=D3V������m[�3���Lطw��vA�� JKK���ڪPR\��6m�j�"9%�]�n6��B��v�8m��T�w��)�.���Lf�����t�x��hTPPgee��Lf3����Ih�tɂ�b����$
~���-�;b�i�bs����j|��������l�Z�'���<��~ط��MK�^�O<�8fϞ��-Q�݆�U�ۍ�¶t����G����6��A%f���n ''6�.��N���p:�H	��pQVVVݩ��~
L��z ����d[Uմ)C�u������j6[`1�@��:%��c2���RZ��mP <^o�APD�(5M����P\ܶAZ4�`��5��2�B���9�+ ddd">DUdQQ
�x'-�n�a�f2��#�Q݋�)A��m�Ř�&�ڱ�Б�d2�|�^�V^OscL ����+8]U����J)��C7k��nGm��f�~�m� ������xRTT���o�]�K�1w�*@����]v����9�`>��M碦��E�p�iLGؘ
���>x=��E�"At�vxl�:i��;�q��;���O߾�FGZ�fmTݙn����+QT\]��(Tk���_�W����Y��Pe{�T�����zЎ���@�����G��e�h~������.���?�Ƞ���ʕ+�t���=�����SO>�?���r1l�0�9@NN`2��f����_�QYQ����r��	>8��4�cbjg�"j��M���x���;�<s�O6�f2�K�.�%:�����r��G:��� �>qqq�(����+�}�h���ښ�����_�k�v�ڵ�|���t��@��}0b��u֙8jԨ&�)���i@��������"�t�������QS�z���1��!+���s_������f�s�7� $�znC���#'�+֭]��]Î۱h�t X�~=���P����ʅ���}[�[���郣F�j�ل��m6Tx=h�Ș�������������mSi�Z?8P=�Պ�x�N�U.bc�پ��&�D-��U�!���`����wW�������rE�u֯��n�w().F「�1�2220|����OMI5|F���b���}�m;vT�����l6dtj��̨c3��HO7��N���E����$�/��f[:n@ v��'MBl\��f�-X�e˗G,�
��m��駟AĨ3�`��a�ݫW�w�;�W�����P�t���ׇ���A׃����S�N=/��g�n�6S���;w�t2�ZLucu,��ƌ9
��r��$�iؽk7��{��ko��9֭]���M�7[l�x�)HLH�SSS��c<�Hޖ-(*j�`F�Ôb��͆�$%%��8�D�޽z�f��������o���\�լ1��҉�&��Ն�1�_��.]0i�$(ͨ׫�?��.\tȿ�
���7�xOU]���G�8���1!!}g�Rؽk76���v۶m���[`ti�ѣRSSbNRGҳW/���� ��%%%��}�Y_޶mX�b�nۆ��b������ܩMj&
���a�4�}�L������ְs�v<��c؟�Ⱦ�
�����9/b�0�7�0u�T���ǰm�j6c��Q�XlA�TTT�/�����m��W_c�޽~:j>b���ٶH�{�n�e8߹���k�j��v�n�Tŷ�z�N��3N�g���/�7��x��G�漷QTT��N-"�hh�U�w�*w0h�@�y֙P���_|�^xa\n�!�2~��Wx��W��U������9g�k3�{�1�32��E�W_}��۶��) �������/t�}���aԨ����$
� HMI��1c�&X�����7o�m�/���|�}{�`������x��yx��'q��7�GCE���!Ҵc�:v��b"�Й���z���O���SO>��^zn���u���q���`�>��- e�̙ga��ͮ�o�>}�h�w5l\���|�8� ���ϰl�2�}���aÆ�ܤ�Ƥi8�	HI1�Y�g�~�%K����X��t����7
���!��W`KcƎAff��L&4��XE�9�zˉ&�t�:�s�u�(�_����fw x9�������栢��u��E���K/��=�����/���)^@B\�O�{L�q�=�*<������e����Vᩧ�Fee��{�2aڴi���>�/pth�5
�F�B���a�x��Ǳw��6������W_ᓏ?6\2>!	'Nl�6�H��Ï��5d��i�pJ�S �Ʉ�.��N��C��� ?���|˭؜��n]m�n���G��O�`ѯ��X� 6.��_0hР���ĉ'W_��ض5�� �mk�>) ���C=�իV!xէ��ݻaƌ�T��UM��y�Gl�:�}��'x�٨t�~������u������� F�Q����C�{q$�ڬ0�-���'����9�L��@zj*n����ۯ?�= �P^V���'.��b�2�5�;�ߪ�^���<�}�?p�����K~�6�L8��p޹���, ���p饗��Y澜?7�p#6l�ܪ���k��r�mx��wO0�ɂ/�C�a��iӦ�㏇ѹ��z�ܳ����BQ+{�+z��q�X��Q�UABb2.��rtJK��{�#6[�!x<-Z���΁-��7�_¶�z�����u'2�d�8�+躎_�	�^s-.�݅x~΋X�n=���-�����+1��q��s��#�"����8�N��[n����P�8�t̘1��}]��>�5�_/X �����Ѷj������E���ÿ_��M����
Ǝ�+.�V���$ux�SZ���/��2�.+����ч�M7݌�k�A�0�58�u]���~ß��>��Ð���S&c�ē#�-�L\|b�1�
�}�̛7e�+~]���g���>_�8?3�M)�}��pV:q�m�#��>�zd��t⛯��?���ݻ㨣�°�Cѯ_dee������NTVVb��}X�b%�/[��K�b��mգ�5׏Q0v�8<���գG��� HIN7ހ�k�b�eA�MAD��W_a��u8��p�93�۷/����҉-y[�чa�k�a떼�u5��[�����н{�QZ�șp≸��k0��Y�r9���T��rᕗ_������/�ӦMC�n]g0\���
y[����c�ܹؼqS��<t����IhR������aÆ`�*�ٳ��z����0` ���PU�B~~�?����Zx�_C 1�|�fo6}>�9��!��_|�Ep{<���b��=]j���x�i�zlڸo�a���@bR�6t�\.8�NT�������P�a��`�1������#Z}����1�Y����my0z�g��]x��G��o`���}�hdee!55&MCaQ��ۇ�K�b���عc'�~o�}ё��	����4q�8�ԁ	 �ł���
�v��K/�T�hӠ.��5�W��nǜ9s0|�p�1�3����Ʉ��r�ܹ+W��o�-�֭���y�|�;�#G�0�Y��=z��g�T���G���>� Ji���ǟp".���%%u�<�����}3j�\���
t��	��+VT�*�_l]�QQQ���2��j*��i�-VL;�T�{�=<p`���S�L���p�-�`[�u���;�g�N|�駰X,�X-PJ�������DGVv�����.�I��e��N �$%���^��z�MA�^/�lڈ-�6��wޅ�j��b�����v�ü��93w�uN�1#�W&ҙq��l;v,�5>�a�� O[ri��(,,DrRR�w#z����yUs����eO� j��̳��+�����<�����	��^��=	w������sϴ[0 M�0s�Y�={6F��y>�h�u.��ge%*+*��x�*ԅ-��!C��SO��/�����ړ �����܇��+���{\s><n*+*QYQ��*Wu�i�|��={��G��W\���!��I�N��aC�5 
�����H'?�h��;����Ç���O>�����b�"p��|\�q�2�T���+���;�����[Ӕ©S���W_��.��	�a�W��*���HLJ�e�_��_g�y&,&Z��[�P�+�j:��}�]x��'0t�(MC�`��@5�K�|���<�T�y�E��y��ͭ;އ��.L�s󭷠KvW�$�WTT`ǎ�ޅhn:zs@��4�����)���{������5kQ\T���Z�խ���̒�����1c������ɓjs9XGH <�<3�'O�+���E�����%ψ��GRr
�=�X\tх�4i��ڶ�n<�t�i��� ����4���vj�_�01�N��K]�������X�����¬�z��rI��o�V@lL.��b�;��}|��6o����=?Z�y��5�����_r1.��|dt�Ԧ�]D�=��ů��~=	<�l{��ߪ���f̀���+W���>_+ۨ�ra˖�����ݙux]g@oV�i�='���:\x��X�r%���{���ö��P\T��e0�w0
���I�ջƍ;�L:�F�DjJ2���
s�p��c�ē��w���>ǢE�k�.8t�N�̈��C�^�0��q�2e
�9f<��{���S
�9�2tX�1�u���ܾ0�ZYj����l2��HW�_G��}`j�H_�@�G��1x�Ph����޽{u	�y�6|x�s]ב��[��v���:lx��뺎~���j��b��(���9��_�ѫWO�Z]�S�f@n.f��\x���������`��U(�/���Fs%Jbbc��)Ç����N�	'��ݻäT����d6UUU. "���T8z�V||���Ғ��/8b㐐�ت�6�L�y֙0` ޚ����%��塬��6�( J�`�48bc�������sЩ:�2��w�ݳ;+��_r)^x�y�m6��@M��"(,,Į]��c�l޼�7oF~~>�N'\�@�v��M�`�ِ��Դ4dgg#77����ӻR��`�>�#u,j����Ǝ;�n�:�^�[�n���P^V��
����@\\,233�77���b�����̄�:��~�ʊ
8�Π�[,$&%Ak�ޝ��p��o�j�"!!�p���G���vv����\�W�t���"�{f�III��p�Dee%*&1�-HJJl�픗���r}/��I+_�Q����Rlٲ�ׯ�ڵ�k׮�w��n���!6.q��HLLD�޽1`�@���=�wG|\��;߫�n����=�4�II�߱���xQVVt\�a����M!P�p�@>��m�Ν�p����N@)���!11	����YY����n{}D�_�7<�ԓh�&4&&f����ڳo���P���]��^z1v;z+��]A���x<�z��z���|��|Д����
{LlVk��F��g���������J�l6�b�"�no�6~����/w{m�p����hَ�6u ^�.�^�70��R�X,�Z��Z�������<8X�>(��ߏd-�fa�! ��o�4���p���~���9�4>#�&���b�u����3�Ѳ�m* V�VKBȠ}0��<8�ېF?��z���ЯlCoo��k?�N^�)ԑ�|?��kᡦ��|	��:Q4-�����p�""��$ 4�ërg	���(J�Hӧ2�E9	���e�8""�(&�.͏3�6t""�������Q4-�����:�E�:�5_B�u�����(-�)�D�˝���;���0¿�h�DDD�>�.��V��0�E%DCm�::QTif��z2�E-�$�6tv�#""�Zv/wщ���VJ��DDDQIDD����Љ����ha������(���;#:Q4����3�E)��{�����(j�7�+{�E��&g�s�DDD�K­rg	���(��`�5��E��̶�Q0"��Љ��� ����ֈ���Z�Я�U���;Q��yl��`�XNDD�D��|l���(���Y�NDD�D���NDDtؓ�Oe('""�ja��V�E�0��Y�NDD���ǡ_����[���8�+Q���H�����Ba�;��#�8Rё ���,�E�p��YB'""�b��rg	����c,�j-X�����Vؽ�Չ���V���Y�NDD�X�NDDt`Fu""��ő∈���2s""�(��ʝ����NqDDD�?ζFDDt�p,w""�#B�m��DDD�,��eX�NDD�Z0�E+�GDDt��ќ��(J���;�Љ���Xx%t�r""��֒��։���T�c�3�E%�!"":"�߆.�r'""�V�V�3�E��*�棵��E��c��Z�)�����Yx%t�C'""�R�oF��Z5�ADDD�R-��>s8K�u���()-�����C�D:J!���h]ס (��4�]���������*�]�+@s�	���jE������U�HD�Q�y����>x<(M�b��d6!PFm�밴�����ػ{ws�U���J ��W�1J�DDD�C!�[�* W�߆v�'""�B���Eo""�Ù���G:%DDD�j���tJ�����t@y5�ie�N	�� ���v��H�����ZGӴ����2-%%�q�Ų������#�aK)����φ��F@Ff�q���wy<�" ���j�U�{N�p0:�%@��iͶ�����pD�g?��������9ETM)��R�V��}gm\�a�:����F�~�w��ի��2"V f��b���1&�ɪ�4��4��4�R�T��`B৪��R5WE�T��k�U�f�.�PX�v����RhxW����x9.����R�<\(T�]�R��ԀR����u�V���o5�k���^�=�:Z���Y�~Ԧ���������j��d}J��u�������4��Z��p�	��ʂޠ��^��u��c�o�5��b�x��/=��WD�H�����9��:{�~���������nHBi�{ͪ��R�4����k?���F��w���'��f�!��`geI��5�|M^�~�������4�	��t�cP��V�p��Vw\��n�f�'�z}���`����~i�'|�P������e��e��FK׻�68�W� ۯ9$���dݵ��p����u?t����������K�Y_��]�j�GR/���\�dX �5ikt\��*e�R�p��I�ɋz���ͯ?��ڹ};�~x�W��]��E��O�����FGT},�4��o
 �t]����߯ ݯ+]~�_��D �_W��t%"�~��s��oP՗]��^W�i� ՜ "�7H"XMŊ��>���]���>k��כ����}{��m�9��g���_y�7���4������]�78�J)���x���q�I'��^O���_��5oIݽj��O ��V��b��Ҡ���"5�RR�����R��$5W��;_���U_���BW_]�҅�r��ȁ?���M��r��7�R����d����/U�=}��Li��i
J��MдڿiJA�(/nKE�c}+M� Д��Ai�mk�Mi  ���;�ݨ�j�,��Q{JNIE~�<�쫇q1� ��)[�fʼ^�}>8u14��4��~�AY4(� ~?4ѠC�I5z�_�h�P ���\����k�R
���5��=�j���5�^[k�ª��5�)S��/uWߠ�cG��ɧLz������-���+��s�|6��0٘PRZ��n�/��r�������#F�87--}魷��ߏ�1���d�l����&��-W�ƥd�hT�Qu�T����7��n+�ꭣ�i�h=5�u ́�Oլ\I��������R��ڂQuU��K����[����_�D�N�	�ʹ�p`E���Hmy]�4����P��nOS
�i]��L�u@��lF �X`����*������t�	�v#..J)j|����Kv6X/�y	&�����D|B��v�G�7p9�� Æ��m;v���."�Ꟈ�����?"1�Xi����*���?�㳟�[��E�05�ک���L8�$�������M�Pغu֮] Hk�a꣏?�?���`��������'���Y看��6�sύtr����w��w��[o뒙���a���Lr�=�8"J�""�,\$	tMh��q�ۏ=q¸�YY�>,DD�XB��23�0c�i11��A?.\��Ҳút� l۱w�u֬^��_	������~�o����[o�S�<�$ŀNA���`��1n�ñ�d2]f͚�ض}[���j
@IY|�!|��Wh�p�RSS�>��c^�~��k�N\w�5�N6Q����[t꜉�cƞc�����ݭ�ye��ڎq������#�=.��xi��O�ظ���=�8�#.҇���Y,�SP����٫���7[,֢`�x�.��˯p{�	�>��3<��cpV��q��d6{323������7�Ήtr��Bb@���:�����:u�e�Z����l�2���V��
��U�qｳ�o�n4�(�����G5�I���6nğ��C��MDD�:�>����k猬7��t����N���?6��""���Η���ILL���#G���8"}���ڮ� ��={�]��A���d�'��}��*�G�w��l1A��M&�;;��"���.�sϽ�>DDaa�;��q���d6W[���b��%�r��j�O?��>�,�n����aC_7�Xٳg���H'��(,�d���>Đ��Щs�-��Ш}���8����T�n~߬�p`�^;��11�srr������G�?yB��MDD�>f�s..�������_�UQJRR���oDm���ȁ����f��٭[ϫ����/��F�����EXB��F�����,��>0�}c
%%%X�|y��j�������G|�}�)$%'�w������S&cǎ���D:�DDD�G����?`Ѝ&�E^�����rE])]D��>�N�A�i4��KX5���t���&"":8���[d�tØqGO���F}��a�u���	���`�|�J>r�a0�X�e}r�] ��}���NpDDt�:u��8�̳�&$&m1z=)9U��u������!�͕f����go����s��_o�!�YMD�jlC�f%�$#77woLL���K(���bٲe�Njuj �׋�_��?�F���0��~�j���x��"�t""���G���={?��I����9�|�p:#^Jy��s�vs��Q0hȰ �~c,X�l&"":�j:�6��f��g�"[�n�h@�����#Gs��������w?��r���]wϊt|_|���O�p��Wh�<zbb������v��ϛ����u�ge�?�x�4qR������й�Kq�Eg''��
�5Q�$�=�`Ăys���8�v�=�x(3���"�Ý9�	��CRb"����6
���˖.���D�ÁC*?��x���vW!�8�f�ٓ�����E��p�ݳP�*�R���DD�c/w
Kf�,\q٥����U�f|ڬ]���8�iS V�]������A�`��BrJ��G;��S�L����x��q.E�� �KF�;�j����GOLJ���y���ED
���/(�v󸸄���3<�s& ��>�t�z_|�N�p��:}P|B��P��<��#�$���x�^y��G�k�nn������� j6Q#�#��),�'O�裎����8�-'�K�.���:$����xꩧQ�D��vMӐ����i�Ϙw���`���8��#��DDD�ܜ� "Z�^}�`f�a������^3N���e���>o�IbRʢ�&��k��!����,$":hXB����J���V��f=�R
�v�Ė͛Z:4 %eex��G��/���4���]�u���W_nY�|n��o��B""���>j,N�xʉ�ظ�6kM3�#�=~�J�^�_�|z�8b���M&��[���������\�;�~O������s����GϞ���o����묬L��^ݎB��ޮϣ+ �}�=�x�	8+��txD��Qc�z殿�����>�L�����(z<�������]�u��xxUȰ�#dێ�ZJ�ۺUN8�$�vsh��m��㏱�c  o��v�����(��߸ 0pА�4�,Fϣ����7�k��."RVQ!�\�g1ޮ&��շ_������{���#�eDD�;�Q��ر		IHNN^n�Z���R(--��+�m�~��ƛ�׿^����oUӐ�)��S&M�{�Y3e�M����t�E��3N�̳�����ۨS ��K�UU��R���?�$��䆬jOLJYq�)����,"":�XB���������p�n�ܚ�kPPXئm) ;w��}�fa�0|D�n/�޽�_9͇}�����HgQt{� "澹�_2`FIZz'��ZUB�W��t����ILf�a�\3Y�n�{>�ҫsmW��Z<=��HgQ��UU �3�:�ŦZ��*��}��U�~y��Krr�W�k�����3g��3���0y�4�qNDD����
#G�i�Θ�P���+/UO�K�""�M�����=c�>�d �DDD-u�5��ڿ\ףS�����Qc�ɞ���.�׌Ӿg�>�q�!K��͓�o�-"��v�x���"�-DD�Nq�*��;��O��!�U۾}�n��z�*��>�>����S
��>�0�9g�9S߱s'�v�u��""���[�[3���&�%T)Z��R����󎤥wY:OLJ�8q�Q�9�  �/�t�~D=z���i��pĹC{՟�������V����G�l7����G��= |2�K����HgQ�qrj�-[�`��G#..n���(v:+;U��^���%蜞f8Q��_X��+�-�Qk��i�ҥ�[����7F��5�V�9-*Q�=��l�~{���[��qY]rdђ%!����̺���cBV�wꜱ����;�����@���������7ބ��G�>�ߡ&j��b���n�ED>������jW���P|܉���7��>�t����{ ��S��d�;ĸ]�u��M�>_�`�f�:9j̸����M<t�c?.��z�?f��g8�9Q��vƙ��UW����^���ēN�����t�������J偗R&�ֽ���xc��睏��^�]'"":r�����Y���G��ޣ׶P=�kwY�|E�������ǟ�G\�vs%)�i�Κy�$ p�uk�ϵQ��v~[�,��1�~0�r��~�?�Ou����_~%9]���jWb���{�	w��魷����|�]&"":򔔕AD���N�b��hG�t��]���{ٴe�{�	!{�k&�<􋧞y���7܈y$һKDDtd��変�\i��xC��%3N?CV�['��j1�X6;���k�������W����G��Y����}��l��\@��8d����h��<!1�s����$"�_~����#��DDDG�5k� �Sgddgǚ��OB�������Ymr�	'~4��S�}�y�:�_��M""�#ߥ� ���z�����u�׀���=����:�\ �眈��8q�46�;>#>!��s%�]���DD��nl޶-һGDD�q|�� ���g���[��f�L�>��=���~��7X�zu�w����c���7��~������̬�ו2�8��cbw�vƙ�fv���v""�����G{܈ظ��-
�J�9b���õ֦�:>�/һBDD�1=?w.�="��=z]g2[��	��"i靾0hp����b��a��""��������N8��8-)!1�悹R&;n�޻��Ǥc�;"ªv""�H[�`  ����{7[�뫫ԃt�-��w]|��h�N'�{��H���o��S�L �쎋�L%]w8�^�<uZ����GT:��N:���@$%�"%5�j����i�FU��j?5�Sv�,t��k6l�t�����1�dA�Ι8pprFf������Ė����LIM�ӳOߞv� p��wG:�DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDG���Nþ�C   xeXIfMM *                  J       R(       �i       Z       �      �    �      o�           ����   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��    IEND�B`�PK
     �8�Z�����  �  /   images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.png�PNG

   IHDR   d   d   p�T   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     �8�Z�Lz��L �L /   images/256658b1-ffe9-46c3-9f0b-70052a8fe00d.png�PNG

   IHDR  �  �   �X�   	pHYs  �  ��+  ��IDATx��|V������E� ����)aADp�m��[q��:�UQk[�u��l�(Sd�����7����wr�Ҿo�Jk�����<��9�9�ߵ��V1� � F4$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A�(�~������c��AMuՁ5�u�������p�.�Gɘ�i�
����1�ϫԨF���6*,�!��3i�TKbX�%66����I��gqBbO�Y����KK���yUʱ���VVV����o�Z�].W�R�Ԩ�j�]��z�q��o��
���w���|�>ӧ�c�b�S��s'�O-=^V_=%5���dqAbO�Y	x��j�jKx��g��::SO��O�X�ƹݞP��v����
���3��� �\ܙ�}b/���o:�Ri�)��.�jL~^��ܜ�W��
k3fLQBBB��/�_�3j*/�`V�رcI��a�=Ag����O������<�ő����&��i�A�\�%���T*s:���t0�n�_�:���~&�|I��{��UJ�w��O��'��>ߛi4����5����q��9��F��dj߽s����ɦ����322�ASH�	��444���?e�Y~�������Y�b6�j�d��g~��!Y�V)��3����V�x��q+�)�������ʹj~'����S*�\�5L��3~ߟ�:�ꍈH.�G�U^����a���Hy�ݿ\�eK̮�>ڸ*""�&6vzSF��b1� �'bX��+o%�~�=ל�89G�5��ydxX����
���tZ5c���|\��Vs�\�a��нZ�f*�{���p�|\�}ܣ��B�����~�F�t������+z��|U``��a�s�`���,<:��t:f�;YO_?;�ޥ����z���ʓ��^���7TTTl;vl#�a�=A�
����j���F��>|���*�d�ޠ5����
��ûf�w���v&)���px=n�G�V�Mƶ� S�A����u��ڮT*�*���+S��*�����v+�����(��q�ݧ�z��S�Z-[RGk����q�4�B����RxX���::�Y__��j�&�tv%lްyv~N���[w�;s���H�*~⇆Ğ �az�{o�7f�g.lom�B����tڠ@�Ya6<y��Qd���˺;Zw�J�tH~_o�(s��`(�<qr�ĉ�'L�Rb4Z�CBܡ��.����yH���������Һ�{Lojj�T]Y1�QU�a���f\�xi�̩��c���T*+���;:���{�����ܴ)z�5�������=A�����̏?Z���d��E>��r+#�BY��,��m����b���hsi���QW�=)q��Y�g6dL��:+,�ʒ�]�գ<�9����{����e�ڸ]���b��'+$6=�X�ľ��q�2��Ա,)>�e9����͊���ݶg�NӾ}�o̟Ny���=A?(����7�xg�����٭�MxҤIL�R���f�ZYuu%�.�[�P��v{��ys?���+����T7{�}����ڵ��s�����|16n���z����6,ٻo��ͧ��5*, c�d�5�^�j���75�Ym��������;�|C����8����=A?�������'�O����7Q�����pQ��9������YG{����u�����Ą싖.�~��%��9��CGW�v.�k^{��%[�ܺ����Ç�����Ξ��,;�kl�W��5��v?`\�nk��,� �����_���B�jժsy��7775_8*(؜�<V���,*�!�]����sK�E�V���[�r����͌uGL�h!qL�炟w��o)߿��M_~���?_ñc��&O͔n��uҞ={ّ�9���3U��>QW��=�W��'�����_��������B���*���Xrr��d���ɸ��:�.{���3>����0c��SW6�4:�|+��\�ȯ�jhl�%�+cΜyA��%�>���U���$*��w����_���X��G�W �'�ƚ5k��{�}�dgg����	ܣW���2���lLac���n��Y�|酯L�2�Ȭ��+"##��, ..�^S�gMi��-_m���]��<k�ܠ�.\�fa奬��-�d2���;vgMMͺ��D#��0$��#dpe8������i�)kkk�*�Jr8���dx���U�0NYYY��v�o�v��Z�6��2�Neaaa����UWW{��z;<o������g����?�:�%&.�x�m߸��ŗ^�eg��3B��@���)�lo��Z[R�v�&d��}�3��CbO#�I����an�#�鵛^y�-cWg���t��>I`2�bc��~��#%%�388HYVV�����^o@]mmLO_�J�R��jGL\tSld\�}��
E�ܹs�������[�j�9�o�|���R�ә&N��ƏKg>���46���}'�͙������{�M�l���%�_޶뺕�Von8YV|��i��5{�t�X.++)P�NH�8�߃G��85}��J�{}� �C���⚕U�?�Sg���[o�ڛ=���2�n������n��`2i�
��U�����9Ǐ��u�\m6�e~�/,,4\k0�L�ؘXM�QL�R�~��wwvU�U7��v:t�=���?U��NZ��3����L�G�fS�G�N4�'�YscS��l�t�+޿���=������n�.<���mDUuŭ3��2���b�֭cN�M}��=��1��w?��?�=A�����UA'N�*�OElڰv��~q�
�j��	�+J*�w���fSPP�&**�EEEI(�s8̨3K6����*6*8į��bw�ޙn�e�,66V2����L��0�����G��pF�w8�W��~�a��1cJ�@�گ;xpm�[o���V���iu2Ʊ	&���.T�{{��*����,[��}�4��$M���嗟>��㍊��㿈��0:���ٸ�Ө7��v������r8 #{�8K�{��k�E>�x��ڪ�s��	.�=���.%���]{�0��1���X�7�V�*��YYI	���c������.��Rv��!�xn.��4Ҽy粔�6~�xQ_͏���e�--��+�qBB?���0U@@P��q�+���s�n�fSNN~�'�!��>��`�ω��ԢINzZ�02�?�kjj*_~���y���o��F6R���v��~��<��T*�OOWUTְ��zI��E�:|��"�k#�� $�q����~��?$�[���ްX���Z�[T�\�L�����{�2��ʢ##Yr�6.5����`{s����o�����d�'N`[�����v͒�$���˂��Xqa+//g%�eb���.*��N�r��o���QoB�z�ԩS�UX�&�ޱ��hNN(w�c�v��s��cǲ��:���ҟ��U�_�e$���jӨ�Ĥ�UՕ�q��)&�^ji�e�N�R���;v,惘��Waq�!�'������/�������*�F��fWO���;�ط��r�a�ys��1cX���{�]�o�C~��z�q�م_�R�$���Ē����l�l޼y,/�۶}++**b�M�X[g�Z���(�w��»��|b�w�R�Z��Aդ��fL�v�sY�)���ň�Amm�����a�ٳ{�_�=��7���ǯ٧O=��d��W�+jOq�oc)i�����GGG��fq�!�'��.�?>��	k�o����8O��K~�u�ٜY3��Ø�]ΔK���������m�^����-m->�^'�vE|\���v���|���6s�46g�L�P_�8�*++E4����=�����
o�ǅ^�T3�Z�=�����o�XXhX+1��&9�F�b"G����?�|=a����,\X�~�`�=n�lz��WH�S����RIY%Cӝ���(��=��~?H`b�BbOg��v�yYG�V*�����j�o{�ܹȷ���J�ƍKe�kdk>Y���~�������=s�f.��QQQ���Ϙ��"
�,Y*���Y~~>۴y���b�j�z���J�ZB؞��l|���Zč�ѣø��Xk{+���#Υ���9�v�)v����*lu��=���̞=���\�ƯsO|b��꺴��pstd(k;��j�k:������,.�G$Z!�8����0k��s�=v�	��e*�JU\lkmme-[��l�����Zzٴ���ŗ]�v���>�0{���)��{���o�.--�ӫ��-))�����F�Դt65s�X]�P�a�?c����M�4a���7R�IĨT:��鄇h6���ec{v�.��r�w9]����j�X1.j,4|����2wڬY�3gN��߽{���>���N53�lT��7r�M�=!'��'�&�;�w��z��Ğ �1\�������;���j����� �ȣ�\HH���رcǘ�a^t"����3��cOJ���7_�s)Nq��ں�膆&��ϙ�.<����6m�Ċ�����
uO�<e�k��V�އ�e����4����"8$P�!��u�؋/�����7�1���
57zYaa>	f���Δ���+V�vⷿ}�貗���W�u��;Ƅ�Eu��������l�ږ<����$#�3�=Ac��zo�u��Å{6z*���#|?c��m��_\\�5k�&��_����$����w�yd�̙b��-[�dnX�neUeU�b�h�"x��o�9zL�CU~l�hӡC��|��5K�/)����������{{{�>��z٤I����/��zN���v�v;�N�c*�f:u�����ʷ�w�2�ӳL�TJ���y�[ZSS�bn�UP(�8S��|1Lپ}���z�j�Z}��fӠ��f�1.�lΜ9B�Q����❕u��5ulʆW^�)Y豤��?x���SS
�Mr�ϟ����?~���c,�av�=!-�-���h���������=\�c��
��m;�馛؉'��ÇŪu:��V�G�7D�\�3v���O�����Ԧ��r���f�nZ���ȑ����s�.:��4<�@bOÔ��zgjC]��\�#���$x��c�;D���yX&ğ{�黹pT�|����/+*���޶���W��O���cݺu~.�L�VKN�������c*m�F~�mŊm�7o����g��o�=&Y̗/_�.��B1�h��-*�}>&���,+W���M������c�q��{�+�o7�Lq�]�a��"rKg?��2Fg {��p��{ﯮ�@)<n��፟<yR�V�T��s�eG��<v[LtL�O�����o���w�!����兾���ɽ���G���Ν+��#G�����FnT���|��ϥ���T����i�9]r�%-۶��ێ�_O���t:%��&
�0��������` �x�����$����iC�w,=��#G���ޫf�����uw	�][U3�߿J�Z�g {�f����9���p��Wh�������eӦMc�ׯ�����"w�j�*?�����x��<��3b,.��7_��¢��'.�=Z�~�駶-_���7^���-['lٺe:7.��{�w_TT4*<r�KT��*�m۶լ�dU�A��ō��X�|Ǯ���³G�Y��c���>V[]gLJJ�΍�����m�L^���֭;8��l6���k#�_CcsC㤎������A|OH�	b��}�������\(c�NC�]��Qq_VV&������gG�������舆��jkk-**8���\?R\tYww��� ���%�޺��s������c��W��S���p�xK�,����Ƿl�ꊏ�WA�!����cS�LFHVV�8G|�������ɳ�����09�`�=;v�?p��ew�*�J�/�^��j�LV���Ğ8���0S��9m˹h��Å�C  �b����0�m�Ν�cǎ5��������O�>^iai��fOs��*��ŋ����?p�.#=����z}'�g���x\>�l�: 4�ie[{�߅�w|�#���t�J��#'��PB�1�Q�`�O=) �?���3��[�ܷ��^y}Cʘ�����:n���Xz��3�M�X1.=�@QA�T�ק������}S\\�:�F�{�^�����q;�?Ey^�=<hL���c��������{��{�<������{Ϭ�ݥ*�2c�3�!%����ݱ}{�/�{�B�}]6�(�����x��w9�>�F�w�⊺�1�UU3������c: ��w�ƍ�n'��A��q�
LP*3��-iM��M�]���Ą����3��kn�_3OhHh�Z�v[lv���`N���d��1�8���0�ĉ����).�K��=����Eg �(�Êu�G�fǏ��;;�~�O_-���{pISc�e���:�-r�))�"Wo�Z�'MJ��Wu���fx�>
�d���
��\�zs�sO=~���o�N���{z�C��=���۷��	C$� �;>>�%�+��A��%�{�fn�$�v�/,/-.8|���_}��7˖]Pο��~\�L�~��߄���`������E3�8���0���(���X�թ�]Cxe��#���zܛg�������i�gW�>Κ5k"gg�����pq���z��c}YYY�7�r�'vc���r}S]�.�J0$�so�+elr��C{��p�܅?/=Yv�Z����߃���xD]*�Q�9�x�6s�`[]����G{a��&��Ǆ�sZ`��qú����e?"P�����ڜN������G�o@��ɳ'�$�1����O�|8D�ox���C8�Z�\o޷���A�!9����+��>�?���"ae:c��0�9s���7�pC�O>)�-..kio��jDc�$&&���'��\�}������r~j��`<��f�<yDpNH`v@zz�0Np�G���xm���|+�lK��ܸᢟ<%s���[�z��/df��ƒ��ǂ�9|>�W��p��%�/ay�L��@bOÄ���<0�{�>�_(�!r�1�!|�+B�\�}-�-�-_�k��C��0u�C[�0���-����3�pv�}w��%ڵ��744�Y,��N+��@A����1u����>o�.G�^�W�\)0��B��&��'O����҄QR[[+�򵶶���:�ýz���>�1���Qp�W��J***F����
>�⦦�]m���S��~$;������Y��@ms���=A���}}}�c�W�G�����v��9//�ŵa�ҥK����޻wop����J)��!���*OUu�%*1�G�B�r��@�Fm��"���/))�Z�VUT�I���o^P\T�4( Ȁ�;l8/DFǋ9�)i�����:���OOO�/B�1QX������5����|���4eҘ�)5�7���3fL/���i��5p����)
%��n1{�{AbOÄ���p.�q��!x��Dq�}9��Ű;#}¾�/����q���EFYi��|-��gφ����=��D@o��!Uaa�h�=d谗�����i��+���oY���cbb$D	P7 oy}L��5g����"�)w�9�(�F�9��ʏ�t�%^��˖���)Z�z�%���Wqv\ww�v�qP3�靌���͛�/㢷��05O��!����1!a`�#�N�Q0�8���0 pO=�T�#.�hӯ ����l��%d����z}��Y���oݺU��K�]`��֦e��!���.+;Y}�]w펛���7~�1����z} ��x:V�[�hQ��/��?���R*�����bw���"�PYyR��s�9�&���E���������o�j��܅6�n��O�x�;׭���ͱ�1F��I�ȩ���e˖��_�F8j�ѥP+<>���}�לi�*�U���K� �'$�1<���0.�F9�P�/��#�����xJ��˖���wO�o߾����y���a�!4_UU՜��s٥ˎ=���b_�:�r�,���ӹ1 �υ����q��w�������)��֑N�~hы�{���[�����`0 B���5��$S�ө�vI�-�#e���ʕ+�{��k��w�Z������H��ϟ?�Hv����^s�Q� �9y����^r�'�7$�1())Qp�8�?��b����s<G���Z�[<\C�333ݧ�����t�F��!�΅�SZZV�dђ]C!�7N�R[[�������,�h��]�;���s@��I�&	1/,,a{�i�0H��������{@�P��40���Ï������SO�����[��8ݞd�f�@������z2��۱ԫ��`�V�����p� j-�y=>{�@bOÀ�� %�̯������Ã��56mas�]~��f>}T��r�-�N���� c�{]]]uMuŇ}������=1��rM��i�]9z�C�l�5k�J�qC�-X�@̫G��oi���
Q=>o�<Q�___/<z�h��l�:����	��أ��;�s`��S(�c��.��r�G��	�����>K":�R��5SkT�Q��@�8���0�j���p���)�W��	�G�^��"4υ��_�]�������wL�O��1��˽oGk���}���-7�6�������h16�u�PU�1�BF�P=��fΜ)�
�����v�m67Wj=��%�?}�tq�0 ��E�!?g.Z�eF���|JJJwl\���S���s2"z���#)�RtN�D<����h��W��p��&�t9�?�� {�pAWq�3Ωf^��!t�",��Gę�;!)���i@Q����O�//-��X�{��t�ݻw;F'�>RTV$﫼����_��ף�c�y��x��n?B�s������j��;\��;233������0�L4�A� !~,�3�	�/V�������F���/�.t�q�Y~�Q�N�3"�!�ɵ�GU���e���T�.����)��?�l�$<{��ސ��0��=�:5�Ȟ�>D��x������3>>�����b���ZMIQ�L�R��v����p��jjl����o�ݺm��w�c���s� Ӹ�*�*��F8�>y����t	��t�>�Ç��vuvy�w����}~N!�@!`tD$�(+g5�UL�|=�R���=N���_]�3f4��o���s�垽0z�o6���ų���Wb��-�|�_A�{�@bO� .�7<Z����G�!�t��[#C�:�}�m�?��T�\.����T���c��1Q{�?~���;y�r��MF} ���0M� |R�O��Ԣ{�ѣG-III�<�̳��SP�� /���X �urQ_B\�h�s��qGLtTim�ߵ��;�q�4�N�ǫ�hD�Ke��E���W-\8r+��5Wp+Oc���E�O�`�?
�=A�e���P�`)���C�\��Փ��:�)�9���x' B �@��\��]x���S��¸�����1�Iŀ���=����x#����ͣ�.??�u�ĉ�_�x�/��xç��uuuE�5JVh��΂C��޾n�ѪXrrS*%OCC]۝w��<t��g���{$I٩R��
I��z=����2��V�X���ܸQ�e�}\.���+�`q �'�aDW�v���"3�N���iY\��z���u�|l[Gg�@�xʠxs1v�]��33�n�Ey�����}��3���@>��<�q��q����G������h��O?���B���@][GۨQ!��_UU����8D
0U��6����暺�+W����t�U�w3�B���d�+�O�gl���G~�H��n�.1��}oo__r��ZFg {����XE^U����" D�vgg��`4vpA�3�ө�1O[^�{{{��j����ڱ���6O\�f��|�p��E��C\�����ɽ�QUc�(� S�zo���Oy��C���с����Q�r8��;���zV��]p�,=-�:tȲt��iii���=�t��?*  @���XJ��SkU����#�P-77W�_P���5M�P�S�B�:��@bO� �	{�X:��	qǆ�����6fS�zEl?++K���/��l6����(**懺M.�����3.���( &�PT�9� �"W�����c�]yy����;.}��	n}C����z���� g4�Ae�^�U��Jtw���u�U��^ii���1���q�8N�N_�w��`�EYYYf_�T&eA��Į�����u0�0{ap��������H�	b�E������'�է{�{x�r���/!!��{�B<O�81�TK�,>���S������Kԋ">n��ǅ���~	�����v��Gm��	yz��Q̱wG�G՛�7�}��]����{zzB�㙵�"�#ִ�r�ǏwY,}�,���kPZP�t��ʁ|~?��\������曓>�����T��at8\������7��z��Mz��Ğ �^.�X��'�Ň�A�e����y�X���t�mwfp����g�V��WUV�_t����~œ�?y>7&b��-.�^��#GDQr��L�:�r"��қr��_v�e�����@�����$�?�(�C�������M{�ۼz�	Xt���ܓ5�w ��q�5�NNN�l��5k֌�ꫭ���o�)X��_	��6̌���O�4)�a��1�8���0�{�{T̋p��fV.�?��1�>00o����M�u����F�ё��T9�۝NG�-��R��˯]���o����N�u��C��=m�q

r��H��ʟ^YϷ�s}��ק<��C�
I�Ӫ��iw��Vװ�s��+���mٲ����s�����|�g���߿~����9�f��}8G��['L���F ����7]��а�_k#���jc����v��~;j'�����"����^~o�rc���{@bOÀ��t?�C�$5ڣ������B=X=/�Z���GtvvMP�����7�8p@�������1��^}KP`И���G��`�:�u��="a}�;vL4��b�z�u�o�{`��y"�p����h��� ����|?7V�E�EM,�0o޼o����Ծ���сB�pN��Z,�������_�p.�3���#��Q�C�Q�)�� �;��)>a����fAqA���o�� �#$�1<�r��6�v�Zh�;���������G���D��߻w�8�Z����^/����h4s�lW_���~�beyy�L�J�			��@�X�f͚u����itj��	6�|a$�;G֬Y�իW;R2RjO?�>�`̎ۖi�Z�"ŀi�2X������ؔ4����6o��������/���/8��=��c�^m2�Y���J.����4q�s��I/�����Ɔ4�+p]N;7j���#���
g�a"������w�����<��R���8D}��
�=A�G���_oV�U}�[���{���:��A�9����z
�p��%!�?�7�b�?o�;w���p��B��u��O���K�«/))��Ǎ��ϡ���l�o�p9���<0���At ^iVVV��ٳw�7��}]]]���Ӄ��|L	
nL���τ	
��{֋}^^^Tuu͵��"���w������������ q���b@�^��Z�jkk����kA�0���0atLL�J��ȋeN���v@^�V���\ҕ�N�F�f�:�<>>^BX��O?U!" /��g�f۶mS� !}tAA�h�s������տ}���̙c����C�z(��r�z����xH�۷O,��*�M�6Y����-�sA�������?�0/�X�Ұ�PMgg���\���=�E�^z�o+����^^X[[�i6����?�R�������%�Y��:�,��BE�9#���=AbB��$��U΅�X�.7��#���FOXd������5-��r�\���'�~k׮=�!���c\��ܕ/2:B��Q���;�`����Դ���.����ac��9;;{�Ag0@���z,��<�M7���ν��믿���q��z�{��	���k�p:X�F���u__�%2"j�UW]U��_���͔���***Z�����h�������3�����QB�-���\>��g���.�FL���=A"�.�J�ƅT�s;8�|h<�*������F�1����y���!������q!�G�9y�O����X� �����k��{>K�?��6~�n��cG��q��'@�?*��`�ϻ��}�`�[���7^~��W�x�}�V�^��ٙ��]��7~^>��^{�]������Y�!�6lJk;�:���(���A�����9�������ǆH�������NEGG���6 �Ğ �	Q�����{��V�o�ix\�z���@����;��`_�5�a|.�C�va@8���<yr����G#l˖-cd-�-�믿:��s��	����?���!�s�
��:t�SVVv�wO>����.///��n8�?5"R уa����p�y��v[�����f*+�����sZ[O�r1��V�r�j1���=]��R�`}�}b?���6]YDDp%�+2������0A��t?�䓅�v.�f��!AY �EEG7pﷵ��8�fwDc*���z{���
�����Qe�p>B�xD�������~�M����#=]\����uu��h5Z-�G�v��>/7
�B��\R����~k~~��W߸����r.�*�"�|}�7�$��~$��mn>2����B�FgF�{�N�s��G��p��%&&��0��Z
��a �G��;M��.F�{�FD��Wp����,/V����6�R�ʊD��C �^t����T�C���=��!��Ə/t��r�<�$W�ᬖ՟�~q���X�fHlsrr���/�)ƅq�q��������������v��c�����Þ��ӗo�rӃ&s�	�z+]]]}
������z033����ٳGUY^<�0i\̕0�p�`(���=�OL��{ ����Lkk;"m�>�?ۋ�{�F�DE�p���B�� @�e��أYG'+U�4.�:�=r���Q�./�q��$��00^Ûĸ������������9g�7�2�322��K�^s�5J�Rc!{� A���F^ّs�����x�.�����_Q~m�q����Sk����8W�V|��>���ȍ�>v��T��N���:�i��`4Gj�zq��kjŔ:�?�z	�O��F�10�ĊJ~i|�~o[A|OH�	bߧ�jQ�?�q9�"�>������8�zwO�V�T�PԆ<�r�B!/�����IMM�dII	B��ŋW756u����=��cor�
s�\{�O�9�w�
�R�p3Z�����}����.,(8z���t��k���&߽��?���/4�L�� 	.���Ғ���)���+y|cgeee�윜��{��_x�6�-�[[F��l䏡�����nJ��qo��q���,�����ǟkE����Z��q�PkU��8�e�=!�'�aD�:֮P)��w��v�!���!��r��Z�����8��Nrr2�I�����vq,���b=��}�����ƥ�����tY��W�~>{��ٺe�e\��X	=��!������1�~���������?���Ʀ��8OD$`��,����f�8s��}��p����e̋/�|eQq�r��6&$8ج����:+��4X,Ex����""E������!&
�$�X"��LLL��TQaq& �'�a�;��c>�E��� �d����y�X��$���A �G�a|x����r�^#|��o�������[���ުU��SSS�&�%�]n��g���f�d
P��M�&�n��P��4Ԯ޻o�f>�\�u�������55�W��5��1"�w9:��w���G���'����&++K���_/۹s�]��3zzz�����G@��O7��op��S"�"�O����߮����x�C��,~�X�W�V72�8���0"66��c�6���-q+������д-�A�~�r';���}�	B�8b��(��^�/==]��_R~��w�=���M�*��ޓ����g)$�����!е�����YTP��G��رc���s/���K�޸i��5ZM4��\,�����x�ҥ�>��'�س�����G�k�{nh%���)q����y�9��Eő֡h���d���,V!���x��`\7�Ԣ�!�����AA!>��u)�NFg {�^���P���!x�"ޓ�!|x�p�'�`��{��F���v�m���`͑#���^r����?���w�����y�%�{�5��p;ЁH�ر��r97���/ݼ�溕+W������,_�f����8_�!�\��⯭�m����˭��x�l�j���XXXxm[[[bgg���0^pO �E�xËG'<��!{�yuu�@�@��A�"�czc�R��&݈Xޗ��!�'���l2�wj�|r��� �P �o2�~�o����@4 �V��?�'��������4wGGgyyY�SO=�.##C|YNNI��o��?&�����5�1]��/7'�yނ���r�-�|��?�bk�����-[�n��F��Q؇���
�{�z?���o�Y�d���ttt���9����#�@n������;�v.�3p�����(����>��%0���1X�������O���A|OH�	bx�lT5��n��yyy]{�����x*��Eoz��0��x��# ��1�i���{�����
&N�X�\t]U݌�V�|=�?��g��IM�4z�����'pT𺫯�z�_?��?��ѿ�񕟬[��	~|rll���?�"������M��|��7~��?��ݻw�jnn���X�Ψ75; y꣜FA�$�L��	���b<�l|U\���O��9�hYYes@�!�loL��������=�.N9t/��!�w�P/�OJJ`��ڵ�������9�J���ap������q�E|��u�u����zl���`��K=\�]ee�o���}>_��Tp2�������Grs�{���/����G���_����?�' 0 	��"��Da����98N������s�}������l�ԩ��Y6�C���;�c���[�<ܫGټ�������=L���@)����bj~�"����W*a(���f�F\7U��u�����d0���/��.F�{�fp�ݪ���\ܱ��p��CD���z�#7�f,�h�2T$�R^w�mq���M���FC��]�
,V�=&"*���Է��ֽN�s�������8�`�C�u���n��H������u~e`���?����1  0�{��
p�4���a����7�|���
ϖie(��ꫯfq#kߔ��i���\y�B<J�n7��6;0�tZ��ao5:���'�P�%�X��V��w��gKKOz�x_J#��0�߇Ğ ��u�����r�b��`�\=r���C8 ��c�6�m���ȅ{�aa�5���I磌�b��-�w�V^p�y����̙S'�+1)%1!Q��s?38(��KMc���e����:t����Γs��He����?���훥��M�s���=�p�>�����{͕W?�«/Hg�����\Syy����͡|��{��"�*Γ�;��
�Y��>�.�#�"�=9e0
�V��6��I��JU(�G$�����;}�a���@bOÌ���ns@@��a�s�^���!
ȿ#��GU�躆��w��e�#�� ,�q�޺������:v��|��_��~Lxx�()�Ȅ���1�^=ml��X�pN�?�/���ܲ3���o^���}1edd��cq~mmm���l{{{��;n���/��ⱳM�:::¸A�ɽz��H��Z�,����2 �����z�퐯��&�=����K6p����,ǔ��;&^��!���3��7 �'�a��,���j��J��A<ރ�8O�T���b.J."Z���N;��$!�V��M�8�A�/����8n�����--i����8�d�If6�E�?���?~�Dgsc���ѫ����H�ǚ�ڥ�A�11�QJx��q����!RTT�mw8�?��o~�r�c%/��;��1��{���}<��«�Go�����E���|��
��Z������d6�˨�3b/G p��\�߇�������1�qC*�Q�>�oBbO��۹�p���������@�[��"=�!6��!B� ��*��9b�>C<_XXhh=u*�{����k5ڡ
r.������%���>]��>v�Xد{⮆������.@j��r��������/y��W���2.��l�_SGG����UqMY�z�G/�C�{�@=��[ʹz<�:c,x�96����3���tC�X,�����H�F��7 �'�aFpp�#$$����O�!,����1���q!Z��""���������9���Od�w�F�<��ʠ��+>��*��d1�3g�X�~�ڵ�ή�c��/�f/>+ί��B{߽^�Ŧͷ�7�L�8~��w-Z$�瓛��mjj:����Gz㪫�j���<s^^qBmmmf}}�Rn�+O��W��������{�CkQFa�aI[T�L��3�܁r��ܞ��	�g�z*�fW��4z����߄Ğ �\��z�������"��bE4 �}��v����tZ�yn=s�B�)�v��k34,L��|�i���R���[�VKKs��K.^�����/>x�`����s�=�0����u���b5���lgQqa�Y�>��}<&s�Y�j[MM�n��o67����@�e _�fJ�J\KY��>U����e�s�>H\ٳ�+�a��Qy�B���y!�~�Z����{�fp��k5Z��C���I�D=l	x�(�Bu�B����C��c��9x�r�544�G�{��ttt0����Z3/�͝;Wtq+,*lY����o���{��펟?��G�9|xQ���IIIRRb�X���-[X}C�������o���s/�:��p�%���u֩S-\[�Y��":���;���x���r�6�}�S�Yxx���ܳ���`��? G������r3��#��ew� �ϷNn�uR��w!�'��dw�Uv�vu��½��!�T�C �yx���0�[]x�UUU� ������k���>D���>lT�-�PA_RR������ㅹ�������u6�Ƙ?4~t�z�ر��ŋ�����A�=p�@�Π����~��{�-	�����Ӛ��2;;;U�� �-�E�IFN��@�q�po`|̫׉��={|����x-"-J���z	��>�3��7!�'�aFWW����%�{�Jx�)))C��x�F7(�۹s�7)��!2z̭�s��!�#*�=t���G_�޾>1}���KD��*))�^z�G��ܾ��/�����uQDDhTb|���������������h(���+ޛ5#s�Zi�G�ʕϞ��nx�D<B��˞���dn�s����_|>��E}ܣ��7Z�F�9�/���N�ch!y<D�}uk��2���Ŀ	�=A3���M�M��\��x�:�9���Ѝ��- <w�tx�XUǔ���\:��P����b�^vv�( s{=����"��9
1W���q?��,sG��OKK�_�H��g�D
l\L�r�;=��V)#�u�Y����@#����9����\�˞��؍<�^L�\bX~��&V���6�x�o*`���0`Lx��*���{��A�����0���6�{�)\$��Bo!v;
���� �F��"a-W'L�����Ŭg�cd_�5��uuup1qr�11�m`����1,<"��{R����(w��fBȨ@aL�r�4}z��T��
0�����*q̘͗]|�>�T�4���q�֮];���ijKK�B�GO)�(O����v�ϓk��Zů���%?3��C�p]���p��pq��e�>s
�
!�����u�#�$�1�@�?��O�v�-���G��.w���=�vx�X�^^�Nn�aF.�fTݣo�̙��ޱV��10 <^�0��G�V�����>�1�%K����L�V*Ĝ~x�|\�F�>��.{�׏?�s�ر}���5��6�W�///_����h	�C�i��j���N}�
xH��mq�	��N?�t�E|
�S���MKK;��{�^HEEE��S/���{��! �N��x?����A��9<T�cqL��x=����1a�D77(�C� ���ԩS���3Ez���$;z�������p�·�硇HcǎȐruuu7�洵�	U,��b���!~�{�,�9�����"�EopM兊N�����D�c�$w��
�8���0�����0���Vͷ�J�B�9��l�EV�w�H�.���s�=��A\f͚%��|��!0�o�����׳޾^�V�ED �&
�0�^?턍
���C��1R�%�\�+\��-��||�I�t��'l$��f���s;;;'�K	Cx�
|���,�2C��=z�v�0�LF��
ꞇ��|ށ�u���Y�V�ɫ�)*���h4�������w�Ğ �\�%�9�-��ur�T���k��=x��@Vi`n=��x�j.Z�0^"��h��ֈ�$%�3����rs��{���I" �A��ȱ\WMMM��hػt��y��4��F0�����{{����q���sys����j�0מ?�<���۩�=�u��$.�A�L9hd�>^=V�s{��`b��fw��>*������;�W�P�����)�{F�{�F���)���2&J������� �����^+C�a ���U�V���Qb
B����S��@����葫�>��#z���C����޾�}�/~oŊ��͛��c(��wtow���&���^^�Nε˞����)���%��J�bA�!⾠�3%�X������!{n b #��>�&�	�������`#���=A�w��ի�r���r��w̉G���!(��������8v�7}�t���!L��=��>B��T�C��G]� �(���ʲ��ח�U���������C5��؏~�&v�t'���+��p�E�{���t*�p�>w�o��s��FBP@ 3Mre����J�"//�˔
>�R���1����N`XF�{�|��WIO?��%\��onn%�B 7^�[����0<�sT�˅y۶m�� l�رbl4�c��L�֋><~��zx�?;;ۗ�����y�z���?�<��'?�I{�c!''ǰaÆ%�mmA�i B����ˋ� ��eч���1�5�hh�;���G�P�Q^���y��{�j��x��x����"��>���̎;�7n���9.����(P`�?���� � Wi#�����~#G��W\!D
b�c�:�xD�����Ǵ2n(��98m6{�V�]{��{�SB\~�~T�q�kNCC�J6��!���@L��`��4�@��~�թ�"((�����7a�9�C���y�L)�-(8h7{�rG|/H�	�$++K��_����_^UUe@!���>�.j��[!����y��� zx� ���c_���ahx���Qe� 7��{t:�W�-_��mw�]�u��q�cK�~����r(
�O���AxO_�NΩC�e�?�}y
����f!�*5*�]n�c�F�<w�F�N����qkDE�yH�	�E��d�M�����!ҡ�%���A���c9[�b����X�.77Wx�W^y%[�t���C�e��#������T�ѣG���J�F�_����͝;�����f?V��4�B"��>�F���l�#{��llP�}C���准�m����%ϯ���3=���8T�����j4�ɔ��U��{���"n�ꫯ" �r�<�}:���nx�͋��ށ5�������v�[�h�"!�X��{K]]����;EO}|��{�6�sm��ޒ��;É�����B)�R�(�P�9�sh�i{J����BKiKPv I d�Ď۱;�۲���}=�nE�������\�T�ҫW���u������߿�c֬Yk
G������������+��A���$���x�L��G"'kZ�R�.>�F��w���j�$��*~�=��圽���6�m3sj~�����>GA�� ��a���'�WYVV&	�����C�jI��8 ���� q�-����q��G�^#r����f�����۝���҃=�ˉ��׭['F:***L����ȳϧ���9��<���e�dL�xN�Ώi�yш��ɕ���o�Ez8'4|ހ��!O>%f�s4��+J�9���O��>'@��GI�����<����s�������AOJJ���͕Ev�^{���O*6m�$~��/�w��b�ҥ� �7o�<�u0 @:t��P0���~�Є	��	2�2i���W�D��C�0�4!�h�v��?��w2�����FM�8#3]�����>y�x�=�������GB6�u[fff�PP���^A�s�����nҹ瞛�\�˃�}�A)rs�E���/1��# �>��@ ȯ����g�u�l�{��d��w�!+���"o������x��+V4
�80�رc�[ZZL�#q��z#Z���>�t\P'�ɍⵘ�W���r�2�#�!�hH�1���M&{ 9��7��i��Ǝ�#>(�WP���s�α'N�8/''ǁ�;Z����e(�9�9n�8@( r�¼�_]���a���׾-�/[.��y�^"�؎;���3^��v��U�ˉ��A�Z8ݔ.Īy,x����HX���U����xD_Ph	�Wυy1�)�l�%�`��fSMNN���t>%(�WP���/8���o�� �� �A�B�Pɛ0~����HB ���@ЮG��s(Г��k5\�ׇ6>B�h�z��%��>���'"!%����3�(Z���kBK�7K��>{�L�ɡz�٥R���n�pP�;f�8s�O����0�~��F�###�t:v���7)!�O��>466Κ?�۷ow ���8T҃@�����5kD��Z1w�\MU�<FTԣh�����ܥ�΀�u�^!H���E�����0І���뮽捯\����@NU�O=��$"�b�����6��� ���O���y�
z>7x�hjyZ@袧��W��N<_O����)�9Ft��§E�

������ם
��b��;wJo��^�v�$z�� ��h�"����?�	y[I[��x��|��P�!QTX$󺻻DzV�_(�2��3�h򠐑����Y"���\d����N!kܰ�(���F����9���̣lq��,fa0�Z�Δ�0tH��A����i<I"�it�����1�~�ʕR@*x��B(��F(�z���Ç!��իWK��cx�rn4"'�AL}�dP��E��s�ٹ�d��Y�f��P����������e��P�>n��#��yv��N��5#!5-E������Ee?�,���2��5�a$���!�ް��v���)B����i�[o������q��Y�+��F��y�u�G��d�-['EU�aI�0 @�x<g��m��曒(�g("`�6��fs���&�3���eU+���V���D��n�녂��7�yrVW{׌��>}8����D�N�[ 
��"<M�8$��^=��Q"h�1�pBa#����.�C�yR��䑣�Gt�o !�����|��c�hOFj�{ӧO�

�"�+(�F<��Cc[;:/��O�C��;��1C�\/����#��@�=nx��_�Ey����^Bhdd6YD*�=�� ��E:=N_k{KkgggD(H�!do��[��ޞ���.c��~g-���� �H+.k���h^���a|��s�C����b�s��p,�?�p:�2s2��§E�

��iY(lkhh�!L��,Ё(P�b.�q�7
�@���ݻWz�����Ϲ�xݗ<���8_zzz���!�W�����ߛ={��ǁ]�:���z�^+:��5c�#O.���D�>M�����1R1�#�Oh�k�?HƗ?1&���t�����RTTT%>e(�WP8������_y���۷�@{�Ƀ8Ǝ+�Cj�Q��U� ��o�!��._�\����dp�8�]�i*m�&�q��i3}衇�	��z�&�áQ���ҫ�z��A�ɹz^g&z����(��i\����[�����[��H��>t̀�f9@�Tk�§E�

�999���rO��Ly�
���5��b���<q��G�=�� =�������5&"����;j���~��m��=��BAC]]���_=2���?��L� j�E�Y�D��O���(���
��]�U��Ď�A�ܯ���k�K���as���)}Q�ԡ�^A�4aW\v��ǏO_�l����xӾ>�p�B)���y����ϖ��?�Y�Q���Q�a�<ue���7
?]^Y� �ğ��7�p�������ZBkn�h{��Y��n�{&e ,~CT/�7̉����@��1�1 F�ܱ������1��v���(����N�r���0���m]���&1��/}�K� �
E���eH@ށ$�#o�#D���f�M��A4D(>�Q�*��v�2m޼uv4� d�
��	�T�~��- ���0���"3;[���	��&���ȫ��}y{zO��zb:q��F��#;~�ӵ�9�W�L��^A�4���9�λﾹ����zTȃ�'M�$�����ر�� ��`T-���AJ�=��D�秣қI(.�*ϯ7�T8�cp�ĉ���ʳ����M��	˵�Ѩ6��s���o�ox��j����,�&���@89e���yv=�Jz�VkS�˽���X	)|&Pd�����������ݻ�ʼ�<ǘ1c�����D:����+d�8;;W��#���{L�CX}0Ddd0qն$�L����&"-�.����#G�L�,&R7#���i���[�~��-?���`�%z�^�}0�5R�Ez�|=0.���С}���9+��F((|FPd����������w.�}NII����I����~�x�c���_,���ң�\{�g1�p�����y�1�'�W:����;�ED�K��򈲠@�ə�������(�L�އj
'����\|>��'��k���rr�������*|fPd���c˖-����雑F�~���2G�ryy�rn=����G�>u0�.�H������dV���DhXJ���.����)8x𠧽�c1����z�!��x��s�G��dX_;� Eyd��yk�s���z�~}x���zͣ�>�W��o�L�D�g��A����g�m6��?�ޱc�r�9�w<g~ڴ��x��g�۶m2O/IF��'tn	���f��Yk�B[ˠ�@0`
��bE�������.#�	�FD�C�XC<���<���[i~M��E|�/��'�1�a;Q�^WaqXjU��g	E�

���}���~���f�ܹs�,�!z����.��@���_��� ��G�}x�<O�=Ȝ{�?^��fD*���&��@yy�������<)x���Ë�&��>ޫ?�7�SA��{�EVN���x`!h�sz �߸���h�

�!�+(|Fؽ{�����ǎ�>}�t���L�3g�+V��-t��ݴi�,ă! �t��*���IORhÞ��+vŧ��,�v;�p8�
	466�7�h<���Ϝ<q�Gق��b��Z�c p��FD����D[x��q��O3�x�}���
_�3�"{�� ��Ֆ���̜9{Vq�h<z\�1�f������ϗ��ꫫŻ�+��<	�d4I�7�̧tq>����2�0�#�v:��� �a�������m&��°�� ]����f�{����ǯK�����*���0C7D8"I�`4�P$,����	h�Q�:d���0�owNN��W����^A�3��O>9�H�ksf�N{뭷t xy�行�|1=/��pH��h%r0�5���Ɯ`,��"Gz?	�!&t6� A�����e-W
�6p��4K ����'�������&������;6�,c"W�) ��������ϒ��~���C���§�g�y&}��7͘6s�K/�"�C^m���/�)w���ٳG@I�HH��.I
]�]D�����
�vù^9v5����`��FT ��;=N�� K(H��Օ45�X��y-}}=D��D�6�����b��zM��Eq�=��9ߎ�=��].a6����C��6�(DF�`P�Q,�(�`����l6k娒q{�8[��E�

�"�����K�Z[ZϪ����b(�8o֬Yr�| '�!܎���f�B:(̳YmZ5=><|x�ɞ=�X��D�����^k(0:�	�ƍ�����q�.��:������Σmٻ�
ſ��Z��F��3��!��v�p$�����{ �Ͻ���C6�AI+�(�WP�� ����~f�o�^U�� �%K��!7��E��{�79��x �m�$� y�n-'O��ܱ^�'��*�qC�v�FJ��&��Cح���Bo�d��~�ߞ��%�.�H� �����y[ D��vڴ�S�mٻ�1ZZ_�V�gНT8�sr����l���


�BA�4@���§�7�xc��O?���L���Ўo~ڴiRB:l2�W��`T~CD�h0&Tِ�7H�$Β���}��s��p4��`�Z�:�����4���`�����[�ږ�A�Xw)cF��c��|��XK�%�{�I�&��e� �E�.�p":�5ԡϦ�鎦���j���i�"{��%�}��?�a�c���N"��Dব1�b��Ų����u�DUU�(..�Ă�<�D���-���z�\p��� -̼߽{w�Tp��j�����V1�A�n߷{�}}}�H�`��5�֒���K��	X� ��5��!��Bg4�(������v0L&����jU��p���^A��|䬗^z�?�����!3do���j9e�ƍ2?�7n��UEa.� z�7A��	�^>HG���h��*�=�_��Wŭ��'�����N����ܜFo?!F(����ݷ����3O�(nXG��s��V��������������Cn��)v	q�6� �����x\Ə��tN�+(�?�����u�)>��{�(fgdd�[��u����!���6���7��=t�S��<���нޠ���'�� ��m`8��Eb� �t��b��xL���.M�P�������q}}���V0�@�-�Z��	��2��I���߸1ٳ�!�5<&W����F[�3����o�s���i�"{���������E7nZE��9t��r�h��g�� z�AH�����{�Խ��a���w $���#g���tzA�PD�����N�4�ǣ���g�����?�x����MF�D�P�.ޢ�u3�,�5��G�:XS�%�� Hσ�Q���@��±����=��O(�sDS9}�N��p��^A��MMM��^{m�ڵ�l�YKɳ3N�0A΢ǅ���B�ض];vLND�����{/���,���=�!�٣�n��g�6�˰��%��AT >9OBb)ج�L]{[{��hll4������0��Y5d�����>��#���
{�ח(|Ě�r!"(h��>��dּxn�������q�]�Ǎ	��n� ++KU�+�V(�WP��@yy�sժU_�����d2��m��,����w�֭[E��:Y����@
�������A҆��SM<'�_�J���	p��+����=����	'��qLNN�a��=N1BA�p�G7n�8@�uԨQ:�P�>�汞3f̐��A��q�"ʶ�QYY)�Y��1 o&�@П���z ����O&�:'���dl

�����@���ǅ��kn5�ӌ�iYq����}�$A T2FA�q<(=px�L  yx�����ω����ٜ7��| ����28��),,$�1������֭۶~�{�>����tD�r?��"#=C�%<x�U�<,�v!����%��0�ൃ�x��D(�]v�0��F����^2� ��Z(?.�1���RSS�
��E�

�l�Pg��.��X}�O��K�m���D^~���#?��w"?~��Ǐ���{N�Cc�$q.�C�����Oa�d�V�����9A2���ڌ��8\�\���n�S��zoX�0�����|gOG�/*�T?@�;���E��>���Q"b�#��XO�=�)tL�":Y��h�3�Mرc��V㬳Β��o�D���M��J�K������x�j��i�"{��@���Ń��j��ڬ�����{�|�߾}��Ӄ����⎊|T�c�]]]�$} �y]L��ų�J�g�{���1��@��!�H���Xǃ��v��<T�׈��4iRpa�{�}���JiM��A�${J\�����h�i�o{z{�A�װ�_~���W^~U�޳[D�M�/*��ė��%i���={9�0fТ.Z;_}fv�v�w

����@��ꫯ������H42��t�EI�[x�6R���+��R�x�����͛�Ԭ�6F5�y� j�'B�1��ᡳz[�.;�˕ݲG�}��كXXl!c&���̴G�WD�P��e:Ru$F�ѣGeX�n�	�.�����_�����Dh���5(#^u�U�k�յ��׿��܋'�|R���O�.��iU��'1�Ӿ� '�J	�(|Pd���	 r0}�۷]RQQ��` TL�`�:u�,��I��C�m\��#���w�5��� �K�i��q���8?h�m�1˷&�鰷��G�4�]J����}�IOMO����buO<���斖E�^FBXKDV@�H�ȼ|����Hb��(+m��<��>�~饗d Q�.���80�9gp�x>=z��Q�\��^A�c �����:kϞݷ����Y�9&x�йG�ҷ���X��*Ty��[�l�3f�ذa�|�a�@���y�r�,��ЋlǋK�&
�D��7�����x`d ����\�g	�.�)��G�ș�7n�l߲}�i.�kC�s��a�"(H� ]����k�� t��aTa`��z�)Ҡ
��r���~<tP~�-[d�������o5�k�W��yA����G@���W�������8'���8��T�u�
�߳w���G� x�<��5o�S������N!�iH����MRY-F�i=�B����1���mq� ��r$��o�?Lf������	TS��U}��<�1CnSST���{����~ЄIv�����g�#��AZK+���0�@�F9w�s�HT*�� H�Ȕ��7��?@ ��`@tt�	��&�>g�4�P��DS��������6���$>'(�WPHB]]���G�C^���yO�x<f���у�Ql��:w�\����J�ҥKe��ڵk%���~x��іĄ�xa{� ��8 ���z%q�9�+���<D\p<Ρ�U�%<z.���cDJ�"����ό&�h��� ��"�(h���\��uXc<�>�t���djE�_��@� �V�555��GF�*�[TT�%>'(�WP�\W^y��U�F�9�.�����KR�^Zyy����������Q���E���\�#�� I3Q |�|1��^9�>ފ�~L�9d.�c�T;��!!���.ԃA�E]��V�{�ba����ڣ�i-r��uXs��#�k�'O�"= 댽�2e�ܳ`\���뜦a�|� �.p��ر�[TT�'777 >'(�WPژ��{�����]ta��葧-))�Ev���C��y �˂�����x�7� "����:�P�9�A� ��A+ �}�G[�3��\��'�y{�=��'�����=V�M���:�ȞH8}�����>x���hD8΄1��x�2!+�s0���O.��������� {�׿��/�w��@�'�o�n��!c�͈�P����^a�^��w�=�w���H$:�ݼb�
�䎪z�c�?./�h���

�@�K�,��*k֬o��v�R�%T��j:ق�cUy�9�,����q����L��Hdb��j�勃��!��03>���K�imnM'0���m߾{|{{�|��ԯ�k���"!9�EU8t�<�����z6����9)@� �#�OF�����r9�̙�*/^���w�Y���H((|^Pd�0�nݺQo�������&�BY}� ���o^4.���m������G(�x `xy,��cpCN!|��W���kgA#���a~z���蹭���wx��B2��Ȧ߅p��i�۰a��'~�BDE6�d	d������D�-��ɳ�9_�G�Oϰ�mxF�4�Pi���o~��}Ng�֬�^2�w�u�PP�<��^aDc�ڵY����q0���4����!t�q�F�w�#���W$Q@<e���Rv����A���A*��>���s�$��{��q�>���7�>Jd��3���
�@b���KD@�=�ga鉨�:�w���#���ȑ#�---�#ak	č��Q�@6�8�V�Tw���H��s��4 �~�����!:��i�&o��W�P#l�((�W� O�����J�o�"�Ԝ�� ��jm�Au��ɭ\�R���K�$�
|L���=-�X��k!xm:�#n�VK�qΞ���d.�c�X�n�{�?l�DB_�s��=0(`���ۏ<����F�=1����Z��A�\	�k��ȱ�±S֚�����>�B�!��F��c}��A����p�A���w�y��Ç3
��Z�q���#d�ۆ��DH=��P�O�{\p�UX$}�Q9Ҷ�<�X$J>�z����l4	��*<.������~""o�7h�RpN�	#��8	�b�h�sѢ��͚5}ǪUߛ����I�nĴ6xz������kD\��������S�Ayy������D3�}#���Dd���z����,����RT���e���[�p�p8�7x�Q�
��8�j#��+�H<��#��y���7	���Cv����&��A��ʡu�P=��8-V(�C�{� n�<�<Q���w/�xq�0/9�Ϲ�DH�nt��k�����;��M��&�1�}�R���=j �#��Ym6gK����kjj2��:���pJF��� R�r�x40�9�����sQ ��9��d��1�ɸ#//�W8��^a��O�S���Է"���`�P�5o�<yA߹s��9���Gn^!���=g�Id0H��r������0O��ki!w��>ѣ���0���h���E�|ii�")��j��}Zn��91�����" �њZ�@g��é���h��乨\3��ɂ���z��t@��M�9}n���=<�Z	2���
�-\��[((��Pd�0� �뮻�⦦�/џ��R޻w�l�CXy{\��ţcly��̙3e ����3�b{{ \��㼈
�.�0����er;�ϳ'ʕ�DZ�/~��0���������Ԟ�^�a`��`R@� ���"����Gٯ[�ζ��si
е��=��Y�`��q-�h��������L� W�'��K�^�3f�f�[�W8#��^a� �9��s�܊���`3� uh�C�}��PLC�0{�l�b=7<h�rq�G�>���P?��0*�A� x�L4<܆��8�ϯ���&�c��\�7����l�͛�Q^���f�ǘ� �E͘����/..�y�zMb`ǎEd��Mkj�����}@>�)HF�N�Ox�X�`((2�� d��C�L�ɡ}����������BA��"{���`��7n��\�`됗E�<�S�s��zx� 	T���>�@�9��'J��y(���ʖ��)�#dY\9΅�ǫ�eX�ivL>,��ae�zmw��۔	����~��]����~�ȇg��9<���o ���f�8v�q<��Da�۱0������̹��.D{X�=x>�����0�l�SSS�ӿ%��p�B�� ���?��s��|qss�sT׃ȋ�9r�{ҤI���6'��@Ax8b,8�y y��Y9d�-Z <�g�Z��e%=��s�����0r\��>*o !��GD@M\pA0������=1L��L�>�����9���zbt�]������b������^e���{"��ρ�1���dy\����.4�=iD�Vˑ���BA��"{�����g��?v5���t�0�}�'N��ѭfժU�x��/>���@��!�Cˋ>��!�;u���/�-�?�a��#	�Z��Fx7��%�B9x�f����=�>o��	�ߣK Q�O����T�,t2,BD�^z�d>?���I�|:������۶m�iii�F��[&��,t��hE������ᝢ��D/=�S�5�|ra��Zmf����B�ꅂ�E�
��W�v=��_Cg�׮G���ɓe����>�ǽaŊ��o���q<.�.G*�D���r8E��bI�}�b��]"=%U��hJ�����e^�{��@a�8	����$�P�����&���<D��U��M�����?������1�y� �K��J�{�.QP�'220��i���������61�y��_���119��7T"��ޘ�W`4�d�C+��P8$�����T��!���ǡPP�8jB=����}�ܹsG�:��Є"{�a�\�ryvW�� � �lmݺ����~����3���p/µ�����e���Q�����$�9�g�_zIV�]zը@�$Ώ>�cx��p}��v���WT��M��#ŀ��
|��!�������>q��SȄ���1��;|�nHE$��RS�-��7�׷g�ܹ�<Z�4���#�Y�ׄ2�o0&�Ӣ�O�ɟ�0�=g��+�q~�ö��zTᇅ��E�
��w����C�Y��եÀ\��\�{��9����x񂣿�ݓ�t!7��Q����$��8(..��:G��jzhwc%5 �5��L�A�����#j�6�uvv^��d��Dx�{��^(�'l���g̘�Ͽ��S�>���k8=UkD�  �63<#Ozj�����APC8����x6�v#�,�Gt���>&K��5��n��@j���?��Q����x��+����777Wy�
g<�+[����꫗�]Do�C����������<�߭Y��Yh����Ё��G����Mk� 0���_]�1�?�Q��9z��<{��A2�v�Wz�1�3g����u[�(�L/^����&�|��^����]�hQb&.}~��������O�q��@�R�-.�˟���lN��n���0�t.��+3�7��CTk��9�5+rQ{�R�(n����"L�8�G�r>���h���YO�PP8á�^a��駟.����voo�h�x�@�(�>��s�7�xS'y�5k^��.�鸈��j�޾^���.�z�8ހnI 蹇��mnт��P �@o>�d/� ������+�m�׋�3Ӹ �G��=qv��uyǎ{�~N�k433����%c#�#<����xx���p��ub�����ݵ���Ʌt�}�^�*_������<����`��u���g^O�+bQz�pNNz�PPPd�0,�6�o����F����pG�=H��^�3f�sW\q���~&����Q���e[���D>w�\���5y��H�'�xB#�8h$nJ�A��i󔻈֦���s_��k���ߗ��.$�p2�� ��H���0�-����뮻���~&/�gϞɌ[Ȝ.�ŉbb�Νٽ�=e�F�W`<����8E��&� ��{���ϣ�Ye/)��6��! E�
�555Y�����>Eёg��+�Y�s?�裏�n��ɭ?��/�K�w!<u\�!������4i W)\����߲��H�W�Cr�l0�d@���A�F��w_qŗ��9�_��Nz���&��@ 0\���^RR���ºq����H�\�Ć���������:�OX��a5~U�/���J�w ����X&{���Z'
����p���	"##��<��G�wWH��Ac~~�eeeJWaH@��°Dee��P(8�.��dnAț7�z�U_{��.kX�~�����Et1���4.������������A��W��}���Q��v��ᱨ8OWw��;1�˗-[ր��}�����qN�t�8/���322�%'L �O �!i�a�}|_��K�8��L���0b�d��C������w�#g�)Yޖ%p���`�Oj�y�4<&z��c?i�C��[&L[>\���+;TWW[n�m�e>�`��@~PE�|t׮�o~��C���?���<�Ѹ�O�6-Q���ϗ䏰:f؟ι�Bi\ֲ�A�(�����B�$�<a�j��<O#+%U���x���<s��qb��������a������9���¹`|�\��D�[===�*g�¼o�q��4�n�$f�B�'� �b6Ya{.��6<��c/�������n
�OOO��r�:����"{�a����Gg.�h�)WUU�:�;==�D���O���t[].�ԼG_=���ox{a�?�0�DΤn$2�*z�<i��p(X���B�a�1c�v:���7/Z��F��s;����b��n"$�G#���!U����y��d�	�b5��P�F��;ڏ��� b�;+	X{��������}�� .�c�c~�N�5��zv�;vX�1*O(�WVصk�����%t�ϣ��9[��#��������Ǽy�꺺�<{���Dm��=zT���'fw�y2�{��!Y���1��9���|����a�6�xcD���Ν��+۶ms����1�%,I�V��xxpz!����YZZ����
ٛ����xx��p8�z�.Q1�@�-���s&�>�o�����a��N��_{�X����D�Gv V��	�&}����ә[�B�
C	��������⿈��#ú E�\�\x�[��~��e9�%��®��M�B���P���8���H��˹�@� �����p%��DN�dff�7n���{�������Bz����%B˜�����N������_�>777D�ޏ�x�u�,v�L5Ģ�.�d�v����~4������r�`ر���-#��)ޏ�Ev�&�ēy-�8&z����rrr���:�����"{�a����"�qmm��@ƸH�'����}�s��m�qZN��"GF֢�|;y�2$��<�7���;njj��B� c�Ճ�9d��ZǏek��П�����zQC���p
����#ud�~�?�+��K��Ii)//�|�O������K��mw��Ϗ� �`�x�/������q!��|Z++b��w0�x$����Y��G����{B�Hb0M��V��SY-v�T=ztњI�&���"{�a��>���h�J��;&�^����۷���n��c�����<L�����GqH�:��#_���+/� �Ǳ��8.�����Rp'%�vٲ���gD�o�=���Y )&h���~���\���Y�W\qſ��B^�b�`_O_,�q&D`�]bxy��,�{;�*<���O^-ooH�=��W���!�1�~���*|�G�VCt�=;���Z����"{�a���Gkk�z�ƅ��������e8|���K~��eD�T�[�.!�)\L�{����4@��omj�ab��A
�!G��d���'�܇ƌ������������غu�l�,Y<��@6��� ��c}�����D�a-�!k�\��z�` ð���L�e�w�͖q��� ���wh&���m2iy\��^=������Rsq��
辻��`�)ST_a�A��°Accc��A+��A�ĉ����9r�Ͼp��ϛ��.�6H�2Q��A������p�)[�� �����E[x:����O�V���;��4d����&�2p���Y^�dOx��>���~/�>9Ϗ6�=� 6��+b�0~Y�ڔ��\�R��<F�
<ϳ1�\��������h����O��á� #ڛ(���˯�J+(	(�W6ػko�@�ot,޾~��Ţ�X��������?��g�?7�\��U�(�7�PT�&���.�sDg{�cH �=H�o�+��:=n���.s��P�h��sΜs�qc#�������;�x����mfE�P,��F��"I@��	
χB�62H>Q�.ә�X�q�����8�������t���x���F�A/��B�F@�K��7��2���A���Dl8����f�1�b���eGC{���m�����
_a(B��°AOw�2OJjZ���4-�������{��ܲe�SO�~�y�g��:}4,�����:.�ܶ�V.x�ȣ��A����H���~�+���x8��l��7/���F���_Wf��g���) 4y�Q:߉iӦ�?���wDS�.�N���w��?�70��a\��@]���O'�ͦ��/:�xRő؛`@
����(Dbm�7"6��9��
\�ǅ�:}L�-2m�������
5�VaHB��° ��푇��v��9�����m���ZXX����7��!9� 1k}�~��� 3�;;�E0�}���sT루���³��t�Y���M~~��e+��>����:��j`$�߅Ea�x�?6k֬�%h�,\�8mg�j{��x�[�y.���YZZ:�G�~������Ydyx� O���fx���=k�LB�`#I����<<�V�l4��~nQU�
C������q�M�|��B���?''G��=���ǈ|P�V ��t�A8#���2H!�.�'H�.#s��yg����S��CA�F�|��0�`�3	��TO�'��;::,��}9�t���=U����>_[��C~h˾}����[J�n����a_A��A�oբ:�S<v �6�.h��<�V렽�����@�u�qO{�����&��0D��^aX�����.�I \�"������F��� vx� ��� �Ç'�� �- ���v���钄�gу0p>2
�3�s�̞=;A����楋��X-V�?�O(�aZH�QK�e ?T��477{{{�6�-!̃4��y� ���z{����!]���o�y1���d��A�}}=�#�}��5��ܥ ϞC�h��M�7=����uQ��-�F�~��z�PP�Pd�0,�Jl6���J��h�'B��E���-��������Z�2��牐�1 n�N��AL� wL��={�,����11"����ª��nݺ����,"{��ᔡg�����N&�{��O���n��6�ɒ�A� ��=�x�A�+���:��׿�������Ѕ5�;4�� X&nV%�J|.ZD��卹=�+��X�Q��X5jTA�PP�Pd�0,���ta6q8��r$.��^��j}� �!���~NN�4��:�����Y��|^"����^+�C��_����w���gʔ�W��ﴬZ�*�7���R�ɜ� ����2�td(���h).���~���w(���=΁����d/ d��7��GCCK	�mi4���1�p��oliѪ�9Z��b���	B�\�g0�N��z�@��1�v{���|b���P�"{�!�w��_��Bg��2�]wO'��11c�I�0&N,�>�|����gAqOA�����9a̺G���E�$i���������tãFm��׿��֯_�����6ł���{����y���DA}~x`��N��mw��5���4������o�9��H�M����Oa`�џ���E>�`6���{��b�":�Sf�'�q+"֊�f� �F<r���[[VV�����O��� E�
�(��s�.�^�1c�l�+�8$.��� !����h}K\]��eO{`�_�����/_.I�p��&��t�� ����oڴ����2��������ɳ7p� �����#GL�!rss?V����Q	d�Y<��\������E������[�������$z(�`d��AZ����i��X�����VE-�oL�<p�s��'�U��g�cZ�PP�Pd�0@\�7#��Xi![\��������F�-[��|;��R/�)ρ0�<�>x�\���?&��A�{�����[T�c@
������=��ɓ&W�7.�_^��߸ 7q��=N-ݒ(�w�Ϗ555�ô���߽{�yǎ�9DPf�>?~�4XP���Z�[�������r1$#�(���_C�����@r����oX� ����}9EQ��" ���6�6I� L�6��7�!E�
��b����m�\|��;̢G�~����
z�1o��r�8ρ�A������<=��A��y���x���퐤��8j�Z�f�V&9��f9xh����$B��(�{�r ���L������G?���(q����\c�~3R�p�}X���;�-/?Աd����׋����
Ӟ=��o+v:�:4,����&��v�S[� ���<�H"�r��m|�ۉ���w��ʆ|����"{�� y�z�u'�bR��s��&M�9mH���+� RS=���E�;�؁�a  � D��=�d<�x�b���'ı�u2r�9^z_����:�x�#�߬�F�~��������k�����@��O��cɞ����6JӃ24�߀N"������s�;;��]<�U<&�$6nܘ��־�$�
{�;[&���m�:���t��v��q�{�ТA��d5=:�����1c�&�^((U(�W�E"1��*|G�G�|��-V�$Cxy<Z��h���^��5# }�x/޷m�6q�M7���<�_�J�v�g-��߿pᒍ+V�8%�Ku19��Pl�<3�����s�|���蘏%����2
���V����;%�y!"�="�@zz�>2v����={&�i�6�}(�ľuww�ܜ�IӁ�OII����s�$����w^����)Sz���0�"{�aV���=�=Bܗ^z�ػ{��z��}OWbh,��}ܒ/�}��b�̙3�ڵk��_,&N�(s�K�,"�:_�^��O�����N�g����|��W|%���_�� ��3x�-���5��;�s�=z����|7���K��2�ш.��@F-�5PUU%SH��ǹ�-�_UVV6$��6l�`��o�\J{�	k�5����A�6w^[*��'�.�cOk/���ȡ|�?����P�n�陙{����E�
��X$ƅX�߱D_5<�ˮ�B9\N����xSS2$��|�FFF��j��R@���/�8(N�$V��<��S��w���}����!�7W��|�Ё��- Cɨ!@��	��}����z�>"�f�1���򗿌߶m��۽ހ�:u���q�w�qbC��~W�����˿T1TI������7���������Gs��a7I�`/�G�b͹z�g	 8������:T�WT/�	�+y�ڞ�Z�����i��s:����<��L�Mdk�0Dh��́�녗^YY)�F�2*�}���d.��W_}Uz�ȋ���UW]�я~TY:a\��~�@�{���k#��x�;U��"����UZ-�߁�:F����s/h��O��li��tӅߢ�K��Aqq�$@��{��W����c:�;J^�'*�� b���'?YH���6V
�:a��,��S��>FD���.�K��J` �g���޷٬}������6��0L��^aȃ.�:�٠����H,,�VSbj�Ao������[TU���(�9x��,Q�Cq������cnEE�0[�◿��x���C=$~��'!������;=hc/�D}��6o^i6���.�q1��@8붭d�X���O�*,���C�5�_�/�~�_��������7���Am�U�qϟ?_z�����X��DtC������r�رgi0���~��G�(����c�1�9|��d�ҰҌ�݅$�k��"BW�?>�H�q���;v��p�0l��^a����̌�ѣ��d��Z$�y���'f͚%6o�,*�u���<=H^#dp�ՃL��@��?a�x��g�}V\��bժ�Z\�\�p_ߠ!�{���_�F�����B�g�}��7��2���Nt\4=#�Xnn�)R�0"���"��<�[��@����wF����Z�Zc���]7�p�ko�{SE�ڵL�B��f� ���)���PP��O��GC��&F�~�����kCs��z�� �%�r�v��U�S�z�aE�
�Q���%yƋ�ሬN�����/��KJ�w��E��ߖ�q�CN�����<AM�QQZZJD�F�>@�ҹ(��Θ>K�:,�o���;0p��<����S!�\��k�e4S����&���3sJJJt�=��d�@0 R<)2�Od���8B�=���{���g�y�n:&��kʔ)�|;w��0L�H������Y3�v��W�!��/��+�|�O=�yc�`4q��߁�>c�./|��"	A#D��|?a��qn�����

�"{�� =�z/��>�%�@���	�{�c����i3�	o$�jo��A�𔳲2d΁s!OD-���^|E�r��bӦM�Ç+κ��K+SSӉ�Eh��]eU���q`ùA8�sG����S���E�&����&ϴ'#=�n֬Y���-[��]|�%�FU�tF�8ߜ9s���}�6�}A�h�i�G��*���֬ys��ؽ{����s.�^=���O o.j�
c�x�L�<����>�<�8�Dt8��s�v�;���

C���<���M�Ĳ9�ٺ��va2�7�/�2��j�裏���뢘�sx^#�Y��I:m
�"�w���+��:d����m�v�Βz�w�q���ן���ה��>����*��u{JJJ:�����@gGg�/��mm햮���z��;����1cc��g/=� ��!{�E_��-.,,� z�A< 0�m q!t�����}����~�k��FE���M^�<�mf3��� brN���=�3b�XHG���" ��w�^H��:ݮ���f��0̠�^aȃ� s�-��.��=Z��oEVf�,�{���Env�$l��dIj�<��z��9� )���x�qI ���z��ݍ#B�t:�mW^ye�_>4�Dc��D"����C:�n�ׯ�ڋ/����գ�L��A�&�q���eZ~�����{�}�8p�2>\c#-C��{�񝠖��s2@�����˖���!��o���>��(�S��{���,�Q!@��K�^�hiD��z�-/��J�A݉W�w�gf�=묳���°�"{�!�h6o�8����d	��1�!Y.�����F�cZ����@a@9���aQ]]+C��s/۷\.���/��ؽ{���ν^o����w�������i�n�m���q!�����W9�x����~�y����&��f�0��a�Z���[[/��B��}�m�v���"�RH�3`޼y�C��¸��G0 `�lݺ5x�%���o\����q��x��]55��BA�Y�D�|=�!�oֶO�c����iam�Z�����tD�m<�!c�b��ҝ*��0��^a������<}��EyK�,�a�,�;�D �mTA���EmZ6�#����`H#��C?�BF����+lV�سgy�ex����o��C������i۶m�:}�?�_]]>����կu���.0��!�gB/��:��#�H�H���/������fw̥�a �!� ��{����(<$c F���r�_��_��oC��]�������9��b`����Է����k��KT�#���?�<��?��7p{\[Ǝ-:*�!�+Y���[�KF,�'��Ē����C�¨���􋜬�q�D�������&r��D8�Uk�([<��a�>Q��( "��A  [�񄴽{�B�NG�@֚��Xo�ז����1YY9���?����;wμ�� �ߵk���뿙F?A��<m��z1!���?��K/�|#��tz΀χ���: 08@p 3�l�qR~�"B�����8CV�֭֊��h1	#���~;�^�A�Sʑ�M����&��>�ɶ�����Ω K�!�3R������ԇ���	���$�mn:V3�����cƌ]�͙��"��ĉ�.��(/� 	�a�k��c�M!MT�'�?��Ri�h��!u�uT�#'��=T�PYB��,�  ��Q䠝��
䂢<y�Q"��߿��������/�477����31 ��mٲ%����˯�^}9}��j5d�3eg ��E�50 �]�=[ZZ"۶m���/?~������dDyZ[[����Z�{�����<����8���އ��0>�����8[�N�ٖw,%���PP�Pd�0$��6y�)taw�������uww^���5.�p�q:�v��������%��A�i��ĉ�(��;�� ��yh�[,&IzA__�$T�����c�}k�Q�uu���>��@2 o�#�N�=2g���9��g�������윀�<�|������42"d~�����I�^"*�6D`H���9Ry�E���~����o���+���A�ӄ=�aF<0�ɜ�ay4-?��	�{�[� ��S�(O�b5XTT�$�)�+������f����5��{R\�ğyD춘�����ȼAj�c���o	�X����$�B>hȳL.<u����ɕ�������AVNKK���b:y.ǁG�ss�<����������7N�<�|ӦMW�]�L�,�*x=�w�� ����xF
��Et�>��wp�ƍ�s��}���{S7
˶o�6�8��ZtF����:&|��sZ�}Th0�`�����R���Tϋvfddn�:u�PP�Pd�pƣ��elwg��F�
��h"g]o������H�1�i�Y��Har�$���Nz�ȉ{��RZOo��h!ވ���%2�&�<O��$�}����H;U������Y��4ѽW�ґ*��1{�0�Ճ�A̘�N��|����z���h$ZH����| �d�^�=<�D��T��2<bt�A��]�����O<�fb�c��ծG}�bz��<Ĝ���d/�x����/Ya����� C,b6��KK'U|tb���p�"{�3���YN�� %�m���2�
sxhG��dO<���pӽEd�d�E��V����x�W�Л�&I� d�(����"�ǃ�iiG�{�2��T�xR��Ճ�qz����-�����UjR����Y:�����ލ�;�$_�y�����e '�.S�}r�-��=z^~����!�喛���A��P�-W�Z5gp�?��Հ5�n
<<��1��Cl�.�CąC���{p\ M��c/阾�TϚ���BAaC�����;�B>�b2�bD�XLz� W�G^x�̭�\��zT\�
��ȃD�Z,6"��Eb2<O��dtBg�B�w�����,�~���|�ŗW���|���C^����+�I��.z��$�cr�<r��5U��$��f�7�#<�� }�0�"3�<"x��@�xm���Q"�n"�mii���{���7��Ad/�֬�m��o<�b����W������X+�'<������aH�:{��O��Ţ�HKAQayYY�*�S�Pd�pF���3��(sX-&�REj�k�Ǐ�I�wh�#L�כe�E\~�e2w��Ҧy���:�����Ga�Y�ۃ'�^v"�O������o]�xeݹg�x���_��ko���dB˻Y9�3�g�����QF�;9˸r�G4�3����B>_�رc12x|���ʱc�>��q���r�1��o��1\������u��� B��<�ֈ�ϳ@��l��Ғ��U�x����o 狷�E�SUa�*�W�Pd�pFm�U�[Z:;�B}����������Č)SEw�8��$�k��A���q��K�,���D�vI�~�����Z��@X�R�Vze>����XR[_�7�2]����c�),|���k�]�Je0�����ƹA� ~A�t���$w�g��H0.��-|2$M�!��M�<9@�n߾�X0�6���9g�<�@��ٳC��z�N�
�#�<2��b���Q�`�/ג=w�O����J��8x.--C� ��j5p���ǚ��J{�7!��~��4t�aE�
g4rsK:|��_zn�ٻvo3ۉ\}D�Շ��8�b�¹�P�;&'�բ(O�������d�m���0v��J�<x�N�C R��:<m<7zt���O������}G�T��D�����Z�$p���(�h@���A> �� ��6MM�  L����Hb�*�����B����o�}Ϟ=؝�������:������+V��y�1q��+�&�����.�K^' ����NN6�<R)��~Ќ�D�u����:u��Q�Pd�pfc`����Y���}ͺp�\����4��y����6���+&L(��M� EƁdNH�	i�]�Ñ�0�uR/��w]��ܬLǳ���N"�hOO�A��ܬG�<�E m$��B/�B����X2��ֶi@D"��w��h�ڲ�<f���( A��q���.gE_o������l\龥g-�����_�|yd(��Oq���Q���g�ڹ��5}�_����9&{`��x\Ҁ�Ϧ�{�jy,��=D��j�(-�]���F �+�����Ni车�D�]����>�{��"FČa0�hL�E=?�P�wv˰m��M��Ou�ǅ�o@�,j��N�������B
�ȃ3Py��$@��<aH��Y��}�Q��r劷
�F�{{{ct�X8��A���ys�wF��yD>z��=zt���ޅ���UWl��?�`���'F
P�������)���cM9\�^=�}��y�G�A�S�+�Y�7 n4x�
׺\�;����"{�3D����7�C�����<� �и���x�ͷE(����lq�X�x��e�}A^�8V� �{�|�"RS��e����>a6DsS��O�O�= C� ���\9�.�a9P�@& ��ɓ�����o4�t��w=v�M7��B���j��{�.��~(�o���m�h2�y�����0sD
�����N2�.���P�~ъu�,�0�su��W�c�`�q�=֚[�p�.��k~��q���=[

# ���8�b]��V߭�H�{�>�\x���'��TMl�k]=�"#=S��o߾�܉�S$�VUUˋ?��A�	�X[F�M�A��|B��yDMM01/sxT�L�P|�J�+�c�'����nw�ߙ2y��w�s�s_��|7�|���������w��;0��x"�q�����X���4�+F(ȸ*&�~:�d�5pꓥn?�8q��AG4NKt9pk#�U��Cz��`NN�q��0B��^�CGkp��7p�ѠˈFB�H4,rs���~� y��r ��E����q�P������˖-����EE�A�M��]D���A��%���G46�":z]L�C�D���"'7K�*�5=��Ύ0�|����ZZ[*�L���o�|�o���Oʫ#����d�O��~d����#Ԍ��4�h:\VVV;���{�%Gye�����43
����"�d�1,ج�ٵ���^��l�&J(�%��(�f49�ι�����р�6�%v��wu�twuUOC����{�?2��w�3���l��P��ԼB�\)���<ʐ�]O�	E)��@�(�RZ�{�s ���- ��`����l9`��x>�yN����hGW{�-^�Pi4RQz���zJKK�","��'���"���AY���9"R*�#�(��gɩ��L�>E�_�~�����2����G�Ϯ/.�GKst�\tG��G�����CtԄ"�y9ٻ���ʽw|����XŽgϞ�g�}�z�N?���*�)�@�u%%c޽��k{p��������W�ԼQ�$ �ޛ'|J�&�����BU;�ׯ�����"z��4���v��hqqq�	8�s��[��-�W��e	1���I9��,fF��܌�1�^WW+��̚5�INߓ5.�޿��2�a�3�S����G�R�ҥK�r��7Џ�t;�G BAa���)�O;�*�
K(�\v���<��G_�	i?��/@����r���=x�����L��6�l���BWwG0������O�?_+��0��'�����[�'4���׍x(s�e�.��JJ�Q@�% ς��9{CAݙ�9��O�����q��uI�U�9s�n��q>��=��	���􏋋�/�j�9�	�I���)>����:��َ�S��=�7n����5�\��]�v-���PYI�p�1򈁺���[Q{괬�Ǎ�@UU
֢��[>܌���g�9r�:��!8\i�jGvV.��[���W����G=�9�[���������`�g0�(�@���J�`�宻��~�ر��^��Ç5���S��h1��+�D�� ��e�<A3���N�'��ɧ���z� :'�*��4Vk�`VV���L��8�s�A�q�X��t� U(F0���=$W���r��:��lݺUN�Θ>/��<�>$��5���{����X�h!v��	�Ɉ�{�� ��O�]�>ڲ����v��n���g?�oi�Ν�^�b��x\j�����j��Ͼ���[o�{<�����O�뫮��p�u�mݶ�>�J;�괫�d�6�l�A�3c�U��^=���)�����h4f���^��U��j{�<����O%B� ��s*�T���)�)���Wj�����|�}��~J ��N��'�vKӂ~�!��
�)RJV���1rږ�ښ����~֬Y��_]�<GmU�@���?�&L�'��^p����@��K�^�e˖�n{�N���Gh��;x˗o����L&sY�S��%���rs�d}qk[[��}�����ʕ+[�4<����E�p��M_���)b��gZ���.�?%��+���Bee��c;v����Mcd�U����+�'��[.�S�Fre��R�#�z"|��n�yt�='���E��X5e��>pp�g�d����A���kM0�/���nw?tZv����tN���:���ӀBC]-��Z�
�.�D��/+-��먠/M.����߾�?�<n��&dg�b܄q�Дe�/Ė�>N���=z��'�g���Z������>P&�XB����==��y�����ڵk�}��7��G�馛r:�;/	BN�2��HFEʒn��g�%�B���v�_�-��s�WЖ͍7�8����6�ݭRAO$��J:c���)�u��*�L9&F,�	)+���c��@d�ۭ����B��8��ɞ�Ԟ���:#.�W�:]R4"d
/C ��?-�T��k���5���TV���o�����>�?���<ٓ������4< '���_�<� �͛'o�l6����D�V��fɊK?�٬��������a�b`�#��d0�O����W�ݻ�"�ZCCk$�ágd,))VA�����CG�r�bD_{��555ن��f���F�������+�b�KPH��OJI�u������d��I��_�4�,`;v>o�p���d��
����y.�DC�L�������_�#A�!�q1���*A���n�4�)4tu�b��ݘ1}:Ɣ�������	��F����5��K����~ʴ����{r�@�t���JKK�
�^;v���n#v��{���G�7�iW�V2��{�>���CV����mj�آ1i-d�CcnS֭T�m���Sf<��^��|�u7����j~��عsg������)S2B�J<=ɑ=�� "��=Tp8�r����W|��@��NP�~�n��3fL388�Cp���_�s{Z���7խ��h7�ٛLde�A�7bh�^�L����Q�{�n̝;"Srm�#�
s�=c*TL�M�6MN���ף�� ��RA_<�@$C4��ي��6���M2-Y��'�T���6��G�������_������#���E�y9[`��10���j�7���S�0=�CL}�W1�g<p��(e�`�#�<��}!���W�9AV�ԺrLI���o9���'���CP���)�׳g�,(�5�|788�Cp��8g`��}�x��L+_��$� ��:'Gd�m�l�����[+4B����[n���	;�������GQQ	J�Ɛ�^z�E9E^9y<jNVc�%Hgľ�㏑�����t�6�2�euG�x��݈;��NLX�Ɛ��!���22s�7��gN���կ~�Ю[�uv�\��ݵD��g���V�G4�Ɇ�/,
fdd$㱸��q���0u���>�`7'����S���yQ,&����Zr[��a+\~	���2���H�0�����2�>m£)�S�z��y`ڴ���y���'{�s����q��ַ��]���EW\�X\T��<|�-i��Ӿ�h�M,+-��>w�l���d�&c���fԟ�Cqq�"��/�z�-�؝r�����߿�"S�6��;p�uס�������˕�ꓧ�uۑ��-��9����)��a����_�o����Xв��W^9���.�y}W�Ñ��[��pD�HK���d2��L�Gع�&���/��ꫯ�����=��C�Her���I>�oS���Ϊ��W
��JG�R�OΆT���&�)�y�{��At8�G��2���8o�ɞ㜀-��7��WǕW̚P9ް��@�����w�)��-��ݭS�Fgn�jLY6��{�U�P��0��>~"�_x֯_���Od�������
�V�+�\��;v���F��{���w��u��eB�<y2jkk!&y�?-]����q�;�v�&�7�W۰�U~suu��[�n�x��O*��P���1���hT"#��Z�`��f����3�<����y:��XLH��M�b�����G��(���'O�%��Rz�O�>���O�a��l������ޘ����9�:�B��پ}��)S�}xݻ�CǏ Q=w�\�֏>���o���nG+S�c�k�^�W�p9K&+�WRZ�#㐛�/�����i���B����D�I=u�+W��xrқ9k��
�`�fyߖLv��;�LH7a���vc�ޙK�~�9R��y��g��{��Gǟ�O���Xt�~e/|����bV��bWnPE���On��{��@٫W0:0�`�IA%�fd����N�g�N���{?�����sg����x�,_�Ύ6���b��%��e+����٢��g��u�\�-[>Duu��3�g��a0�A��.�BV��7l�.��ys�y�f,^� ��{�l����mr����_���,\�GW!�5M�8��i����6_4��ߙG�Y��RLpB'���%�V�?�cfH){e����p�]��.��i�*x
��'{��
��޳gƾ-����Ю�r12�)�7s����'pӍ_Awg+Z���%=-�T9O���M�?i�$����eE�w�^Y�_��rD����������l�2��|R�V�o�� =�ƭ�k�+��O���}�؊������򅡽�����p����I��!��#kq��~t��qkF���	Jk�g+��`���}wq�O�����;����9�.��r�{s��N�~|ie�0��d3���	�ٹGEL�0�}��t�mj��2Gd��L��b�V�c��c���[������l߾��݈o~�<���DSSNT�¼ysPRZ&��-��ǵ�	?~�G�|q��J�'�3�k�bb��������/������kh��ș�s���)�<E�+����n�͑	�O��g�>1R�GYv�M��eecO�>��N�g�6I��o]�q�jօ+��Z��%�Bȇ��<ԝ����DSs;����x�t$��`F����i����w֮��jh����.b�����UW���lD�@?��0#�b0��w�yG&��˗ˊ��nwR ���z?��u
_�mۦy���gF"�
"h�"�N	ڳ'(����M夊����(���F���+�Ur��&����'??�{�s���d�q�P_��Ě��}՚LX���ƬU˱�?GɌ�8��F\T�`=#��q�Qs"��S����I��K��vtYz�1e~ACS�L��ݽ��Č�r��땕�ZP�tm���o3ې��d�A�{��k�\�So6�U^>��/,p3���Ng����@�n�]��P������x�(��p8��L:�A
(HT��*�A� y�3t���(..��8�{p��8+��%���ܽ���g3
C'�pD�"a3�]���[��s`IOCcoZ�[����@6T!�6�>EZ?��@% LI��pJ����x
���#����@R�m��n��رm;Ɩ�ˋ���4p���Lf���%���B��А�Ŧ��~���:���33�(��v:��'eOϕѵJ&��+ǆ�_��uu99�m<����ɞ�,�����=��.3똞�A�"R
C���:�Au-�.� �L�ee�ap�j�zxQO�$�^�	�;.��<���V_�Z��ݶsZ^��;���.F��;a�Dy�A�O���36i���.���p���cG���¡1n�[��j�#Cj0*���F��+�NDOY]O[��GDO�t��LIJ�ع�333�����d��C:tH���%uO��4�Zs���d/�L��$���9K.@�͂H�(t&�ly"����O��䨾k�V��'�v"��#���+@�i^y�Ԟ�����.̞3v�,@A^�������S�O?Q�W�LM�`8�P���?{��X,�A��(�4=�`,.&�d�}t˝������r`@cp�3���F<{��E����>8�s�lx��y���n�`A0 ���u�
���D�Xr�eP�co�If=m�"!$e�.Q��*�N�g��+#}� ��ny�F@Br�rI3�(++�g֓�>��]|�Ÿz�9���ځ[n�
v��ӭ3�_q93����8�P|��%M��K��)S�ݧ�녑��B��uţ{��!Z*�����93	O�������m�ƕ����C'{�Rs���[n��O��I��$���[��zF�Lɹ�ʱ��I��dZ��`d�uj�7zbX�I�{�
#����&	�j?�'/ --is��<q�ܞG�:�+�J�\���|������VpS�/��պ_?�����풧8��w
GG�~��rL9�*�[CI���k��~��<�ō�EE��̙��+98��ɞ�����K���U�'�N�#ЙL�"4Z#�l��(�?�:Zq2�C��}(��Pz#n ���0\C%@.ؓ����]�T:-�X��555�+>��V��b��y�54���.\�$���9}�̗K&�����ngoo������ �q��՚���хy��:FirK���J�>�W�p/9��?<�&�7���򨷞gr88��ɞ��Fh���Ck߽��?X�Tk��
1b�9S�l�����L�;��!Db��u\g0B����@���`v��~��N�2V�PJV&�&���'Ґ�3��j�Zv���U(��G��CT�o�K|����t�f��O�S���;�L�B�D�g��Ϙ�|�@�@
�|h�^5<��@��t�����ᬀ<�^dǏ���.ppp���=��W���ˮ���fJ1����0Z�Q$l�b��;o�'=���!F#@B�kS�*j���lh��T�=[���L�f,蘢��c�PF��HL߱�Ȕ]\�����ǲi����/��Hz���/[sǚ믳����c:{�ҿa��?�j����S~���䀍�9��)�c$��M,̍ F;�Q����H�ç�J~,&ʯ��%��A�V+W����e��)|�O��=�߇�5ى��k3I�6���^�c��uVjC�
s�#$�ň~0�`1��cu<Ĥ��Խ
��\�'S��)g�Gi�4�!1�Q����FRC$����A/��{Ŋ��=z�U�Q��O�j�������_�9}vt|q���C���Μ�9��Ç�}=sC�U�Ǖ]���+��	�$glFϲW�ut�2�f�^��~<�w����z������O�sp|��9�fH������W��=�J!N6�v�<h-�I��@�S�-A�@/��7�:g�2%�f��Lɋ�f�TU�'T$���ר�fO�,p�l�g?� ��z���e��8[����r��ɓ'Q�8r�
���	�Z����"-7����Oݭ2�]t���Y����{�ر����e!#z�o"�Z?��J���%�S��Iœ�흟��OeJ˝V��\�텅�����3�d��7�����ۙ��z�keP��Gധ�
 �S�g��:�c��֝;6�bĜ`DO=����s��W�-zqUR&�$���r�32r���iX�^�8�=�֪d�F�6�	��=�9u
����s�6\0m6�O����`����nn�̙��G�K��~SIՁ�6o~f��wpg�s�7�|S��ƍCAڳ��������1}�D��~{2���[��=�<FW�+A A)̣`��+�����m3gΌ����S�d���m��oݐ�HV����=V���5�ad��q`�ŋ�Q�I�L*&�#"tLz#F�D���O�Q��S��{P�{ME���|� f�I1I�[���@��g Ɨ�`���x�g����X ��~�^pL�K�u�-p�g�tga$��u���Ꞓ�|�p�u<�{���t/Ť�T=)u��G�ᐍq<y�"T��</�h4�-w��=)w�����r������pEEE888���9�6���	�5.��鍶pTN���~d8���1q�b����ڷ�HKg��@�w�w^�Rs��u����*ȣU>A�L���*�u�O��O�E��C��:��}������g�Ñ��1���A�tv!��@���<����A��Z���;��:���-�vl�z�C�c��hgMMM�b\,g$/�)mvr�]�!w9s�E�y�n�#U���1*u�yL�*�|�^��uG���<����p���ܐjwYw���s��"kB��-S�z�� "zq� wȏr�c�����ĈVԨ�*��|#|�G�9r�=��'�i��s*آ�-#����Ħ``xO��� ���O>��CQ������Ѐ��t67ëW�{?�!tY.`h�������sĤ%t�X��(�qV���lx������L"x"d�g*?U�'��E�+�w�IN�E1姐��#���Ϗʽ��ǈ^b��PPPp������98�8�s|.H�6͇w�p��M��R��]
GR�eL�GĘ���q��SV֝���h�,l��h�XfS��\U/�"��*��/I[���V�Ĭc�@�q�84j-S�z#AX��3��p�U���~owT�\,l(r����uj̚;��hRR�׍�]����p]G����sU���А���7���GG3�������N
R�T�G��*U��<{��0����S����������5����H�]t�_rp�yp���\��>��Û
U�<Siq1�ɌHRD1h�/!��,�ۏ�{��lVL@I^.j�C�E���nA �{�ML�",P0kHHt� �>k=��1��0,:-t���c�M�I�=�d(��9:�,��K�� ��Ӎؐ����1��1�T����N�����͋�㬁��cӛ�[f0BV9��NF�vtu��}�Z�}���|~y_^ٛ��=�V72 �������9Ԗa�m�� �p[qe�888�,8�s�U�����͗�'�<M`��)��J@T�"��h�������i0�M@�o�?����\.HYd��@�É��~8Xp�6j��c|�m��-⌌��I��$t0�{�1v�9�����,T,(�aJ�X<����R[3�r�*-��
�$���Hǜ�b�[�Q^���<l9��������3���)^�v�}�v۩�S+X��Rᅅ�2a+�x"���z�T��J�+&:J[���?zBc�'�s�++�~��sp���d��ױ?�V�ޖ-��#
C%����O��/H���*I����d
�����z����"�����%����N����q/�T�F�jW�c�}�)<2�a�{�~�6�A��a˺���u0�i+ S�N��x�X��F|��������a�9އ
k��ڋ���s�?�������_��W���I�wvv�[1f�F�CCC#=�"{%�����B�)�
:�#
_1��¯�=���qp�p�����2=�{�tu�K��-�1F����0.f�:�Ic���n1�֞~�ldk�����(!�����(�Gv�X�XX�Rn�a�S�4�\5<�VE���������qX�z��O��&e���`a�O�$[V=t���ցw��+�b��DK��9c��W��ѧ� MMM3���'{\ڟ��xrϣ��˙&��w�(y�hW<�9��+����s�)(`_��h6�*((����'{����ߟ��]-x}:���9�ŊPԏթ��g�Z��`1�^c�Q��MG~A��Z���1A`�^��5-�ș6	j� +��	�!Ђn���dG=2ۡ����\�p!|�	����0��XbOc����AE��"��q���p����؄���Q�s�Wn�$p������>˃>��������SjTYOi�`8�h�
���ߓR��(���l9��j��۟K�3§�����N����/��=�������/`�]��Թ:D��{ �Mph�SU�4�Fk4˕�RRD��
wk�ͩ��*��=6j�B�y��a��) =��t3ә:�B4�&��x��(W��F*���*	�5����?����*
F��I���73�0R[�����$.%`�X��P����3�.��c��������z{{5���)�Ge�&�N��������◯J���4���z�v�鴺Ccǖ�L�_'{���{�N:���/�q�[b�x%�dp�Qä�c�)i��OI{bQ��Jsm0&t�GDH��*=��_oЋbv]9S�C�����5wCJ ϙ7{�S��Qv��d���5uZ�ю]�����D�]kW1BOƐgʂ��65iEĠ<(�`���f�A�"���oN�;�g��պ�k�.bd^��\y��Fؒ1�R��̰?3�N���{�d3�g��"{ń��ܜ�����1���+�d��g!�Y������egRS�FF�l���P4�|� kbq��GR�����cM�j!2�ՉL���b6 ��4F�1�!���x.�����/�@Ʉ	ظc+z���QT����]Vڻ:��S ��j��G��Y��5B!�d�&�� Ea��b��Ϧ6�Q��vњUo
K��V�s ��Ӛ���Yi_�]q���ϗ�=�u(���S��Iy?e�ٻ�Կ�)�|[�J�J��f::mUIY�>������ɞ�������
5�����S�M�g�Y0"�Ң������ς���>L�6BC+����� S�aP����:�M�A�&z�C����6U�����@o7�i.L�DiE)�l�/tf�矇.���>c��K$���fo��X@ARJ�j���}.�I7d��]��[���K�8���H�x��~o`��l�z�>F�є-�J��������@�A�����Pz"h@������Ke�=����j�muu�v 9�%�ᴾJ�9��ϟ�	��
N������~�k	i�iL��#�fG�٠ż���6�V�q̘��OWcǞ���~���ǔ�VH��!���t,8 %����8��j���?r�j45��qX�T�E��ݡnL�1;�n���q�� �mv��503bW3��	*��г�"�f�6k¯�\��/?�U�9����c� Lu}}}�wL�(}���%�ߩ�^v�Y!�R�r�}B��#P�eZZ�b_I�Sʞ<(�O���){��<��jݙ���_'{�O�))����䂎�ǖ�B!!k�L_}1�ڴf��%�^���VXCa<���`��9��و��|x:{��ur`�j�`՛`�Q�w<	��d�������|=x��8��g+<:������]�]��0��`6��>$�	L�(�,�a�U���� �eD@%�C&���ǝ��:::�n�g��Аa`` �!�<��l5�)|�����<�Q�&���*|]<�G�~�.bo �2�^I��[���ugd�6����s��=ǧ�޸%�z��[��d~qI!�LmG|�șR�.1���}͵(�[p��wBm1"��"���I؍&�),���qh�@��c&�h,��M�̠��#;�ZSu��>{z�A���L!���Ƃ��<���(�O��&-
�f��F사��	y��D�B]�3�7���ԋ�87����
��en�[=88(1畔��U���N�����^�W>R���SE}�<g�4g�YO��Ba�N���4g���9F�Y�/�ϻM�f�u��4�K��LXz�L��[��>fO�D81Ȉ݀�˖`�@[W����B K~�L��ۻy���A\s�W�Hwb��c�H�E_,����@��G���ŁHЋ>������^FN����q";/G�b��	��Z�xL�ۍIhi���5[��N����6N��4���g����������{'%N3�+**�Q��5�������v:

�ј�GǨ
�Η�r�Mt���T�~D~�j����1%k�ϟύt88>'8�s�����	����\s_W;��ۅR�
e���l�����`u2u�`��	X�h�����@���L]k��Ű���x�&X�
��`���>F��	�%�Ȯ���Sh�:�XR���e���ԝ��F��Aw[�B�*����42D���@Cu���$@��"&J�1�0�I�������>�ܡ��.���w���1�����X�UTT�����V9R��§{��e�i�aJ�S��<a��^��'�/ʩ��VM4�{Uiia-888>78�sȐ�3��?�U���ѤE��J��(���7�<#T��ɠFg,�~��[Z:p|�Aح6\�8}�[�Va��8��=#�0[����F2͆��s�Q��Fğ}WO���l�D�TŨ� ���JMM�����S�F�Z���gU�N�e��$S�b�ݘ�j4R{8�b����۸_�9#b��?<�=�L��,q��-f���ٽY��'������zGEy
 ����R�#��ܚG�(ů�j����&L����N�r���~<��P�-%�� �� ;�P9FĞ>�>x�J�J��7�1S'�����S5�`ϧMC�g
~9N?���A��"��Bm0bWc=Ʀ��>v~ߐ3'N��7ބ��Xt�7����b�:��)� cn�T��Խ�hE�N/���%8MVH� 4:"�ӳ�R�C&���}��M����8�hii1755�a$�Ni����8�)�M�N�{�=�V顧牄��ixJ>Aq�S������u�Qppp|np�� ��2������*]���|�-��p�Ɇ�����֏[���t
ƌG~�x���W�c����+��f��QZ���v4>�lW:�����3��׽q�D���3k6��i��ݍ���x�ې�*X���12��$�E���L��XС�@�f��@�����{�&F�XF�>�Vl��̺n�Z>��ܢ��7��ԁ�-��Y��gΜ)��yX H{�{m��_&te�-�Q@�^7n�l�C�S��T��b��l�f����9��������ɞ�ΓS�qq�ZJ����� aa���=�x8�>1� [��-� N� �GN������8r���o1a�8l��#T��E�Ǎ(Si�������?"�t��\H�=�)������ً};w�\2������� �ՅH ,[�j��Qh�$��sM{����4:-��<�'�U��c_���o����q����:�)�2�ۭ����^XX(O��[���z�rP�L�#��Ey����H��ݏ���=�C��~v0�t;
����������<��k�����b$\@��^���:�H9m�}lq�9��ӊt��|���L�(��`AA7�z+�UVⵗ_1ce��+�����xo�n��]8��C��h�p555�058�nDYE%$o ��2\{�Mصn#�-=0	�bլ���h
�-Fxt�����X ����OY�_����㜁��|�ɋ����-�����|�
��~7!@&y*�#b'�V� ���i[&I�U���'�Oj~4��{���J-i5����������o'���j��Vu����,	�7^���߈��&a�r|��z�{��j���/��#G1�r*�}|mu�h����d�H��/���HӚ�n�z�U|��;�^Z�G~���b�[X���p�u�aΤ�8��c��7�=0'#쩫/cA� �������l��0�+4�~z*�X �`�d��0��%��C��kgM�U��G��bD����ƾ7JߓBW����SC�H�������P;&{���H�#!�@��>�y:GI�#�^���m�����j��N��1b[��7��ug�N��^RӘ���Op���W>x��ړ�<�����`z6�z0��%���h-z<�8q�����o` 3'O�ą�_�
�ӎM[?�Vz�z��Hǋ/��1?�n��x婧�I}�4��r<�UG�Iu52�:��p1B-��8T��'�F�D��S�Z5�L勌8�ZU|@�ٿ�꫞n����C����_{�K��x!1ͫ��͕�܉̉����<�H�+�{��)}��*_G�O磻�	�>é{zMJJ�`~~��ٳg������S0U�:��OC��9���+.���U�x��[�UT��>�f�(�b���ـ�s�c߮���-���fX&O�5˗�ԡc��_�D ��x.n�X��\�eW_	#i)�D<��-�R<���짰��(����_��~�^?j�;7�P1c:�w4c~��d5"����T�q���Z��,���̛3�ŉ�=և_��Ξ�����c$b�on����e�N)yJ�S!��Mi����'���b�^ޫ�L ���ޯWz��}Rs��O&.���	8ٟ�oښS}���6���z��� �-^��;v!O[��U�p��	\�d��!h#X�����F8���.�D��{�+�QB�m����Ow�D�>���`�"���b��&��׶����k�b����e{��i�:p�8#�/!1��؏V'7֫9���x@%�X8s/��>��͵k�3��w"tJ�+�xR�}\D"�����%Fz��:R�t�hO^)ʣ���^�[OCrT*}Ҡ����dt���'��RU���~�M����_�<{*r&NBҠ�����~���o���P6�^���]l�N���U���%�k߾��(�&uf���d���7�E$܆ۯ�e���������yyX��Zlٲ�y9�����XW_W7�L���6����r���Ia��~2�($e%(%$DTj���i옷���6p�kh�n�����ⶶ6���YY�:w:�2��+3��\|G�@_o�������qii�����ʜz�*��������+�u��^����w���y�jw���o���j��b�}r�A��O��b�PgZzZP�g��K��0������0Tx��M 㳛�on�L{!�?73[�?�P�т4�f�	[�x�'0�����Ĝo���w���^u)kj1�,l�pfWNFz~�N���ff�����C�Pn��SA��O� 1"����btˢk�	�;O�c�>}:���a�{�cѨ�L��PQ1��m��v�(�n������o���Co4�$y0�	�$/Z�a�'��ק�xD��>�H	xR��(v�)++�U�'8ٟo8y2�cϾU�,�\=S[*[��*4�؋��.l�څ���Xq	
33�t�&�qU��B}}?~�ċ����?BH
�����g�^�k��
'ƣ?�	��p�b�lJG�������t9d�w�m�w�t��@��[�����cժU�� b���FvZ����B�A�R�:�ԃx�o��D�C�> �s�}�Mlio]�ZG�u��N:�ꉔI�S��q�nw�O���L���6����"�{e�!��O�x��k옘���w�ܙ5|���N��H�<����5�;z���� m���0T݈�����U�P>�'��ഥ#&i�*3�;�Ŧ��C+d���ٓ�S�=|~/l��hh�E�`'�ҌX0k�`�!��0��D ߾�<��S��DB~X�b���19];{�,?U�9� �Ȗ�����֋|��d��e��"n3�"ѝ�gL�v_ ���-�����^�7�=�(�:,������S��R>�t�le�B�D�t}��V�]�@!{:gxܭ;/;�I�&�*|� ���#t��V��'��5;,f���BC5�j1�`������S&@ѡ��1��M�Z>�����Q�h�F=MZ��'N`FY�q��Ǟ@��c�2�����^��}�ǞaǓlש`d~��	D0&���9����t%B�A��&�p�0҈S?}�$��3�cq�j�3�pN�\�U�x������\F�3��7����a���#S����	d�C*_��F���\��'(��}z���I�^�:���/��������<���c����K��7;ML�ա L�>iR"�:�lF����(/,Ee^9�=ܭ-w�1�t������/�3����-�^ܺ�2��6���h�sN�	S߷��m8�DٲE���{��r�X�)�)*���߇��&�{�#����Xy�J�@Yz-������дw�� ,j�ܺ��j���IsF���K�^���v�=�
���_�
I�+�m����"{E�S�>��Z�f#&DF�F�/_1�F+R�#�k4��V�=XR��	�����b�-;K���%Y:�Z����OF�=�=�d6�
P�J���;��A$<���"k>��s�cby1�Z��r����E@�#f2Q1ס�i��bHC��jh����a�X���E��=����|Ҽ9h�s@v�[��+�XY&��WX�8�����dd�E`4�JH��e��X;��+_��s� 8�9����������������Փs��O�T�O
����>�B�t]zz���I����J��p�_b���l�*..����'����6.MvtNP��0����z�x��N�D_�&O�-��.9��#����''k�S1v��mMx���a4��'�Do�������NǬq����K��Y#�~�	�5����ݘ66}nDh^��͟���L�6��;�y�Mٱ�fzB	�1b��}�J,�ю��Ϥ�y�]e˗��8�-(Pܽ{wQgg�l�ۭ�=�hf=�Q�='�&�O�}"v�=�������@�7*�@@i��_O�A2)�ߎ��&�;�^�������y���'�������FZL�3-)!���p��^�ńc�>A�� Z��0�s)�O�q���B�_[�n�o��Y\y�W������MX4a".2s������WA��Ę��x�n̞:�FZv�Eq�3�#"����=�
�	���*�`�_+���#b��%�4�GQ�k�ҥ� �h�k����Ocd���<J�ɤM$�8�QQ��O)��ޙ�����4��h?|en=='�1���t����z�����!U�Y����K#�1i��`��*��bf\��������a1��]{b"
��_��р�3g�^X��<��G�`�c���k��bÌ�q�ho��(�eeX6c&6܏����1x�/c܄|���6�_�ߌ۾r,y���">¼���e���GN��ߍ�Ph�tZ�=�ظ�7=��cX��t�՟^�H�^__/+���rdff�dOi{*�#u�<&�'����'~$�I��^I�޳��t��d����SY9���>�Y '�b0��Ş��3"�i����C��j2�PF�1O,+S�#x�Z�*B���iC0�Baa9J��Ǳ��f�^����=l��́��N,[��]hb��Ѯm��8�݊L���dӦL��7�FwW��>�Is+�;6�փ2G>:��P�h���K/ƲK/�{�y
��hUzz�����Y��ma��!p|!h�oɋ�#��n���oI�ggg�*]������2�F�E��v�)�)z�k�=�{�N����ƍ��g	����q�x����>렻$-)A�A'haЛ �pGEY�1Ro�����ȵ-ٚ�e��0��uڏ�������";?�+/����ɝ; t�`�/���3/X���BŢY�~��������Q\��?X�S�w2��=�_�e
.�H<����x�-�o��߾q?tV��%��H�H�QuI�{sy�(~�8�=h��G?��<�ϛ�����Ę�SO���>G�M��j!�L�K*$>��i��T=�<Ai�S�U���	�����g��Y'�RЬ���~�����%���a�TjyQ�3"�ZlLF�a7`�M7�Tu�v�Ĥ�BDݽH�5������C�#� 
C���UR��� �N��)�J`S���?���R�3,hcJ0=���̂(Űs��2qԒs��@$���'|a�v�AҐ��h?z[7��%��èCw8�2��tWz_:::��4��m�<��6){"l"eJ�+xd�C�F�^&~���C$(d����{�5�1�cz}j�����	�W��q�����{�oz��;:���^�H�J��7E�-�A��:.���a�h9渣�s�ux���K��?�Gw$����-_�ӿ�d�Βb@-`����N?����׭��GPs�8�����sp�U��ц��&�X8��YH�����ق��?��Bxs݇�����w܇��0����Z�x����xz�S�����q�@�����%׺��܁��)���*�P�}^^��ꉼ������
��N7e/�������ze��r����G�(}o �Q�������Y'�B�-n�W��7Z&��զX6�����V3�z5Z�>�N��� �p��7�Y�|�_F�ı�)-A��=Luo��f�;����5UL���GIn{�s��p��	fI���م˦�C_� ��Z�w}Q�h3;?��ӽ�����i(�d �]�`�|�nSg'ˡe�޺�+���cǎ��m�6�����p��������˔y�=Wmܸ����񝝝��<�)�*��8�Y�~J��?�w��Q]VV���OOmw�:�Gקz��=~��2ҷ���v���㬁��?!:�z+���A��봈	h1��"�*5�� �qyXx󕀉�I�������L�Y��J�1����aӻhmk`?s�]����۲�X�c/^L��o{7�{z�%̜8	S/a�Ϗ=�B�% ���)CGM;�¨(/D�ۃ�ن�ieк%l��K��7��5X1s.^[�.R4}��S����,����6<��=�q��p4Z��N,��s����Ү�.;)uR�D�d�C�����b<J�����Z����:N�Ai�S��z�H~�b1��0qҎy��qd��N��d [ܷ���[TuM��i�*C�5[K%�gu#~uI�}�8V,����ٚ�4��	����ʟ���
�ܻ��n����]���>��4 �3Db0yp��4SyQ���tL �q���n�Q��@<�̂DX�0�G{U=Ƙ�<؁�r�/����Ħ����l�M�ok;:���7��1p�50�����?��Hz#\��������>Id�HY�T��t������8��RiO=�����{z�L�S\�"ј|�*�)@����y��Iڿ��}��)y���삓�?�z�㵗+���\3Q͚PA�D2��V�[�@�&�q��qх2ы�	�8_p�%(--ƺ^B�ѣ�dz#Al۹�p�K/X���+Ͻ����5Z̾����n�GGWz`wA�;!&$�[���Z���GQ�*��=��?g�sTFHmh؈y���3 �Ӂ�Ύ��.}vQQQ58��w�w��
����~&��ࠟ���_{�e�Y���s�͡n�R�T�J9�
��%���#6c0�IM3�z�a���E�����4o��al��	焓d�V�\JU%U������;��.z�z�V�*��Z�{�'պ���������8l���I��[%��!�!:{����!��㿱��.%�X�ϰ��0�e:���ZX���0�W�ul0�mt��r;�,��ϙ3Gj��#b?�8{֕>v�C�3��4�4���d�)�[��!+C=,����D?�P��vP:�$�h����ӕB����!��?����/P��"7���i�[ۨ���ʂA���k�]E��,�'�C�G�Je���4MM���P?��'��5���Qf`����-�3���y�Fz{i~y�*���Оg��ʊ*�KgR�������'��},K¥Ĺw�����/c�5�����Y�v�|��W��}b;��|OO�q�4�O���F�ά7K���z�����
uҩDa�*�������-��ID���E�x���ñ�R���im�-7%���ӵ��K�UK؛O�����Ѹ2���D,L%��t��R&����'�+��#���l ������*gϝ�׬XES�Az������!�ˤ�W��e�����T�fD�����a�h�b�Zn_?�n�@�	�-�ؔB��r�s�(���Ϗu���_,��@�"Q��vx�e�L����qu���W�8q�P�h��0��s�QZ��N>��[�������p��|��c��g# &�!��}z}�n����w�M��@0� ��  LQIDATsŊ��I�K���$!����_��5�CsB�������S?{QC��/��zZ��������ƀO�٧�y�����)
���G�-]��^�%�fO������ƃT����}���(�?DMQ�/HiJѵ�L5��Ɩ:��+0ClP��4��GӲ�kخHRWo?yY <�E�O%���|����ߋ��o��m8F�E�Һ={��fa�5�n	�BS�;�������ٳ�СCt��	%�p$��TU��"���������0��� �_^fGk<>�2p.^MӮ��!��p=��1R]]�}˖-��ˀ��$ ?�g���6FO7����R��"�}���x.M�,�g�4�y�z�_qJ9�Y*ğN����`L(˥���5{b�l�L6��5t�}�<l9�;z���I�h�k�+�]�ޠ��ar�24�b�Yu5��"���s4���޽���x���IM�C%?Y�,y��%�aQ4&����|��D�u�]w=���^�ԧH����]����%�Y�+X\���
����o$6T�{�G/������N��[@�H��Px��%���W���I�PI��Wv����;���Tv~6��7o�!I��˃��d�ĉ��#Goo����X����)�f�=�6���"�5��|�r�)U}�ٵ'���^~	%Gh4#�iQ����o�1�a>�^W�����_�7z������OZ�y{����m�R��G	��k�8r��}s�>
yC���;&�D�`qIE��J�!ᰔ1��`�}��h�k��Ŗ�|�O���g/�����ֶ<|�ż��oCy��o|��)%����J�1Ŏ��_��WJ���o���̙C/����_?00��v��iǚ{��n����=�RWoH���o���'��վ�h�Ɠ$�eA�~0����]6�EcN�2��i8�\(H͉$�yt��[�f�`O*O.44�)�"��y���N�J�Jes�m�:ڤ8C�_B&�FF�����������l���+�k�(�7���B��)t����T��h"M�N�����)g�u��X�S�9�'��-Y�z��Ĺ[?��w"�Z&����=�����Ͼ����M�FǎS	vH�;x���K�9��a��]�����8���򇱀P<^�eo'�2�����~�z�l��>���H4J��-�I� ��	N�嗫~������'����I�(��R�=�c����{����S�ǷR�ᤜ	���p�L����h0.�?�}~{#p�œ�yK��K')c�(X]�~п���Q�_���O��wSǩfz���<���$������ө�����oQ��O�d�����7	cv1��Ea6z(qΚ�����p�����`Q��[� �pdΣ�-j瑅�	v}��/\�P��Cԯ��5�]��wq��7Sgg����w�믿N۷oW�#C.y0�������������=�C```�Z�x����-C� \rD�'0h���{?sO��㆔a9�^9��=Yy�d�.]���}yׯ%r{	e��0)Ͽ����_�ŉ=�pL�Ϫd�DJyyx������q��}�G�CAʲ1O�����t6=��o�Rt��7�%t7$��?It�Z��f�:���O�\�\�,��>6*���?���E����y�������[�ûH��=t�6���YAv<�� �H�Ú<������_�pA���Ϡ���J���ÇU���Ŵf�jl<BK�.��Y�h۶m��oniQb?{�lu]҇�Ó�T<?.��	@�����l��ۿ����:u��S����'A.)"��e�����i?����b5�=�P2M�l���-�5}�FJ��q�ay�[5[���R�_?A�������v
%���}���X�M��s� �\�M�]�Е�t:):<Hފr
Y����W���C4��EK?{��G��Mǆz�'��),�x���A~+gR�a�p�=<���?_��C'�O��1<<<�_6�߉��!�\x�X�?~��d�<w��9և��[�ѣG�x�-�Ў;�{\�g�Q�"o�ʕ��ׯW��+����x�X.@��1#��*
�$>�27�:����MM�������_~������{/� ���JW����?zGo*v��@���RG'�3��3���9�O���"�=)#ς�!u��W��kQo����=�0A�����̤����w�ʧ��ھ�W]���e���"���)��Q*���y��r�Z������%|L��z{�r�B�v�*z�����|��`P��clL$|�|��s�_���n��"Au{��ث_��gx���_}�U��~��i·�_w�u488�߽F��XC���hT��/_��������vr:���tZ{# �:�p�wܡB��<~tݛ9c�J�;w6W����Q��Bk]���YoY֗�;z��}�_���y�m�� ����W'��vs4�ʬ5�C�UT;��Z#G���o$Wm��اJB�;��2��S�L���d&����>�y�Z�|)���>88@������,��l*�Q�yND
�ȉ��T:�B~r�}��&(���T�������0�z跏>F�/���Z���R����#M��z�B%>vR*^U���~��K�?�L�aϺ�5�e��G�_�d	�8qBy�,�*K���6�}���ݣ�{�޽��7K��a0�:0 8�^���	{h��0��?�i:r�Ha ������x�cru��B�}#����)��g��Ç��i"��p	��`�k�_����t��Y�M?xd�Y���F��v0XE�7>�D/<�,}�O�LXwO籘o(�p��Zy:N������<B��ϥ��7��u��H�Pr�|6�T?�&���,��	U����}i~�c��x=��/��S2�!��K.��S�>I��!�m��OM���J+��/~�v�x�̝�o���z��}�������,�[X�}w���<x�$��²�J�g͚��>^�T� ���1������** 1ǵ����k׮-v�;y���QPYQ��0n�m+=��������EK������2�.Ke�Q1ĆH�w��]����h��U���Cwgۺ�۷����9+K��sӷ-����c�G���iŵ����h��k)P]�����cI���8/Go���l�J�D��}�I��RE��E���p��#3ȞJ/,�R*���Z���x��$KYexY�3�]l8B�g����)�w�m���O�}��x�q���6����K�ϛo�wy���ܹ�$\4��F~����v%�yd�#�%oȜ��#	k�0ZZZ���HЄ1��v$�uu�(��x��?���:���# ��~��G� iɁ���'T���?�9��z?B�3g�P�#�d�f��{aٲe�$�%A�~��3�]����?�ϝZo~��[��_A�h�2����fh��E���9������R������%"�f����Q,����A���4��V�C�c~��7i�S�Ӓe�PiY%�.x�9�����(o�?�d�D��z�d�q�$����G|�{��t���^:�{/mٴ�FF#T?s.ݺ�vji>E#�H��L�}ߟ~�uc�J)�����D���\�����;���3�D>[D�͛���Pbo	uC��08q���UЖ-[�10 `4�S�z��C�V@?��̝;Wu惘#�F"��c���6��DO�J�{��w��+W]�B�����7!��	F_w����ӱn�*��Q�$�%c�A���z�Imn�����~x>��e�^8���R"t�M�/kR�J�N�T�=��E�ۥ��t7:��G�В�+���=�ӭʪ��4���G��q��=�L2A��M���h�|�<�#I���+tӲet��~Z�z5?v�V-[K�dJ5��s�Dls��V��R�K��L���i;�v��%p�⏵y���:=�z��F�^{�J����?�q�M���U���S��'q�������V����7�xC8��=���qH��Ӄ~�n��f�������^on������9���`,Y�������HOOo�ʕ��O�9E�Σtx���Mᦓ����i
%(�P��;�w�E�~|+���/����������C������ZO��A��%E	�UX�������L��.
JiZ�ry=��G�]�W�o�$��8%�#��!��>��G�{����
yN���|����Y�Rqz�׏���5u���/�{�/����-�Ҁ���g�b�~*^���X�;��=xƩB�q��D����[��&7�L�>����q���U%�!L
U��e˖з�����?���jI���F%��\��\|̹���u��믿^=��0�n�q|�X�7�����xꩧ�ŋ�	��Ȃ \4"������}�7_���g;ܞ��]0�q�^�cx���Inv�=C#TOn4B%>��:�����7J��,��x��;L��>��w��6����/Q]i�DGh(���=�l��L���p�������jP����;���#JFh�L3�ycUEbԴ�-jm�G���Jk/����g�~�Zj��7䣷�t���#$\�s�d�z�'W��P��Y���;���ec?�k}d��sSS�||�Z���mW�v|��C)���D��>�|��� A������ܹ�zzz�}����jG�����Z�:�=��c�ә�����?�8	�pш�O0
^����3�-�H���g����_?����P��,9=�]FU�C�l�B�rJf�T�-��H���ұ�MK�Y�S�����4�Y:wp?EK\��?�3j�YO�L���{�q�A��R�C���əs�af��uQ6ɟ1�6�?��m��S��#���R�R���3��~D3gэk���#;<kN�O6}����$\<(�������k�k7�q���|��k�k캄!x$�A��Y�s��"FX��W��#����nR��{��GR���GT �A���X:@�=�G���K�Z?Dp>�e``�.�J�?������� ����b��Q~����ytǶG~���=?���/�9�n�tF�q5���X�D)��Bn'e-���)H{�.���hw�~�M_��FӖ.�]����A��뽪�.O_?O��i'�9�<j6=E�t��Q���32�������g-a����:�K�\�нo��D�H���~�E���؀�C�!���!�h��� ֺf޾nm�����A*,Pr#�r��qm�5���;�nܸQ�cy K������c�y`ƌz�l����.`�����u{�$����I�� \"���M���;5uUg�O������y�����%�J��94J�\�����)��L�)Gy%���ᗲ!O$���-�6�/��G�ɯ|�zs�7L��믣�e��ޡ�T֮����s7_7Of4J��NӮǞ�3��2~<:>/���=<d��a�L��lx�3������)	���썯a!vA�5���$<�-�� �{��#�nѢE��F;]��57�*ϼ��L	9�4���Ã�~=�߫ɉ��D��#�����C�-u)@8���w�0X<OY<��F2 G.�I@!���?��._���)/m{�ɯ�F�+��ndh��磜�I�In�aMb���N�{��=���E�a��#Z���/�N�ۚ���OK�l�T.I������g/�4�d��N%�D�H�η\��om�� ����I{�/E�	ʲ�����}���7� ?ޗd����n�S1�^��^!���!�]��!����GX⌵u��#���������>O����j��{�z� "�`����ذ����m�W�>DQ\y �իW�e<�G� D!��-h� 	��p���O"
���/�=������x[��}m����,WI%f*<L�T^M�˲6����<{�喛v?�"UMo�ֶnJ�wR&ߙ9r�X��9�N59/�tP���4����Ҍ�s����F���}���=�t,���(i�mhd�������Ei�r	ao���q�WϚ�Cf�i��IF'�A�!����e�G�<��^�5vlX�G�[��!�f��q!���x�׎�yܫ��[�K�͛7�ny��_5gb���{�nu�ҥKURD_��{��:	- A�(D�')�����?�?�'������xd�;_���ͫ����ϳp;rgs*�ޠ,=~��ĩ��9��G{{��⨳�<5��ea@�d$N�@������^~,��ڰr�8r�2�M�i���P8��t�"�>2rd����?!�2���,��zx��c?^!�z6�ܱ�������� C��ec��n��Wd��ٳG�GT ������#!%ur>�	<^�����ڸ@� 	z0& ��40�:B��� ?K� \"���BRS7�n����~���_��T���ps�@"QVϘ�L��\��.'�Y�=�
��w�������t��>��_&�/&?��S��0k�Q��s���M�L�Z�3�Q=��r)��D���p����L�����ϐpi�&�9sf3�w=�
�Z��a�w��:�Iy}=nǡ�^Q@����,z���X�����Bo�ٷ���<��o�Y	<��`�H؃��8ϴp�|-���q:��}r�x���W�*}���� �?���ZX��v�x���Oٶ�s���ٜ�v�MJb��;@�X�L�)A?u�Q]����6ү���h�֭���O���s���E��ˣtæ̈́HAogY�~�u��	r���_7MV�����m_���|I:�]Z�,���o��B@�ސP��ا������b��;2�!Ķ?U	9r/�4�s�a ��!�il��Y�z��� ��!� ��q�7������m}���u{��1#A.�}�!=��e���_�u��W̌�n6ñiN��0�)#��7��Xx��,'��hv��O�������ђ�7���*zy�:�����VѪ9�h��Ô���@	��)��|�R�}�k���ύ�����K�(
�ϲ���6��}x�j�J�!���3��c ��GZ�b�s��䧔���wc��x�b���s��/��'�T׃� �F ׁ`# �	��&J� �ol� "���B��,�����l�A�hD�?`B�a޶�w�9iz�g��O75����(�+����4J,7��}�;:B�(�I���㴯m�zM��>�Ij駇��_(�NR0������!��hǌ\2��2�Gl���}�ÿ#����А`��Q�JY0?ς���b���Шk���d��T���-�k.\��]��}�X /���ux��q��<��5���C�`Ŋ����Vw�h�wp��#��(�9j�Ø(�*	r�\�T �k#A.	"�`��sG����z��s�������}g�r-/'���Ȼ{U?�
���dR�2)�pS6��$e����r/�M��!*���XW/����z϶������Lrp��OR{��ŽL��F:;;�^>
=�B�����	�ZO��	sh�OB�p;��!����	/�K� �ا[�8p@	��q-\az܇������Z�Jy���X ��������2*	��a6Qe����!b��X�a�����?���x�®׿���|���{����@I&a�����2�I^G��"ar]�_��]z��)�~�}�֭t����������ٟ�UVW��3j_�������M�Q}aA�g��u__�A�f�y5�"!��B�N��C�ui�}x���Q��o�>\C��!�ړ0 p쐑�ux���l�� D�^q<�A�!�}\�/���YY����p!�D�K����0/��/�<�h��]����ᓻ��}3��kj�|�ᘙ�')ef)���P.M����7��J?�գ,��p�����t�L3��f������}�1Zu��6��8&Y�/��v�3�9�Cxa ��j�!���Gh"�� ���G�g��ޡ�u$�a��"��=B�h�c�z,	�hx�����V�����O��ב�}�� �����hw��gI�K������/�_~��߹u{���w>���k2��~�;�_�STZWC;������J��=���m�~�5�=0�8k�M�I���Ų��w.D]���g�b�"��@��G�>�w�̙�y���ݣ���#�8C�u=�E���k#j�n�:uMx���z�
�#D�\�Ë���t�觼n�!~�$�%C�^�71�n�D���m�.�q�����~����{�\ޙ���7�[i�U����(�?�&�T5w���}�FC�0	W��]�о9*��.�U���Y�A��k���n��b�'�x�[��M��s�*!>t�(������C���wTI�p�ѣG�<����: ��� q�3��П���9á��n6P�H�K�����J���y����[o�\h�tx��{;[�/�ҝwz��Gs׬�)�uQ�U�Gé)��v�'?�:���H�b�,�Z����S�F���^���Go^z6�V�;���u�ػ��m{Z��ܮ��\%�WT�� �h�������Uɞ���}���&;�؇�1v`����y��s���~�ZJ��"b/��E��{������?��k/���S�����s'�Py٠�K����ްn��9s���
¢��=�}�u�Y���W��6S����ִY��w��N���S!z��}�'�_R�j�j�뮻TI����_%��<B��VeU�=sNs��f�"��A'�[�s�f:����n�c�k� \bD��_����~7�Ҳ�O���3���_��K�jk�(ga�2�l���w_z�soK6����500���.`���^=DT7�ѥxz��C`����j��b�0?j�\��P#555QKk�j��5�x�L��O�"�N*�V��ݦ7U,��}a�����1 ���<n�{%%%R�)�{�߅�А�뿊��T?��/ozs�[�tww�͙7������_�B��p�`�=���X��������#�u:�� |x�h���;��{x�lD�>?�x㍴a�Fu�?�񏩲��jjj��Su���a$��Numt��Y� F��l��?�����t:w��(�{��M!���"�ćܶ-=����TtΦu}�}e��b����R~�*̂W�3����";f����uw�C�]OQ���~�ajb��3���o�a�:q����,%wXǇ�q�{���08`T��~;��ϐ�L�']��2 b/\4��z]$\5X`�`Ne��Mtt��;o���#�?�^��X��1ɕ�>������*�qq�>�yjj:��%������$=� QG;^����q�`x�ؐ�k#1�D��{���JKK%�/�{A��`�~ppp)n@��k��C�uB�ڛ���c��ǆV���¨YU�O%��#D�� �CV���a,���,]�T]Kx\���s�v�<R��[?�=!�y�py��	j5�x7<g&�z��02�-h�i���1��"�����%�z.�|�1�^Oj�U�?�)�B���&������q �A������)��A��?:M� \D�a�"j�d�_��i�[�@C���m ���;�!daGb�q;Sj�]'�A��v�C���z�Y����t8�CS���6 "���a�4�x�^)��˄�� Lhz�������"���@`�v���V=UNu���Ľ��!ji9�" ��ܲ�j�_��9.*/�P"��.�3�Q0 p�������1�{br�a���Tr0�H�e:].���}��qo���	�pY��	��`~&k�r�N��!s�,�t����KɄ����;�0��!{�ӣ�At ת��V%v:�����B��Q��G ���0:p~�K�S;}n�_TVU����t$m��V�����^/�{A�� ���ӳ��w1����b�����v[\���>������fW��{�;�Yw�r$桕.�z�ǆ{ٽ��O�Æcp}�_�٢�L���)���7A�������mY�jTȱ�b�^�/�đ����z�3�u/z��������H�{x�:R�kB��Gb�n��t�
ײ�p=8F�æ��ƨ�c������� LPXЧ����֯�m�P���7���W�����(hnnV��;�����ΞGx%yH΃���|y$���CotW<����1����3;H����� LPXL�R��,�
�:�!�@����:޷]n%u���{u,!=-�ډz
��S}����Z����tZ���E��!܏���uo|�w��s<�M�� W{A��tvv�X�7:�r��!ϫ��]ŵ{-��$9���dZ��,��F8�i0n��0��'���g��TQQC��J�ޏ�8�."��fЧ����TR������{�֏nhh�� W{A����>����,�N��'��w��x]v���
����qlGGG1��-�流�*Va�s��v�UT�qz{rB�������"	c��n_��?ǯ;�5I� \D�a��Bj.���YM�s8T(^7�A��Wg���d�ut1&���vd�,�Q�D�1��\���� ��8�QQɷ q=4�щ���Q��p0� �u�p���	F���{%o�c�q �{|��H����a�̠����:��r��WT��SL܃�#_y��|����i{ ��O�ؿU^^.n�*"b/��X,v�['���GV�b�v{U�b�K��}#��H��Q |�Y�0�i��u�]_QY��C��E{\�0pǲs��"�;��|60����Rr'W{A�`�����u>����HC�!޺�]�����=ްN�{��u|x�8������(e�Y���B��%�`Py&��yC?�v�D �[}>'�b��#A�*"��0�`q������o��s6���cG��å<z��F'�AرQޤ�����cϜ(�LQ*�Nz0ܔHإ{0jkk�����A�=Nu=����!69;1^=���@�O>��i���J]]� 	�pU��	�����"��A�\{�hd���A%ԺE�N��z=� ĝ���(��aNII)�>9U5U������H�f3��g�i؆�aŵ~P�M�!99�������'W{A�  ���w%�������=D�v��+z� �`C�^M�Kf�w��7X�G3=��H8��%�ej�M(T��^���������cug>d�Ó�A��	��@(��>��5� W{A� ����X\o�!��^M�c��������V'���G�$Sq����������S�<��z4.&��k��bY�}tb�n�S����`P��a b/ T������R	��=��G"�����M*�F�B�ʇW��w0T-�i)#A�a1��ReE5UUU�~�0�P�8 �D�ޣ������a�¯H�K� W{A�8���r��ZP!��XB��c�;�l&�^��y������v�/�#�abBh��q��w��U��y}o��c���·����(?���q��� L ��p��z�-�b�Fs����bR�m�b�^ͧ���c�٣��ԩS��G4 ����*����*��<�ao��#�o�Y��Hp9\
�(�f<���!��{6FI�q��� L X@XhW��촽m�
�#$�uxL��b���T���{[[�j����t�Q��g��zH��J�g��{;�O�����&>8�}�ٔ��5{~���r��#A�"��0�A>���Y,���c��r��l�=G�����u��9�^},W��N���?8���!�H����d9��N̳,�݋_'��������_�I�q��� �s����X�ob�-�_��Ղ���lѵ��L�������"">{��x�>*++UF@6�&#��C�d�Ϩ����@C��ɥǊ}������ml4�I�q��� �s�^��L&3�E��]��Ycv=�������z0N��:��S:��x,B�m�)�*�������u�iUS_W[C5���{�˳��?ٌ����Q����(�I�5��% ~�c�?��q�rI�q��� �c�)ohhh=��B䵨#��n�k�љ�Z�1��^{������ȠGV>J���qhy[^QF���ʻ�d;��l����fLr�P�,���|������H�q��� �cb�X9��gO٣��XZ$ۡ�^���	x���Y���ǱX��{;d�S�N�Cb��� ��\�^'��8]�χ��������1a\!b/�4�aQ�ϯ� +Og�c��yY��C��N��~x�z~��'��ɓE#�N�S�g�R ��jjjT�=�~���^���(��0�B�;���]��8"�la�!b/�'��Rަ�e��C������t�; ��A 1�#d�u�3g�(�^>�������A%�(������.a���=y�� �������lI޵�����Aw���8�������.e���Zx�r���uz^-����D����-Z��x�|�rjiiQF�C�B󕕕*���)�����ņ=�_{�|,z����$¸C�^�),��,�+��Ch�f�Mt�
4�ƀ���+<���{O��z���ު�=|��jx�zs8mo��8�\��'��w�C���>���g��ɝg��	�0.�����l6[��z�:��l�=�_0�W�=<����b��Qc��#�(O� ��^�;���uFq��^�G2 �^�>��������`Pz��8E�^�!gΜq;��U,�!��T:�7D�����:1O;��}}}�z�`�^�8=����1���5�X����(���Z8��'�!>� ��� �SD�aRWWW�7455�8�����׫�=q���^=���zz����t��Y�F�� �9���@�Qc��zH������z�G$ a~=�~L�>���s�K� �_D�a����###�ǎ�kllD����3��+��?�ʠ��}]R�0=>#��#YO���I~s|���p h��Q�٬�k��A?���׍����ii�޾`0�I� �[D�a��������X��^�&ؑ�>��B�;;;��>w�|%�o���=��z����{x�ix�ا�`�@7��_�||�F/8�!�n �{Ag�jkk��5aF��n��~�]��C�!�t������Z��~��� �(��q�JJ�Ƅ��O�|}�q��?����u/|~�<�s��; �la|#b/���<�lxxx1����{<��y/<qx�}x�x���:#a}9�@��N�J[�lQ��3�<��}ÆT]U���c�;�~�b��y���Y��\	6&�����$¸F�^�^��ױ`��I�F^g��>�C|�L��D��q�y�_��uO��K�����O.\�;vЂ��+Qk����|t�>�}=L���o�d �D�a1222��z���k쑶ɤ=7�9�� ���� �Ç�s𾣣���c������@�㣃����y��U-�Hȳg�ۆ����p�H$�k���\�|�1a�#b/�h4���>%�G�>J�p�Lv�=n��y�L�`0D����y��z>�;�m����Y�!�yJ�P�Sǖ�U�sϽ@˖-�o��꤇u�}���v�������<�:����� N�CEPq��(�#���YRR�E� �{D�a�������"Z�˲��s�D8;|�vy�w����#ń:�<<qx�H΃7�s���s�x�����w�}Wy��Saz��-��:}al�:���_X8���F:�0!��q ��ΌFc[���H$�0���Z=k�v��ϝ;�\.���X��j�ew�d�b�hqp���\��o�]�t	���<��n��Şɲп�F�Q������� ��,��~�<��H76q�z5D޷^��8�:�l�.&ёQ����p�ڽ���=o�ޣc��.�-ίg",�;�u�A����8�Ž�t](T�pc^7�v=�� �0�I����V�s�D��L��lB�H�C�u�:l��཮�Gh����~�V��4��W/{A�7��u�:]'��!�:�N{�y5D�~�DF�X�0�T;��C�a \@�!��h���U�s�a|��1��yݰ�_3|�}|}I��	��� �ؓ_�b[;<<h���cd!�z�-^��L�A�e��M�h�� ���v��\���q9���|�kc�^7����xD ��t�0~N7�	��ﬨ��� {A�������y��ի1����,N��{1ĺ��V%�%�v�^=��c��5x{�v�P� �8"�A��붍����!} ��?G3o1�A�0���U&��⻄�Z���]C��Y��Nw:v����N���#��M.���������ʋci3���ܚ)S��r�k��0"����Լ_fGF�����]l�!A&"��paAu���m��=�/��ա<z�C�!�zP�st��~;
`w�۷�Zs��mn�V�X�j�, p.2�a,�v@�ҫ�=���r;D�u����A���	��� \Eb��J��6���c���wo{�Z��n̝��iӦ)qF Y�k֬���V�d�<g���맫�?y�*��|>����>�<�]-�T���*�RCv`4 ��&�%���?�n��%A&"��p�������E��Z�=}���d����a��{�ֱi�%s�� ��ɓM���E�72��Ѳ�K��矷�,t�˫k�q�0"�< {\��ʇ,|�����" 96N�w�$C�^��L&��aY�Xojj��m�cO\7�A�B��t:C讇jwx��������l(��ʕ���/ӌ�j��o�U�s��lA��c=_w�Ch��{ C	|��?�F���0	�0�����iM*��1���F�P]r��g�u�c>��X�Z=������@7�$��^`���o��✥u�6��z���ud�WWW+Ͼ ����'"x�=��4y$�!9O���D�^�,��i�e����Z���,�x]J�Q.��� ��ɛ&�dhxh�֮Y��ollT��z�)�3g����;�A̵7�ͥ)����m��5.��u�N��/�r9�c�CB��0A��� �뻻�o`����j�ZG�<o����ti�;���Q߀{��ݫ��o���1c�>�D�����R���h@x^g���#j���羮PY�vU� ��d LXD��*���_âzC&���n�h�$��oϡO�أ��ݠ�-�n�ۥ�����y)�����t9%�H�[0�M����!���~6�iw��=<x�.�V!~�6$�mx�)����@8�b/��a#b/W��,�sA��'Nۨ�91�5k�����ىv�b����h\��͟?��ꦲ�ۣm�l���B��y ⸆�a�A4 Q]ۯ��@5��eS.�k_ h#A&,"��p�a��n�`x��Y	-z�g5�(���nw,��l�2�t�|�w(���4�Q�-�v�
קRqU����ӧOS��7ذL��8�����=�ǽ��}�>�M~�� {A��$��:�UH̃Ȟ<y�r�p���X����SCCC��=j�u�\|F9��l��^U��sb�(�㠖�sj��`$@�u�<B�^��fΜ�"v}�Ul�[H��9-g#�?*!|A�؈���y�px)��,�F,��Ǐ��uʫ/��E���1?88`���d��#���R�$���V_���f���s��)�>D`L؝��b��ԩSՆϸ�}���a������$F�^� �A�����[{�F��j��/�W���y��Nvvy�YY��;=��zx�؏D�\"N4P蚧�X�uh���P��Dt. S����������^&>"��pa��eA]���^ho�h<ƞ�=V6
*oay�
����(�C^=��,�r$�l&���UWU��=��N��C��`ƀ��g2���+���!|���i�0��3Hm� LD��
��<�i��ʶ�Z;��!�g�V��t(]��W�W)aƆP�^w_�d�j���t<$��[��S�����[�Y�À�����z�M��r��d��G����0	��+��GGGo��2x�U��w��:s�h2�V�����.%�n��c*a�?�%�h�e�������pR�P�уm �I��{��z�j�5o:�^q_�L�9��l�L�?�L��I��� \!�+�嗕,��"��;x�g=DY'���y�������I��y�:_L�õ���]]]4�az1L�����z%�?>�þ^N���Y���:���I�	��� \XD�H$r-*z���t^{�J��cg��9� C��l{��Z[g6�O�U{���f�!�Z������S�E�i����{-����a�`���A�����|oe��]��e�F�@���Y�_��E8^���8��^�������r ����������PZ���;=��وhv��>E� L
D��
�L&kX`��Z:�����-��u��!�(�+//Ueue�J%�V��
Ǣ*�/��R4�8o%�J������P@��2��M9g�m�R.˱�]����0�����D"���v�i����;�0cB�d<�zl�oo��T=���S�p��t��*Ͼ��\gΜQ��z��3�3錪�G_-Xv���V�׵��ޟ A&"��p�񰠮#���C� B���v����c�M0�W3�9JgϞU ̝�9s��ҽ!7�GF��vRww���Ӈ���z-�0ЬG������?�B�d'A&"��p�aq-c/�Z~�1���N�C=��N��'n)O^��C�[ZZ��W_c�=E��Si�����_��������ww�T�{3g�R������È�>}z�F?�ϑ�{x�l^?O�wte]�$¤B�^.3,�؋F�1v�p:L�OgǧSy
���D�T*C�HD��Me�4��#�᡾�Aj�-:x��֬YC[��H［�%!r��d"a����d�h �Mu�@.]x6t�ͩ�r8��nk;y��� L6D��2��gtttK&�)����� ��u�z�_o������6mM��I}�t���:::�y%�R��t����c�
��J�`M__{�����d�*����5����I|�5��!A&"��pa�ga�������@����y�=�u��I}��t�=�г�>KO>��Z{�'�PS�][_V�-����s��0vN=�m�A�ϖbc����"A&"��p�`Awna!]����s�{�n���ܘy������^J��t���]wݥ��}����=��U[[�"@'�\�R��z��nΣZ���q_�������d���D�^.~�e,�AݩN{�ڻ�r �v(�Th�q4z̭�9o�a@`-����׬R�q���U8���(1_�p�:fddXDV1�?v��;��~+	�0)���D,��⼊��	�Z���7=Rv�Z����C�!̨�8	{���j�Gƾ.�[�j�ʺ�>t�ӹX�]�q��e������Ʉ;A�����e �tXt�V?���Db���C����p>�u�XK�,�DGO��=��;�/��X�M�q�긇kh# Ƃ�絽x���	N~�^p�[�Z�d� L^D�����d2�Y@���NϠ/���)�N�^�^��Ko{�o\���0���BN ������GF?^qm��Y�o������'A&-"��pE�x���3�������y���|���>�Θw�쑴�t�!�,�(���&��L��.Ky��j�-r�k��v���?�n>}�A�����e���$9<<����8��W@���)��̏-�{?��+���[�������cjǾם�������Cp�_��4	�0i���C���Yh������5�����aD=]~���c��$����yfq��h�=v{�n����SA��u�v/|�8���[e�^&7"��p(��)l�����x<�Y����nĨ[����Bnh~�p�^�מ����1��t���s������5���Ǌ}���a�į��I��� \f���GX������l�������
d'D����x�B�<���!#?�B/��z;�/�>���U�>Gw��՟�{� A&="��p(x���؞J$���j������\.3�E��}���ѿ�x���C�}(T��{$��>��� ۡO�I�4����C� LzD��
ShIۊ����h45�����Tj	{��,�{ �UX�7� �N�����&9@��떸��m�Z�9���^RcmA����U��;�/GX�["��,�Y�o��+X���|�^�Gy�o���*�����Wo_����x��&$� �{A��Y����,��K&��D�l6s&���[y>o8Y���g�9�^?V���')���(��#�oYv��4e��$�{A'����}�X����_���U,��x�2�y������=w][�f��xSzS��w�Æ�0	���@�^�),�ht�Ƣ�944���6�N/f߄>��,ޡ�u�@���d>�hgL��q���!A>���8�EYw��G	�i~}edd���/g!���E�5��PƧ������+�/���'�n����"��0�($�!�mn����X,6��o`��Z�����Yd7��H�B�>�����7ī�"��0A)��c�� ���h4�{��xC��[��Sx� ���og����v� (D�aP�����"��_�L&k����G�>����q��"A>P���$���bc�o��b/���{�=�@`�A��!b/�~t��,l� |@�A�I��� � LrD�Aa�#b/� �{AA���� �$G�^A&9"�� �0��A�I��� � LrD�Aa�#b/� �{AA���� �$G�^A&9"�� �0��A�I��� � LrD�Aa��� :ⲍe�m�    IEND�B`�PK
     �8�Z9?B��  �  /   images/d18021d8-4522-4af4-a3c6-358ee97fa8ad.png�PNG

   IHDR   d   a    /�   	pHYs  �  ��+  �IDATx��}xT���;��$�I�!�@M:� �4�E?�>D�+("
*
"��HS)�JH�$!j�I�dz���}���|?3��}�<g�L��9��k�w����� ^��x�ex@���!^��x�ex@���!^��U���v��dRR��H�q�Lzt였7��Wo� )1�~���;�={�l�C��B�Z�����j�\.�Q��{Z��`)�r�bώ]����������G�ʒ���/P]u���0 X�3�����|� ���E�3.&���e�kBb���sK�w�	�3�����r��m��V;��\����DF������aE玉h��r��mC�4�F�Z̗]k��i7[���'E\�
���n����.�]�����KHOO��u�!�̌=={FTD(U��٭�]V���!""g/�@��=q��e�X��Q��Z��&�Q�X���)�7���$�1�L�|���eҀ���r���iZ����>������!cG�CFF/475�`�*�� rS{�'&�$3_����b�r���SxX�*�bl�u����3e���sxj�B�8���G"��RDF�]x���~/�+�����ov}3l�ƭ���s�>�"d۶�1m�TT�Ԁ����J>���p�����/^&�a�����&FDx����i-�4M4�ٟ~}�����ԙ3݄P2(�̙����X����`�)����ܢ�z�n����5�!�}��2���d��ox<��`�~�f����:�9��UӬn�{P����
��f,����~a�K�e0݄L�5�|���q_\�����M|�]R�B�pc{[�߾���mc�O��5�!aaa8�w�A��N��f����k�=B���K�nN�Je�m��;)ݒe�*U��sV��w� ++���W�`%� ����؏>:���8w���;��47�`N����O^�O��܌Ĥyks{_�g����fs�&$X.�С�즆����J'�5ӵ�h�ȸ��N�322n�������+0�ᑔ�����j�.��!���9v��j48]Di3OI$��r�l��u?�J-��E�U�¢B�͒�����D"�TS[5���q�[o����\�
y'N@��:��,�?	�9,&<	�"��p�T�8ď��F��������"�hm[[�;^MMK��d�����m"��PKs�cu��q���_����D�?	�X��T(�@����2�<�"�h
B�l6�E��p8�X�@`-))}��,����Z�J�5*��
{�;�[[# �F*�C(���_}�5 �Jb��[6����������k�)B�B��P[V=q��@���	b������P*�%�~�[�P�~�U���ş��p�Q�c9�F?�~�}���1_Y��V��������������1<55�W/=b����'�<v�>E�H(��h6�-��� e̍7�Z��q�		���p����Ψ��o	
{��,i`�r�N����W~�ƍRL�>Ç_,��ݧKC]����*��C�n�n�� �<v�>E�D*Þ=���{��[,���Ga�j�I�[z�ꕼ�v�Y��-�Wu��å2�R�t�V�k���Crrן�;xp?bbb@ޓp��ݥgG����ۧ1S��ݻ�WVV��z�}���h��.�ܛ����y�V��]���z�Ţ�z��͞8��gƅ��l�r���ͦ��!����:��x.$fNEH����`H"�	�6�����/(,X,�I�k�)B�N��u﯇^��#Q9�P���<G��
�E��^[���1�/ڜ��\6w��lF[��/��y��۷c��%8p��xΜ9���d22$��=b����g+UַmV[����g���FYi)M�PBD4""~��	0P��E�:u2�[��[���b����ׁ����lH$���;w�<������F_b���,6��Cb���Gm�[�O�0�m��}�N�!���j�1��1Iv����@ppJKo"H��B.eZ���N���mokAQ�_~����Aѷo_�[�>�����r:aqX����c���$@�^�f�}ᢅ�N� ��$"""@u��=��7�}��Fǎ!���??�º��g;%&�Assz�鋏6m�����*;�0֬y'`�'����,b�3����A���R��3y<rsOz�Z}��g���g�}/��2}����|U�Af�Q��##"�m6�0.����;�H��p�;�k��{�娩�b�YC8�\�Lf��Ƒ�N��syܸ񅇳��~�V� D�����kx���r���!�"����6���*G�Ѫ+�*0g�ll����$�ζ�}�m�~�n]�=�$���8m�t��	1W|����u뭋_^��k�zB���� �3zQ?0�d4�S��ħԃ�
$&$V��eb	�[>��w�ۼi3����ʒ�!;w��d0IP`v��nݺ�ࠝ:wW@�*��;�����S�zB֭� Ç�)�@�1�[�\�z����H�cgU:z���5�q�ֵ?o�����FS�#H��`��5���L���ù6|��Ϝ9�.]:Ó�jB�xb
���P�/���/--C����M�<�F�QL�s��i�m$��=dee��B>^}m91O)�h��b���b"%5ŝ����6�����/{����k	5r,���V��ǟ�������	��6��$G��H�!>_�7�јN����s�O�:��'&�B�����whi�)���r�:����JBF���
���:52*�s��¹y�&�-fp�<���V*��h��6O���PQY]]MLMǃG	���y�qy��L���!��Ξ9��$���2v�c?�q���v�Ԩ蘭D�|jkk�X������q�III����\��
��N���tz������ʪ*\(�ǐ!��~k����o�_"���U����"�����gP�<>**�s����bb $���!��rҧ�J���555�a��ȑlXL�7��V��L������kո]Y~����$>�,�3�^C����q��5�&��bcc����s�B!tZ��K@��l��]���"3e��h�_�x1�j���^��Ν{q��!l��	:u�<�f��~uHH ��g0t�f�[^^q���Bw*�~�k�<y
�	 ~�߽{�����[�.II�&���qTTT���sMD�mw�I\.7�|������9���E(--ŨQ�;\�v����A�똘ZS���^��ֳ�?�6k������}�7HL�DfI��
�"�DT�ёQ�6T�*��2���^��e�$���r��t�Č	�"�^�Gxx�o������Hk��!�QI3ƴF��hi�����7J�k��/x!�21h��l������v�(jF\l,n�A����*H��$,}������
2�4Ԥ� @J}K6���o�9����ضm�s����[�j!�6��E�MS2=D��Ǹ_�
B�eg�V�ҐaD����*��i#5��'P������
*�k��%/j���XrC�4�jn��:RN�>���bĈG�IT��B�D$$t�A Õ�u�p��)�����	� $6.y��!66f0hJ����AgD{{;"��Qt���-Ӡ�+�R�.aVFG�Ҵ	�B�2��\*���?�t��C�Kf�nss�t��`Ђ���y��7K0g�,�Ox!����T�K�-j���;w�@ ��l.���ۚ�[��Cn���W��>�H�'$�m�5��;��!�Ν�[o���{�ԩS�PSE˵QQ��h�f��GD��������իp?��Ь-5K�<<��t9��k 	hM���P���Y��`��n���m=a\�c��Dҿ'U�p7�C�/Ʀd����ҥK�I8ݕ�\h�Gf%`�=q�eʔ�����;!M֯�ȭz��M�����
W��a��t`Ҥ�g�y���q�:H�u���|�&�QE�;w�/Ɵ2e*�͛KZ�I��p�]���3��?�B�H��+������ע��6F>2����;�I��EjJ2��ݦ���|h�5q��ȓ���I��!��K',����:M^ޑ_���	|��Z���B1�##��۝�r05W$l����8�B�N,�Iހ�J����' �/J�S_�ڣ��&.x�e��(��"7�*�Iy7o��&b͡Ѵ_'�njl��ODd[{�ƚښ�#����[6���_~���9"++�Q��`Jw�/!�3O�>�]��Y��L�7��ko���k���p����pZ�)Q��xxh�)::�ʪ۳��8]#1OS��M����O�^����u���?��!���Ν����8��'���+���@P�ND��A�A8}ʳ����ښJ���M��ň��6H�0�Ӷ�6��tO���7�N;K������8���tM��xs�;����E�z�m���\�Z�
���سg��4h�����H�!��$��|eeR�S����QB�Mټh)��$]��[�FL���N�)��vΜ<	U����oj�QR)NK��)Q��O�:���������xxe��YڊY�f��\���
6ף�U=�h4�0L�	����X̴J��С,� --��rd�h,�댜��ֈ�=ݧM�4�l����3HO�'�qr?�z�̤a��V]]�.�"�N+�O:N��=%㷐����Ǐ7��\])�P(!��O���A^�)x<F��Hh���?�%@5��um���a�XwJ]��>8s�,��\�O�(T���B�_:�v�SgʆJ��Af��#G~�\k׾�}����S��=6��`���0���!�Vь�
v�����xq�s�x���I����M����0�/��D=͚V�f�'v�Fg��h-�����6��3U��u�Ug��	0!7|�ÿ�7�ǎd�p���P���.l�*$�բa/	�_��Z�_n�x��#�8Z��]��H�I���_���rd�!
0���(�hh��ǵ2��^9uZ�&aW�JE���?r��H� ��:�.Y��C�a��n-����6G��R��.�7	o�G�=v%�;��R���P���5UqQ �,l.;�Iȹ|h��		���_˶0��w�v�ʕ(,,��I��rs���2����z�&�Bμ�f��+�Ā��m��	i=����������ዬ}�Z�qe%��
h����E~��w�aPt��x��[[��|�n���w�Gq8\�'�ݦw���!{���O�g�����m��	�"a�S���k�N���6.��W�! �Z�`�a�P�t"�ھ�s9���#�n�ٿ�]�����_{�y�ݒ'H$R�w�(�w��t%n�����)�q��wEX)!g��/�
q�eh�e���D\�����h��䂗y�
)b�L" #��b��\cYBG�����x��?}���{�+nc��Y]

�z�����I��.!đw���I��3����R�� �:�Ln]�d{b$��p
�и��NLW|U��G;O�=��a�ޤ4�w-[�={����XxX����݊J̕��v��tEi�-x+�2B
^y��霼���讯��Ҁ���VTZ-H��C�䉈��0���l������l���W��|�#eӦMx�Ŝ�'�	
B������w�A��٤P��ۮݺ�-���BC����V)cq,Z2]~�| R����D���f+T\��
V	��+j���.���{ ��-���_m݆��,��0��$�IlU��-9��j��'��kxb�̜9ފ���s��x�(��K�s��Ke�&��p���O%��X݈l��r=��a�j�jU�����:������ڶm��ك��F_)F�*hBpp0����]Js'	Ỻt��˗�͸焸���12i\?ȫ*�,���\���as8"�Ƅ�kj��aCTp�ւDy�i�:m/�kEƌC_<Hu���#t�4]�OM�\.�:����cr�3�c��w7�<�{Nȷ_FtZo�	RG�Y�3��Bf��<y>��"�P94�D4���ok�oAn�"�� ��Y��5r2#�N����ҥ�>�<�h�"]$�^��p:3�\�����@��7��J�ú�D<��
[ޙ�Epؒ� �߼��.Ȃ��ED���=}�|c�ڳ����^������s��Ԡ�����Uj4�Ç?]FLR1��jܦ*,<��l����D���?o
���I{�-����a��� �S����|��T�G��OA=�77�@k���f��}�\���$�KQ�cȷ�t�ass�{��2t��К��J�\t������۾�-�)!F��`�ۂ�3���n�2�(׫a���id�(`(�ui9\C��W�UՌڿ�����Q�<t�eB�)TWWO�~b�ȑ���ށ�DWMMM���$$t���_�RDB�
x9�)!��=�I�3mρ��K��jW�����Sш�S`7�pk�68O�-/�]n��ٳ����]��>�o�N
���:�%�ϗ�"��@��j)J^\\��4�wg�帧��'w��k�E߽{�8tT��j���ij^5wt���-=K��dm��M�J�ywA�YQ�En����lIh�����]^@�҄"5kV��e�X
��T��{J�O\�Q�;�-��]���&��8��l���C�+��s�g��>r4"-4�~w��6*IH+�5�̧���FP����&EFL�����͔fx	qe,6���!�v�%�0|�D����?�aovL���S'��'��'B*i��B}�{k1�0��i����`2;�h=����϶����y����lGɡ3�juc���o�%ir��� �1�0�5D�m���O��_oH�� 3g���ˏ;2��t�@���.�DB^��^e�^f@�J�,�X�K���칽���HŰǊ7��������j����w_��]�nu>��q�1�/�ŋ�Jt�С� 00r��V�)7�it�#�	��vx�(:����t#KwO/�d���EL������HI�A�\�a0�T��Mz8.�ޟO͹�����z��Pw�V�S��BTW�����Gl|$	�t]������"���Q��9Bh_�"�j<or?d8Dwg@Zj/(2�'�.�u�
D_�OB3�4  �S�^�w�UB�uA�y2#��|��.�����ʝ
��[��m�)B.]��.�Bz�������������QQK�tS��jʢ��t�/�g����ĺu됚��x]]-f̘�^Cͦ���fter�٥�X�,�X4�z�/�g!n�mz>��>�ro���Vr���q͹T*�+�v��w�%�!:��m~�:�p9)cc�&��nXI7��A{���o7��D�{�#&�%|��=�f#�O��8�j��C��z�&�5q
8�}y� t:�'��*�^�s��'�a.��FAAA��}��*�W��ӝ}Hlq;u�M��aߩյѭ�����>AM�Ӛ�	#�L�,9%�]��qY���bh�`40\�l�m�J幏����	B���d4�tKIq��!�aе�p7�m��|8F��$!��zBh�DkZ�&�Ӌ~���>t�%%Ĝ�?I ���ӹ��`�d5C�����P?@��q,	s�t��ś#��^�wD�p���r���c�9�Ey��9�%��
Z�#>�49�@�F|��~X�|L(���D4�-:�D�.L�*������9��j����l6k��nK2�n�l�^&�᮵�2��*�=�l���h4� ������i�3�v�D
�b�I�o�Z�ex=!�3B(���.%����B�X.�Y.�+���W?�֗������Rm�S/�=t�:>Eȿ�v��'�g	�O�������$9    IEND�B`�PK
     �8�Z�IQ�H� H� /   images/a05d3615-68b8-4f26-98d6-1aedf7f6d878.png�PNG

   IHDR    �   �T9   	pHYs  �  ��+  ��IDATx��y�\wu��\s�y�,k�lK�-� c��? �uB @��n�{�^�������t��u:Ƀ� cc�8�x��³$��,]MW���C���޿SuU�Z26���ǫ\�N�sꜪ�����ۃ
�0�0�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a.A|ߗ�)���B�P���J���0�{ ����@a��Ŗ�����r��������`?�5�0�,����N�W�������iZ��z����ҳ�|��D"��a��s	1�߿|tr�s���Q�T�d2���{�?p���ѡ�J6�}���)�0�,���o���r�Z�POO�jU�T�uatx����mKW,sS��\o�$IE`��5aq�0��m��gδ�Z�J-������N�R<����v��=22RD����0�,�azz�xc���P���ƛޖ+����4X�}p��q��7����nKO���p8��$
�a�%,������~���N���yrl�s��+���"555������ٳ��}�ۮ޾�����SI�>n6�0�s�@^ ���LM�<����=p���믽N�,��L&#B4��Y�f�'�����G�����0�.`q�0���_���O?�[(����r�
8v��>�&�-mm�-d2((v����a���a.!��{h쇮�z��v�ڵdrr���ѣ�U�VI����b�

P�_y���>~�6Ӳ?====�ۜ�
�üSX0�%�����=;�$
��7�|����pgg�433�d����=�vǮ���3�C�P��f�a���a.E�!��o~j���[l�L�ڵk���_���aX�x	��g`rdL>����˷n�T>�'��K(,r�0�+`q�0� 4E��n��������
�R��C�گ��r9뺰a�z8z��42<M65�_�jտ<5X�H� �0����a.Qj��W]]��K��r�����Ύ�XGG�l,Z�����'N��6��^O�3���Y���?`��`q�0�0h�4��g&�r�С��ǎ��áX,&���B�P�&&&BG��v�u*�JcR��3q��a.����)^{�5;�3�ec�m���j�V��֬^�bQ	���Z�?t˝C�g�QP̼��\W�,	`�}���ĩ��^qŕO�\*���������-�_~���a��+��*��g�Z�f횛GFF�6�^��>E��|�i�=�t��f�)Y��p
��aq�0 *r�F�����O�8�r���m���ɞ�)���͛���#����MM���ݝ�'''���tc�|2sfo�[,˺�Z��EQRUuPӴ��z'�9�t0�`aq�0�&����t:��jV���߿���I�D"���
}=����8}��X8�A��"%0�ܜ<͹\n�U�nnFQpY"��9�#�c��y��m+��n3�E�f���a���r���'�� ���7���~�5׀�H�b�2p\K)r����ݴ�MS��ər�l!C��߈F���lB��ڎ���@UU߻�4�2�=����q\3�a(,fQKo��k��;/�Z�u�\{�T5�m��v�
��B7���+.8a�nދ�.|�,+���wM"!���
��L�R����p��Y��8`�l�#?:|�p�i[+���W�\)�E���Q��t{>_���*��Ln7U�@@�!K2�!�hZ�_�l�fڲ�	|}�Yp�8`��Lqr�J��M�f�099����CC�.i�&]u�U�
%#�0(�*)�"D =� -�s/|��8��,�
����)`fA��a(���ɱ3g~���O�I�ǩӧ;.[�B�m[���b��h�%E�a�1��s}N�쁿���O��{��9��,0�``q�0��KO_�e�c����Z]�������)�|ŀ'��y@x�ބ�A�=M��Վ��Y(�p�����a,fa�ߴi��KO$���uv@"��R��,) 
���Nh
b�tN,4�Nz���u�ӦiNR $�l`����Y�DK�ܒ�7o�VJF"�$��A�l��jb��Q�����I���=�&�$t�ԋ��#�ju�q�Gq�)��0�>,f���:�N��ˊ�E��ׅc�fߗd2�� �\|���g ��S>	|V�Z�B�!��Z�"a������f�K���FI�J����߬����Mh詎�䐁o�6|�&	�c�#��}�����\�P������\ڰ8`�f�X,�D��m;�Qej�1��n��3p�}�Iel���:5��܄���;����e'X 0̥��Y �AVL�\�#�O���Y|�j��뢠3@4�=_4����q]�������Q۶Ǫ��p�wpd�K�p�8�s5�[Ѽ/�Q������9���y��ϧ�����ɟ]�:�ׇ�N�P�1\/��s���a+�8/S$Y�gУq*�h�v��B�`��hX�e;h��Z)����S�D�|��\R�8`��YlŀR�������!���	i|o��|�P4� �J����(�+��4.����҂��,J(��>7�Q����+A4U��9q���_�B��O*~�{n�뺷ض�U�����0sI��a�H$�f�Xڅ��OQ��>��yq��xPh ��|�0_0ԧ*(������J�eY���3(B����r��\�8`�^�Jk����x+ǹ�v�����Ms��������&4�CC�@��A6
=�oe�a����(�r�5E�uY�J�&I�hOo��L��M'�/ˡq�����RE�!����m�\.�p�0sQ��aTW �ϸ���y�qqOc���8�B����Wy.�H����]߻��g�u�ه�W�a�����	���#�[��[�{�'�u[�=�ι���[5��^�z��Z���y'��
��MӜ���ZE��(aq�0*]���UV�k�NG���&Y���n�68����d(�w�����qD����j��(L]���b��0',f�R� ��d�Xf��y�qq$x��ޮ:ⅶkܶ1てj����{}T �X,ڱX�Ǹ�Is���a6e-��]{��x]�z4�[�$JA����.�/.T5�͈J��k(��`�;���MMM��7ib�������Q~��/�phE�ݥ+��i
�@A�2躮��+�4�<����yu�K���`�x|ڃ�������r�/����g��0,f�S�?�,�Ǖ�WU�8�o�m,�BA���(�}�`hl����4�]�y�������xy�1����ɑa~��8`��hpM4�of��ߗ,���ֿG��0��l+���c �>ض='v  ����ynm��ϛ�|��|��a�r��Eɕ7>��ݕr���Ͽ4���Y��q����	U�*0���>������L����Rp�(dr�׻5��Am�s�������iv�$R)UEQ�Ȓ���������t:W��F^3B�nLƓͧ��O��L{GW������ӕij�͵��J /����yoaq�0��8�����3�R�r����#�rE�Ѿ��a�1�V�5��*��1�uj��`VC#�י�ڲ,P4U��׮]�����{��}wr,�y 9z(l{�p��(�jF��ɐ�G���Htd����=�7�<9�޾����apX,0�o��Y����cp0k�#��?���N�ON��km�X���?�E�Qa���
TiYUE���&J����k�<[
N4#����ʦg`떭��'���Q<&ϰM,��_U4ח4K��vX�z8�?v��T,���G���@wg�Xϲ��^:8�bE����ms�$ü{X0���N��g�LF}������gϞ�K��z�f�öݶb)�������[o��L
>$�@�MSg�dy������.Կ�B�R1!
��I�X�=�̧�3�w�^(JT>	PH�l�>(��)P�"�}q��\�j�u]�:3tf�8:�H�ɦ����S?��g���+�[���m����a.q������`����-���wMLL,��J/.��K���j�Ҧ)jҶ���h`}%��}�1i�������xL�"�N�#O1�Q?����<�;�q�zV���P(��*B�x��p���3����8z�$(�g�Y���B̊Fb��U�Y�ͪ�W������bq��"��F�N�'�"bG^K&�wv���w~4һqe��k�)�P`���a.A� ��n:p�`����ok�F�7��ٕ�Je)�4�8��c;�e<�" בh��� �-�< _��W@�Chl}�90���۶)�Iz���|S��0?�1v��2�TCx(Ц�+�-|��
��c����F��2Z��>�Q�+���PJ|�mEQu躱f:����������p�T��7����{�����yۦ��M�*��0saq�0	����<ff���R�Rq"�J!659��=�tb||�����.,im�h���	�1W�#zڶ^�@���1M�22�U��R	�=
۷oU�E�D�N��yεan|��i�0���8��%���72���>�� ������
D�(T�.�V	TY��b�pI���a�D %��V<�'u���^�Y�W���Ux���O��b���v�����+�w�cgW�X3y�5+˸>m��N�a(,�wL-PP<N�)�T+��v��X�Xnʤ3�\6+�*�b�/�Jm�|��j�=8:�r�-W���M�eEhXMF��zH�sf�1P�"�����T3�a����ˠ*:\��*0�*�b(��{p.��x���������x>�J��1��d�e0t<�H4
�]w�9s}�Qp�*'�~����Y�$�*:�O�k��b�(>,!�$Y�D
�,�QUU��Uh/ds˓���:2����斖�Ͽ�����W�=p`bfӦN����+,�HMh���J>�)�܌��/^NNOdZ�Lrb|��b�ڊ�\K�XjuL����}�˄�Q�uBh�YQ4)�U�T|�|Գ��QxN2��xVE�40MsN�CZ�(�� mB��?ǻm��(.p�n�q�툔ƹ1�ԹPm����gI���b�"� ��ڶX����;�ؿ?4%bP�V _.B<���5�/�dA���9!O�Lr�t��@"��-P6�G!611�k��`e>_�ahp���w^�d�%˖}��7�-j.,[��
�>��ü�P�����1:ZR���н?y�9�IwOO�:��T[�Xn�V�N�r��i���q��vÎ禍�+�窾�ҳ��XW�?�t>Yמ5Y׫�
S(�j�p�v�aժ"����+>0�4�wl������~z�����]��7�S>�e��	��8��q���>E�Z��	ρ$����j�H���?��?���I�h<��mUA�h�^|���`n�%(��~�c���,K�7%
I�Y���b���	w�������N�<z�С}�]��~��cG�_�%������	���@���q����F����?읙ʬH�g�Ke44�.˲�M�jv]7����8a��T�wd]�4\�纒C��vJ��PEc&Ӵ@�u�!a��< �0����Ā��{~�?E�hov��D�ׁ2r�|����/�#�(�b?7���7���
����H�F��P�`9�8� ������+����������T*�$�(jtm�{iv�z�sf>�x)\q>T"�P�
ϊ(��Ir�\
����IF�����m�|qpld��=/�z�����OO�^�Vb��,dX0̻�����MO�F�����\��*�έ*��+�k�eU[Ӣ��
���9.�G��8��GE��/�A�U��L����퀋�Y%��	����;��P��%90�$l���>� j�D�PB�q]Q��R)����r���0�{��կ~U��M�U��ޮ���,t~��H�j�!�2���]�m:p�m�é�A�� 33I&�Z1g��ll� Iv���et�D �{W$�P6F,�/5�r�!k�)I(�4�zPmɑ���^^���㓩}/��煍���{饃c;vl� �,@X0��PL�ӑ����ӧ�7���X<16�%�/l�Z�R�v�Mӌ����<ϑ|r��άAT�"˵�THH�Q�d5�'(�-o�*!5M	Z)S5"_RE0!�m���ڲ�B��ߒV(��؎%�hz��I"��VEݡ����@#,�+�g���������g��c�D�2��m��G��;;o b�������2�~E�$����)����*��4�N����c���ۣ	C�< �H���<�WM$���3@ъ�f�s�߇�S(���sS(g�+䄩�I+�]5[3�j�m�k��ʭo�y�����_|���¶mW�رe��͜��,X0�<�=���/�>����S���^115�ɬV.3��b�b5SQ!�qu�����y���P!�"�00�´��� 9��f�$QP�k)�@)X�X|�rA#AQ�����P۷/l8}��@1V�
h��p*"��rac���M��ǟ|֮_W\q�a;��W��|t]���˵�<d�g:�;���	^�q�@�B��h���1��p�Cc�Rׄp<�������o01>��hӪ�?m��!�C�0�*� :N��ǎ�A7T
[������Q$�o��IU!�h�����[VJ�Q<If�q�Ո���K������MG�ϼ�kס=�]w͑aߟ��E�EsI��ajPa��L&���cǏYy�����c���ʆR�؋>��@㡋�;*%�F���|`(�3��ED�����hZ�|��ʂ����9(M,ׂ�$�Z��E��#v?�{�����?�.$J-eq�O��]����j (� ���-�SY���?���X�d��D��A���u�z�m�ߎ�O��<B��h��д�iZB8��9�������s����N�ڣx)�NQEVB�hq Y�cR�#yKW�o48*�OFa����#�lQF����x"�����.������a�Z���ry�L*us���W6�]��͛��I`�K���z@�ٳ��?��G��422���-�1-��X,�H��5U���a���k�
�b�.QF@��G�pd�g�.@)���z:a��! "����G�	NCϠZ��'R�%:����uP�lց4�3]׶�2��O64;���=����k_�Y}6f��5�0��eatϥ:J��s����A��L>�룔CD�\?I� ����J���F�t�7���Y
�
���Z��:��!(�����Bpn{��,-!M��=��OB�Ѷ�k��M�q��Wh��1H�tPtX��B�p�%a��Hy�����w���g��9�窫֥k��撂��o���`6���ϵl�*�No)W*K�i��+?5��@B�fٳ)��T�;0;�f���y�l����{�za�Yٟ5�AL�$�	#������0�s��8?�k�( �yhA�HJ�͞��!bD�(��W^ރ�}�b�vA˅�u���_������
�8n�!���g�@�����ct�@p}��O@�����C���%!À�U�2kͣ�`��V��i�8�����bʄD�n���!/�{ �`UM���9�E瘌G�T)KN�l�pn�<99�慗^�x���������cGV������os�0!,��d�O��h���^r���fRS�s���R�ԍ7��iV)�PRq�Ǹ���l?
���8��r�fH6�n|���Xw�i������O�����?w��)���v��3�l&���~|�K�4%�p�"KA�������2X-��:�kqO?�8\�b�y�P(�D�^�TA#���P���e��9N��\�>�
�7C���{T�� �}����/�Lz^|�e�¢_D�PD!��Y��7J�9[1��C(l�QP�e�h����A�b�@A�a%,�8�A^��G�� Rׂ\���CXā8�)�U7i��_S�VV�3�kO��y���<��y��̥�f�CS##`�����5�����\5���ʢ�UIKyݱl�^+@����Oƀ *���`����s�z/��X���˱���{Pw��s�{�'�a�����Q��W{-��{��0u &+j�|�e��p�$P��є<1M����b=C�g�@��o��r�y333�T���������|Ci;��@�Q�A)��Na�9�Ba����կ����#G�Vȗ!��x~�H��oצrPp�A��-'����s���s�A��Q�p��.*���N#��PE1�P�ExT��S�/��Y.�Z�7���=��={>���ھ}� ���A����f���I�ƞy��%{��_sj���B��r�\\.W���h�]��H����>$�f��A}��ڵ�B�TC]۴��9��~-Q���S�c	eC�`��	����6�C��h�f=� a�w_��O����'�1RĜ�^��"�h(tF�Z�őoEb����r z� {����_��?��ŋkM��N\H�c�k5/ʹs��AD�����EJh�R�d�@�2��[��������߆b����A��F��"�rD삅�����9A�bѼ��i@�<�p�=�� ��bP$���Ȯ��z�Y(��R��� ���D"1��PO�>ٞln��jUW}�_��a��-��r����;������aq�,8(��ԩt��gw_��k/_svdt�������k�V�0��j4��-�T�Y����Q��f�����WRɠ�ѣ�@Z^�m4;Z'�������@BW4H
�	/�7���TaL1� ����T�ǥ�*%��a��$ȭ=�W�e<L��?q����Y����C*�R�Tq�h5|V4J�-Q�@��Lqd.�8q~�!��~^mk됳�4O�m�
ޮ0ҬGe��������I���*9�s�\[(�@T$��\.7\w}�n����=X�h�:m�YAQ(�#j8t�����w�D�	�޶������"���V��jMϚ��H؃R�(Ĕ�W�T*����6K���n�U-�p��l��ɗ_|u����3�����TC�"���`����g�?~��e��vxx��\6we�\�T+aJ��xj���ԩξO���1d�E�M ��^�hnoY��:��t7Yֽ �'զ�Z�Y_*��6�F�D��N �H����Z��r��pc/�)�d��*�IV�h�
��U|��--<N�r���2���G��LU�|Yu\S��C�\���Q�'\/��ƣ�$�82�*���T��g.55����?��><_=v��=��H�,2ꁏ�쌹M��ޔ��r��1�Y�q[��<t='Rig�����ю��>|+�>5{�|C|_MI�a*(�(2�f��������N"p?���@b�T.@��鐔�IS���`jN�&T�}8d��J(^��uܠO��k�6���ߞ���V���u�cz}#�Μx�����׮]2�����fA01�G�ӟ/~��Wn��*W7U��b�Q�mQ5��W�H��Ws�����_��Ǒ�"��~E	��y��A����\z�Z ����BR- P�\?�J#�x(V� �"Db�Zp��ÆL�>���h�0��e\���D��U�d�Pȷ턌�/��*�Ȭ�)�~,󋉢���rY�UcR%Z�����FU�]W�ѵᙾ�z����ѷxqxj&�t5����ζ��7~j�U���������$l�Q�\����^���3��0�=��x^E���8�O�]w��)���x��7�ﲈb��2�T�ihjjq9\�4	�@l�ۢ_��X��]'͜,�W$i��(�^%]x(2^�������lU�%
�pmoQ��7�}�������~���pW�T��`q�\�P��������������O~�Z)o-��}�B����BU�Dq��\~О��A���sN�� �M�Q�?(X�#�-4k�`BGt�skA��۟�����i���ȣi�-N�R!赨`XE{4���jŪ��$�L��=~!�;��躨}��Q�?��_��ըST�ď��_}]X�#G�H�j��f��J�ӌ�J�T��G>���������x^j��-�)�AT;Դ��&�|i�S �@�Dź�o��P��(� ��
@����1JX�PP�ҥ��;?�>�LMM�o��Q<x�g�Q���<��B1��R�Ez$y'DG
�tqb��8Ӵ�g�~G�D��/x�/�¸O_�Q?a
Y�M󅸠�J�xB���JUA�8[._��=?{�E�O<<44�Ғ%K�_�{��s�Q+o�����������������ƶ�K�n�4C�dD�!a�D|�hhd�g��A��J�6d����p��mhI ����IRP�>I�����%�I<��	C"b�*�khZ.��'�onjy��s���ֱ?��g��W��}��"��4���zH|]@� 9�̩=�wUn����E���������X^  �|��է�m^v��j"k�^�Z�;D���xG��{&�	~�BZ[��hJ�,��*XK0��.���B�jA�Ԧ��v��`^Q^ڲu!"Qb�D�a��@>_�!�e[����-��DX��K���(b�����R.��NO?�s��O�x��<�20��	�%y
>���+�nس�����m�Ym[V�q,���Z��h�a��=�0<*l�(��0ƞ�\a0[���jufk4�B&h$K�Ĕ �M��
�!"�3���w2�3�I�g��pKy1��Gc�Z�	�a��4����D�iWgk뫋W,?��������4'�������o`����t�����e�����e%VdH�.���-�#�|	�S��R-�VtH�RC���r0�	�B�Y�	7�FHgf`���� �~E�!��bV-�E��k�l��j����E�E�q�H��=�oL�^_��BH0">!B�!SӦ	�����b(�`h(�~�T�����QI4Ғ�R�Q�hR�`G+VeS�,7O�R���y�̙�+K�6�$�E`~�8`.R)?���O�ڽ�����?��f6y�ߒ��2��pT]�J�$"��0QC��< 
��R�57�*�"���wj8�r�uA@�r/��!1@��6��e'��´�6��'�E �L����P��dss���Jɲt$o�ݷ�gOO���ɮd���o��q��?����������{���h�7��Q�,��J33�,Ղ���Jsl�ыs���S��_+*����.+�(loi��n���'���~H6���B!_���$�6<Rc"���LĨ�!�m�l��b�=�**_JjKA�.�E�U�𷌻� 5Ҥ�K�&���Bq5bb�T(�@��>AҠ�ۀ��B��4_*|Ҵ�%�ӹ��n���x�3�����aq�\���Q�}�o��7o9���L���\.�XV5$��Q���i�������v�FA��&X����؃���"�*��C���u� !ewk�pBAjE�Ӄ����'u(2��+̺�ɕL��.��B,�1�E"�#�D�)ꌮ��Q ��hɢW�-��Hk_k��k�����hy��''�3��"����{TU��z���;�;7���P6��p�R$�|�E6	���)p�h$��?�}�m�����hSgO���*"�0�=-����h8h�q�^�*�\�������~;��,���%y�MOA�P�b�ԕ��(Vb�5��"�!�{CQ�EJf�v�Lu%�\���bW)�U��j�fs��ڻ�urb�k��|���X���‹�9p`"�/����W�������ǭjue�R�;���t͓/�?�����!k ��J`|��)r�Q�ߩ��E�cIt*$sF��*��Ǔ�PlO	'Ƨ�  �@Gt��FA� ߝ�y
JyJa�@��M�c"���B)�0�;�ڟ\�n�e��N�A����VZ����{�qQ ��G�����Q��Huό�/@��T���[������5n�7�� ?9��[���"C���wͺ��?	?���0x��vt�)�1�b
��u�MS
���JE��AmI	���j'mU/�Y���G�ñ)V�g����A��c�C"pQ��e��+D̄���,��z	a�钂?#�Hd�N��-����x��͝��,������]�?��;&&&�ڌƶ(�M�%o�
����\j�d:`��0�AM����O�=�f�TE�u*���e��3�lK��baHă�d2)�����Af�u�E8�o
���4W�ɦf ���oh|b��FK��O$�n�S($��t�<ӽ��卛7�����x㍮t��-�@�v��yptt�h�ۓM�$QuH�Y��<�$�ZNC�9�K�l*�X�X��k��8/��������p�n����V9R�ѹ;n��������B6�CTKb�!��BaP�K�׌6�Ēq�.�H��G�8Ma�*e!--����U˦	���&~�[�"�b���@!�Mf��k����ɢN��RKQp~򹝿hϗ��ʾ�xq2+q�[��sQA.遁L�������w~2�/|o�K*�r�����֩����oǱE����D�]2|ZW��6mP�F�e1@�r!4�Ѧ&HD#xS82<~�x��n���Z����(�8P�b:����I��H�z/P"{H�E�zKs����D&��M�Z��_\�t��.[zjˇ>�_(7��n����K_3-�>�=�Р���VI

I�δ^Itj��|�[cje+�3�S��*�`�uES+j\���L*���18s��~m���o���e4��ۇ�a O���N
	��{:;�W�Q*	�IB�zo��us{+�RWd0T�Am�z�J�n����O(WPp&� 7'�ukj�D���$*����[�"��l6���-�w��E���c�(5q�.��o�Ey^}���Ǟx|������Mss�TmF��j
�bޖ�J0�o��,5N1J��63�Q��uZ�>�@��|5@Gk�XF���itK7���q4�i�z��i*���ֆ�aH(/��ffҢ�yL|M^g�x�K6�MCקp�C]]]/�Z�b禵k�mߞ[�7�;6e�>�|%ި��gP�u�m��F�%(��[�qnan$��i��M34�;������k��?�y:sΞ=+�4� ��UMa���	�0�hTą��"<?�"���G�L,�g�g2����"���,SLC�3M'Qf�ZUA΁���zkio=���ɐ��T���*���W��ײ#3��K��;��any�����m����Cu&''#߿����~m�S�K�dW�4�j�DM~tQ�>�"H��4�o�x#��Q��m
%:R��2�� ��:���0mM�D��(Pd�0p���	Q�+�X�ǣ����d�ZZq��(sLƁK�F|���

���h����k��� ���֬[��UW[�}]���`����Q�M��24�7���om�tn:�Nc���x޺,ض��<��o�o��߫��>������o�Q��h�wR-ѫ�
D�d�P�		9H7��lTJs�,!(���c4�,^?�lJx��Z�h����k��)\i*$��B �,�R)(�K��� ��<�a��Ѝ����|�)[�߇Ǻ���y�aq��^�i�Çϴ?��/�<|讱�����b:�([�M"ؐ��m��_�j)v<�zȊ���" �J�����������XBx�V�,�Trȥf`jfF�S�Q]kK�H3L4š��]��(��摋Ŝ��g�@PZ����h�PL�<\/g����z{^X�l�έ[�8�#�~���������C�m=��<�YK!%�!p�@ú�k�+᭍���A ��A�OC�[7�rIu�HF#q�Ƹ}�v��=��?��?
���f��h���|��2q�^�(1�%�9wIp��Z���X$
�x��:���C0�Ud����S$�@�H���,6��rU?�~ҥ FEdWě�Rl�����V!_��i�ų+x���1-����h����?�Q,~x���Xƙ�{���	�_�b�ҧ�}���#�*�JWP�D�H����61�K鉸\�/�⨝*�ջ'J���R�o��B����� Qmr�8J=pto�HnbbB��R*:
��!F#?��Ǜ����]#���M4tL3S8��S	�H����� Q�e�9����V<z���;/�X����>x/X��;3trh�6��Ԍ?Q����|��0����*+�g���oXQR��Pp
�M�ͧ>�)�?v�~�9���MO��� �P�K4̎Y��U�dSb*���j�B-�mk4�@�alj����J �#195�x��~S���n)`U����9�c�Lq����G��0���Y-�EE�H��I�T���车U�����5H	���ݗ��yaq��^���w����}{^��������2E�B2U����pТ�J�VU�򫢙MtHq
u�U�B�� 4W��6h~D��FnY>2p
�PP� $j�4D\/�A��M��557���/j#PQ�RID��(�<xS�D,m�-~<�ú>�D�.Z���[�z���݃�n�-�O#�)��b��c��u��(��VZNn6l��l�N�A�՞ˁ���Wj�"�7M�U�a_L|�K_����0008[�PZ�ق---҆����L{S���c�G����orrriT�]���}=�DE
e6��kp��A���B1��,�(b�P���1��)Q�Q1���E�`�z��G�iV��~ʐ��@8��q$&�4�RU%��ڕ�f>�п>-�$^e���W�8`~����������w7?v�+�t��|�؆F\��w(���tC�n{�X���V��"����h�d ��T8���MUՃ&9$
h�`bj�SS����J�bF�$Ba!D�MM�l�GK��|jDF#�J�:�\FtdD1 �j���X46���utt<�n�ڟ_���S=[{�>�lٲ���؛���_R*�-�H�� ����_����A��x=D��^S�B��������+��TV����<�z�b�
������Ѳd�kP�Vn���Rg{������B�����%�+��(����L:
�L
r�?�4�?;x'MS��2SL���SC.BTJtA��N�B:�Ϥ�x�7@�Ϥs"��,r�U*E�q�m����_��B�\*~�����d~cX0�3h���7��>���o:t��=�ru{�Zm�TCҍ +�R�(�����q���U�C�)�V�_��� ����zb�6�H���C
B��w
"�M5��TD4�7�HD���n-�{�5��Y&����)���J,b@K"�F�6B��X��u�.n˦��_��ʴĩes #�>���Ǥ��h	4�78��.j�,�g14"F��[c�?_|B=��\�c����J�B�p���'��<p��P��W�-F��׮�[o�.�|tvv�`��HV�2+����E��S#���Ã){jq$֒���D��x=����*W�05=->kzb�[�`E�dsi�ΒA��f൙�r�ik��r!�G!
�~bA*ff&hU�
e���@\x2�K:�*õ��}����}k�7���;���/~�g����Α�;|_Z�#�D$�$/(2S���R*�r��`�m���*�b9U�S<Lr+2$��%D`���(L�S�k@�k�ǥTE�#)*t�����FH$�Ќ�Z���FL�]~vpH|��b$��M�����'�蛫��xt��5/,޸q�F���������D�%O��4���	�1ly�R���w�A8�v���yQ�P
�FS`�=w�G�ݯ�.�_����[Dzbooo���	W�s��:�Wo�;��3����JQ�]�4�D�K����o
��j�S��a��P.W�U[k���A�X�X+�����#�F�MiDs��l�w��j7-I!1E�{N�X*^�ƛ��O�����f͚0̯	���<��S�=���KOOo�+*�J���C�Q$����W�V�T,���4E��l��Z�#Q��v�W�
�)�#�ֆq�f���a�HMC�Z
B�$#�����(���Ơ���DZZ[EZ#��IHЃ��m����ɸ��r�p�Dww��׮~~�Ƶ��o�R���\��@��,?��vX�?Gc��1�������Wm,����=�'�V,��~.���_������Uk׉��E��i�&�K%�U �V8	��/����涎�.Ӫh��A�j$%�Q`$arr
�S3�T�3�NCgg't���ؗH8.�_z���c��Z_��������6Ҷ�r���N���8.�[��~r|d䆗_��W�����y���uaq��V9y�7����޵��/�R�����Eh�d2)n�� u��f9�b��Y+Xt��)�P49��8�
�<����tZ�Q���*��#>2 T'!�Bkst�����o��m8$*�Q.;M%P��4>���CKS���`�9���⥽O^}��=�V��K�]Ɓ_�P�{Nf�3Ϣ�nſ�������lj�AO���=ۊ�����z[�����H �s�=��栫�zz{�Qi����"�S�+��J�H4��g�ݚ������`(���*^��/�]�3�����@�e5��/����
�J-���G��8�\A���k�>�)�[�8�CA�O�I�%�vԞ#���k�Ϻy��o8�iW��n.���:�8`~k���=������_����z^��ky�b�i���(R���ܰc�J��"�%"PYY�r�D�#o�F0�k[�O�ѠO��ii��4G�Ũ1R$�H7W�p�����6Q렊�L�.5�ނ"��ɝ�ױ�����DN��5���˯|��[N��^]������&����p܎C����.6*1(`T� 4l7oGs5���m�C�
��3�0�@ ��iPEF�4&ZZaђ%B�E|@�I��>*�p�O�*�JEZ�ti�=���|��+sz,�LLNNJ	���8������)zp�x�ҹ�Q,dr������.���Y�,]��#�K� ITM[�%U�L4��n��5�MK��<�Yʰ0��Hu���Yv����-��uos	�}ü[X0�9T���ё�'�������1��?����PHr$#y�%q��*JQ�����s�7r����Φ�&�b\��!5(n�Q[[sRx�xs�75�͸Z�;D�"��e17LE�r���Fhom���ݜ���45������M��-7ޘ�)�����O�ZRz�Ԋ��{А�p��g��{n���ȉF�*ivu���M�N��sx]R�B0eЈ_�J�I���Y��n���O������泹�h�c�T�h?�{hʀRjQH��3�xPnPab���������C�P@�x��I��J�I����D"	==}�#QM=*f��K޴���$��Ԗ�?�󹝠��7�|��@`�,����0xꩧo~}ϛd:�v�v�B��7���F��V��L�M�7c���be9(��	$����bDA�VQD}�q�_q��1T�8��\/� 1��mCA�ln�ވC8"�$�͋N}cg��G1A�͉����R�e�$��g/߸���1��~��K��~ń�q���5�ؠ������~�B!0���!����\i�����B5,���۔Q��x�eW�Ċ��յH��G�7��Q�X�u�O�����3ӯ��{H�B�����zH

 �bz���:��@�}���$�q(��(N�X�x�;�6L�8��ʒ	E��Ŵm{�����"�g����Ԥ�4-��{.
˒�1�,�ʕוn{����d��,����{��=����gO>���{�o\ۊ�R"2�կ��J���aP�g�%W���=t����uP0hF�&��HoJK,�3�T�i]�Q���X�JI��koȝ�d�r���t|�ː�Q�t&��#��Ql����M$�S!#�ڢE�Ol�nǋ7~�F�|g󞂣�bz,�G��9��_��~���[2]`6�^��ܶ�� ��ߵg�����[�(6 �pT��긌�rR;o�>�uG�����`Q��jń�D�����<�?16���-�K�Ñ=��c������#(X�,_!�FF��3<�91U@�eہ\>#�=���բ�MoC���P�-Q�Qx҂΍P)�xܦ�.�l�J�"㹷ONx����?OK���Z7G̯���q����{����O��Cײ��Ts<�Cx��(�J��TZ��+%�e� �y1� +AT��A9��0A�4!��9q���1�j1���D%��S��h��f\���~�
~�%����������)lP�i��������Gn����5k2<���A��'S��g��V'�0@Q������*	�F�T��Σ�u�<ႧxѽSt�đ<^+����zA�B�L��<>���� ����0��4����d�+6o���g������r�L�$w9�-Qq���ĝ�؆<Y�P���x����!Ը�L4�߄g��R��Q�+��"��Jr^Tdlk�f�~V|o%�&Ź���"�k)f�����/��7��O�8���f~,���]�N&��ɿ�:8p���Ry�m���V����M�Z)��xT/��[i�&�\��%Fs"��V��n����A_��M��5E��4"�Ij����!a�N�b=}"�Х�
|�r���FD&B&�7Ԟ�Vh�F��*���xp�5W=�t�Ɓ��a?��54��N����Q4�[\�]��M����S�l_	��RC����/�Y���fcY��3��P+�$I��	�Ul>�܉���Oe3��;v�9;��'?y�4HjDV���TiBrŜ�	�ðQ��:�'�	eR3щQ�	c:ƪZ���f!��x�����ق��6(����Q �D�䂛w�tL�-T-�+��k��g���3w�noo~
>�6�8`~cv�������x��?3+�ͺ�������H�A>�e�i޶~3�%i�R^0w�:��>yHDP�"y
��R�!M!��)��*�QUCWEg<��mjk���KD�!Eo�h��f'�'`fz*��ՏE"^S4��C�+֯���mW��eǎ	�;ZZZr�t�5K�~�9^;.j���_�]#���Ku��w�9(���z�g���p�}�/���5U\t]OLM�����O]q��ɟ�|�P4_�*4���d⵬�A�hQ�و�؅��6���6I��Z*G��[j �u����H�¨悸��d�6m�򐸅���!1B��1-�N�H�X�|������ӹ����-ZT�� ,�_
><x�t���<��cG�|I���8ĉ�-�qӍ��@:=#F�d��P,�"E��d�k�4����0���΁�Q�WX<HtP�c]�7���"M!�uuAK[+(�.�f2i��LJ�<�����4c��YUU����k~���z�n�b1�B͡��x�1��7�.���DqQ��[�����{'�`�ƿ�S�u�͕��_%�����(v���0>K�x���_�ⵧN�znlb��d�2-1l���#!�����D !e��	�DCN��Rx���(�Si���H݃fh:����B^T�	jb*�+�Z�&j!���<ω����=\~��D���cj������;�����?�����f�Q�)W��Ǫ�*n���'ρ)��l�� Ӝ��i):�JےV��t�t���t��4��p(x��iZA��+ ���Ǡ���{{!����BXP ��� ��g�ÑT3��ڛZ*��nkn~bǎm?��w�.�Nv�/�@����4����mh�/C��{��*���5~�[P��h�����ނ�b>t͒'³qmR)�U�/������[��֞l���"]VTJ7�������8��M�~�a4�4��dG
��z��k{x��-���~NE6M���M����,�!�~��\x���NR�EV�8M0+���N7���]�fz��S��qNqd�����ԩ��'~���ǎ�Q�T�RӴX(�(�F:T7 ��S	Ԅ�~c��r��94�#A��(r����g����D4(K[�ѫ8
��3��wQēI�E��''�a||\D{��ш����D�����_}�U/�������q���ڦ3��gM���� �F��,T�^��?j����ԯ��؄�)�:�����F��hFA�xݫ��r�֓��?��Gٗ��C�X�C!� �y�c�"Ж*zRZ$�
u�1�LԲ�����	l
F��M�8��I�ſQ4��j~-�!/E.�#����U��MkEE~�/_yi0ٓH�M �̃��9}:�|쑟}��7���'yW�m7��%��Ho�(���%ciO7��/�_��=7z#W(b��<�t�bh�5�7=�g1��H������Hih]�����"����X*��atd�3)��]�ns"���_[����[o�q皫��qJ���cccx�����Pr�׹��9N0� I 	�Y$MQ��Dk�D�lY�]�ػ��>gw��d���=��dJ)J$�� &�D�����9TW������`8����<�驪����w�w-�����f�<M���=�)s��@��W��4�s�/�5�i����$ЪHh�=놡'���UÃ�����oӨ�s\�jq3��
3�c2p`Wm(
GX�, Z�	8S�MW��X׉Qk��*�-W�x־+�a7ʺ5h���Vh��oA)��aҚ%E�M}��_8xp��+<.ONx��x���j׮]_w]�JM�B�d�#zWR���&&&��N���	x�
hDj!_�����,�!��1���z�)=!<��Q�5�̤�I����C���Q�7�F��x�SCP.����x4f��*�g6m��Om����e�޴��Lh@z�{��x��!������?Wja��F�������4�A��sE�٩����0��j|��!i�W+e���m�׿���\����I+�+o�M��rV�X��@#*��@����yg�6�� W�1@C���w�#��ڠ6O�[��s,bA5?� �,��5551�N�J�y] ]�l˽��ɓ[_z驱c��K���'3����������#G�QU������8a�2s@E�F<��'�D�k��o'��=-�q0�T��q�5R��E�A@��)�`.Ԕ2MV��k;���Np�A����gs028 ��)0�{�#`�E#�ϯkJ�[�q�/.[š��fo��y*�x<_(^�,WrLK���*`�Y�7���2W�!g��0�y�F�<���s�T��\���y�Y�*�j����}�+����������g��ѐ$
+�%��q�Dj�47 �A`��A�_g�4�ltԁV�Z[�!� 8�녊}��]�m4^\S�h��T��K�]�Y�UR�Zշi���c��]9������O�IPq�����e��F6��Z7�H{k�g@!MPm�a��ZkOtL�G@�&̱v��O���K����yJl�z@�\c�|,��2��Q!�'���M�&����(>N� =>��B�E�"�{��Z���MOn��a�2���h4���(F�ڶ���jܬ�4ڳyQ ���#&�@Ñ�ㆁX��<Mot�R��ܰqÖ�\n���/5�Q��P.�[}��hh�� 0�z���z�E��x�M�%���?_ E����TQ�$#�f��b��LhGCl�T�2���E��y\{-�c��Ύ]'{{��L�'��<9A)>��k�v����Sãף��Rȟ��EY�r�����L�ͤ'QШ�n���d
�,�,���@�X��Ǔ$��&�C�R��-)Ik55CKk+�tG�i`Njb��FO�SթF�M��զd|_s"��[?�O_~����}r�Ax�l�f��w)����s�ϰ�UCp.���Pcu�BX���Ԛ0�� ;DB�����n�n|,��^|��Z�X:���c��������Z�C����˯�`Rˮ�9�>���B���{���j,8�����A\���g�U8W Ө�'e6�E��z��'n}ᵗN���/��q��x2��"�_y�ͅ/��ҝ�L���Z� �4Ԉ����P�qǍT$�
��,m��1���8 �0�����C!Vk�HE��ӊ���������l��%H���Xj�
��MNS,VD}��w��p��ǖ�[����>yR� T�um=��~����S9S���ɹx�g*2�y�3������t�8lud�����drխp˭�j�����������p����w,���"eHӘr��p�fh|��Rn"�n�Z#0N�6I��4�T��EAv��H$�p�¬e���s��D,x��6p���Zu`ߡ���}e��^o�x�O�#G�۞{���LM�o/JݡP@��l�+ f���$�i��%�D���q�z��>�N0-s���>f�} �e�F ��5�	�$���%���\���k�.d&3lp�Tz
ˁ�d�s>Yپ��e^s���-_�<�|b%�e��^���;�Z����Ň$�I�?��/�)�1!Ζ������1QQ$W���B�~��u�&�|�X�/^�h˧o�퀪i���Z �^1�(W*��a���y��b�p�bm���X�Q"�C��PR:a�1�imj�A��B��B�F���F���Ǉp�my	�4(ҸSCЁ�'��~�+/�xtq��!��/z���'g��a����?\;1>�y]3�P�ȑH���?�Q��9fƞ�U���V'@����e�ުH�� ���R���(� K��,(�t���fhi�fT~�`��l� #c)��Qↅ�椃Ǧ�>��+._q߭���jOO���>�B5"ccc�B��$>O!��|.:q;�v����\�Ϻ��sKF�|RԂ��gy�9�d�-�� ���/k��ַd�7�x��o��_�j��d�W����E��
���N1��29����g�AAD���Ã�e�ch�M���}~�EH�,0�&]g�����.%����S�#
��`,���O=~��1��{��x2�P:���d�}_�2�@�%Ʌ���\.���0�E���Zk��h^("I�H��R�hF*$�� �0 ���%�Æ�2kii���X*�66W���4�� ��0��O:II�D�ϯY��g�m�����U�B���v]�i�&ovl�"A3#�(�٨�2��ώ�9����H�k��H��.��$|��4D��ժ��O�/]�f�pM�}BӠ_:������dv��r���s+u2 x�dкe������LjS��]� C��G�<��X+$p��Q���3
eZ?T��P�a�c9��+�4h�3�')+�p��}��}�ҕ/ⵎz酋W<p������S�/���[��ac���vww�}���LMM@���{6�|hc�y8�	OS_Ԧ0����P�Eh A�Yޔ��:�a�GD%K�	�J TQ4�&�����(۶5%�ONE��'֮���oڼ����&s�T�vE��2�~q�G�9��p6��ٌ��s�������x�2?�P�6D��٧�]��9�2:l�ܲ��o�X.߷h͢�^x�e4�[�#7��-K�m��tH�AQ�#1	p�N��'�@�����1Xй $EdŊ�|�Rdb����pMj�ȁI�RsS���8j�9�Q9��g^��ݷ�><�xrQ�<9Mhf�Ν';_z���i��)�R��6%��
J�w�z�8X�����eT\�H�&z%T@�q�"��S�F�� �H@��>f�y�hDԨ>4-��.�H�|�0�Aҙ<>vʙ���[�3,�c������+7n��M��p� ������_�N���~J�J)�]�]$����8���-����ѧGl�N�	���]�D�?���&���4Z�qE���M$����_:���w���{���s�;��SA��D�ӅRi���~��8N�����n�I�@�/�HH6ہ�w�>3S�
�a#p�AC��ń0�1(�� #� �Bu?<��6*"h��E��j+ʟ����\��^��A.B���'�ɡ���o^iK��~�P�w�C!Vc " ��>�L@Mln�˭ԙ��N���x<Q'[ӣr�� u'P������ĺ�uk��0������/���!5>	c�	6�Avl��f2�|�]�7ݷb��}<v�>R��/pm�v|dnA���$���4���}v����}�{�s����Z�A#��
������g��_��O�V�t�}nY��$���������WG�+�aގ׸�X)Gx�f$ctMAOE���&����$�pj���L��F��"�j�Z4/�cdd�Db�&���m�+��� e��OC��b�|�������{��'�x���i!��x|�?o��r���dV+��fYĀ�lt1�}Jcǭ�:�n��0� ��C
���P�4��-@��FU���ԕ�J*�Rg>��@���b&�'3�8�G��OK�Ɵ\�ڇ�ذa/�	\ B��b��/��UQ�Ÿ��0չ���i\��|�0_+#��}�
���p���9��z��Ӳ8|����/_��R&�7��ƽ��?���/�?�\.��oUl�Ƕ������u}Ӝ ���A[�\mD:�h�`늀:q ���P��10q}R���:l?���+
���,71>����[o�X���3y�.2���'L(��«o-޵g�g-��dF����#jVRn�t�΀X���x	$��&RBTkP*Uj�PA��u�P� *��p��B�Q�c���@<�V����A5m������L������cQ'�S����V�]��W]��kk�[. �T*M��}����-%��F�|�$���LN�s-8�-�sPd`�ɐ��5
q�k��}�e��[/����Ͽ���z׷�]�ƽ�0�瞓�!�t|X(j����V��m����"sr�E��"z��@��^$c�����N�\,�لSA�Xd!S�WY��͟���I~�����7����!�<"��K<p�	�#�tp��oo.
7�����<u @� d��V|\-�i����+V���:X� ��1��\4�:jԲ�4m�K<47ǡ��A[;�bq��,�k튙���ɦ���Qߓ��Z��5��G`��\@��W�W��ތ���i���y=�����>ϙ"���F�5�,j@i�:K�Q�o�*Y0-kQ[[�/[���w��g��o������!��}����&�|6{�e7���J��9�
�"E ��cP]��{&�P�Aj�h{<akZ�x��AVÌ�ҁ�nu]ר$�i:�j�r�;���{i/q����F<p�	����'oH��>�ƽ�D�� T63a&''Q�TXg�H<�|M�V(�6Q�6QXmA�'�FbD�ց���zOlZ#�O�<
���B[G7��M`sd�yM����
Eh��lY��D$��M׮�ﲵ�y5�d�Y�s�E���pB���H�4@i��fG�&�*��Ԩ7`y~b=�Ghm@ ��Ѹ/Y����֯\�F`�&�X�=�ޫ��W��;V�eW��7R'�cY>�vj  �Qv��Q��"}S���>�AD��b4�
	 ��a�^ai�bEeQ:�(Q<�Ʃ[�e�]'O���k������=�x������u�ݹ�NK7ע�
F#�!*����t��E��Ex��V�R�a�u�Z�H�RĀQ��CL���2P����h$B`��]��;�B��N���8��
��noMN�«�7���m�7�z{=`p��$\��`#��
H�d��"'���L���Ff���]�ـ�N��|��L��qjsl�e��m�T4C[�������d�A|Q�"P�׻� UFR#i��Ԫ��f��t��CAF�L�H��zQp��=�``����E��em��P B�{����a�� K����_"~C��ܿ�-;w�<���O.
���E.�������۹��1R��i,ɼ�B����8��b$��*�Uu�!�1r�A1~EfǓ¢��Xl<3!�4*�dS,��d[Xhr�*L�O���(��+����Ӂ����W^z�m7l9�y�V���,d���ك��B|��%}p.sf�	ӄD��5��X�_��.]��x�� Fm^�k���S�Y�v]*;�����zz�����`��U��\�\wk�Q���C�����X.A<�L.�
y��,1�O>Z����l��a$ _�LS�ӽ2�S��~��'�߸{�;�⵶����/8����|��5�_(�*=�H\�P#)�b����&i��T�:���F��jh�r�B �ʶ7�X�b0~�<]ţ�!Ԯ����NT�2SB�Ccp��10�\`N�-YhN�__���t�U�r���.���T+�-�^��w�S��e;	|6�����F~v��iE�g�7��쀘}��=�vl���kk��G�����N��65ⷬhZO4�}��i�7o?3�'�{��;��|��G�c��թlzm�ZI�M��!���>��4BA?�߂�����6=��h�u�Ba
j���,������j@ׯ���;x�Э�{�0��8xr��.by��񣇏܄�be�P�����R��j�qMU�ӊ��>M\����AY�QkPm��J'Ќ��� &�T��Z���Z�;�tyTZ6�� �ɳ��9���5�\�a�C뮾��Doo<����zQ&<	�v���v;����m�L7Լo�L�s��M3��Di��g��L3�Ck�~T���d�i�W\:|�=�<٨? ���V���_������ş��|[&ғm�y),��Z$�N���:��#pN�F�\_����V�&���L���S��H:�'�����~͞=�_���y�H�x��"��I7�m�Ϯ���܈ʸ��|f�яQ�(����X�Ljdݨ�\���L��Q#g���~{1�N`yU�*�h��$tu�@K["1��x/Sp�����A΍E�Z4ܹf�ʟ^u�u/���UI_$�ϒ���x�)��6i��e�u�h8y�FV<s*c�)q�9>��3�Yy��@��b:-�@��?fl�hm�h�kJe�B��>��/X�����V�!x�{�'�����w����������x2���X.���C�0G ��,�E�y��<[�D�������>�@��
"X�׹%Z�d�~�UuAŒ��]�oߚ=x+#��-8��ڡ�}���C��"X�޼H�����A�R	�Ji�WS/2`@��6�̈́F�4E
(bШ3�Bc�"G�	G#�����e
A�R�t6'O�bʀk[��ζ�=���f��g=`p�	U��s3����"��W�9[L��z���%|\l� ��{��9SsF��S&�v8\[a�u�^��?��������H��:v���屩��߶>���J��j~���&JP+$����"(�+�u/� ��Y:�R�D�D�Ih][��e���ٿ�5����|�x��"��å��{��5c.�p0�D�c�~
A�"�0c0T3���h[U���R.�|�sD�BdITo@�	)�1R�x1����4�)�hbۨUqphғc��ez8�;ҳ���n�ܯ��Y�O.J��N���/u�C�ao�m��W��D���u�҇�3q
�)}Ј ������������'S�N�h�iS(���+W������?����N���v���hJ5,�N<�
�>CӸ(�M215R:!
2�NM��b���t�"E��e\��
�-1`/ID-R4�88�o�[{�Sk�7���\dB��G}y��x�:�r��Ѱ�
�k�z���F�t�U�5�Ivd�x"^�1�HWP�1@0#7�����:ēͬ8�fΧ&�a|t*�3x�Z�t�/���ǖ�Y>�)��[�)�cN�y��c�����D�Y� ?��~��C�=O��s��3�G�=�ZS�'�2�Cl��L��jnn���V��;�y��f_���sx۱�,ٱ���/�spX�O�1(6~W�"�.s �>�k��e�N#x�8����KjcV8��bS����|}êeD���'�x��"���x�V�v�E�O��"�Z�>�M\��D26��7ڜ�
�Z%}���G*b���(�@�eO+���������c�ɤs08x��YU�2�c7�4M.ho~���nxl�-cޠOH�9��q��+��n�F�q�qsdf�����������\���B�4�3	�Y� �OT/@��8�h�W�/��j1_��$H�)ĉ��S~���}��`×}��|>r��h}A`�fԒ^4Y��u.�Cl�#��@�B�MsX7ݫ$ɬ8�49ɲ쾣G�^y���Nܗ�@��)8��2���O�����I�V_( �B�уC/~r������A ��+�j �,IQ��d��E`U��^F-g�͘�H_J<��l.聖�%ӆ�L��� �� ��N��/�77�yӍ7�r�u��X�<�)\WA�Sp���� ���bͣ=�Q�0̉g;v���4�s� �y�s ��O��7y���S
���#���X��X�yu��e��t��k�̔������#��p�L�G���T��bl�a�:�cZ�t]E������bȌ=C<�d����"	�H�O��o:v<5�Z��Ё�������O.8���E$��ڷ�З|��� 9�શ�X�B��A�P�JYC���Kl���|�R��*h�Z��T��A����1�5���Q[:.~& r��`ɢHDc �2;��T����\Ƀ���D$\Y����-�7�|�ƍoyEN��%�x<_*�^��#��z3n�EP�3/E��1��ϔ�=���5�[��l�i�M��cp2�a.6G*44�VP����D��r�9��f�ڕ��K��Z��\޺����l�[_�ֶ�����T*_�Kj%�߃#zR��|���@�AH�lSkS3s�&��JF�e��8����4�\�W�ڱw�ƵW���f��N<pp���'�\[�T6����ēWb�v�b� ���?R+#�?Efu�Rqzv���eI�h��/���;/��B��8�rF7�0�6���	T:UW���2�P$�h!Eٽv͚�ؼ��6o¢'�H8���rO�����V4xm"��9�y&/�\230�K=�|����1��\ a�m4����MBzr�#��|i����������������Z���w���]�l6�DC�����*�*�"�&7R��-���a!���i��e<	��@N��k��O�gE�e0t=1��^ut���x�w��N<pp�ȑ#C�ǎ���N ^	(l@R�R�tf��M��"�4� $@�U(�Ҍ^/�`�&�qHě�@m�o1�7J%�V��mmn���E �B`	��eH��T:���ۖIď�߰�W��ly�g��"x��Y$���r�G-Co�l�N�\����?�y�}g��G~���G�4�gjc<S-B�wJ�Qka4�Ы_�`A�W7�Y7���qbM<���}�������>�X��o��F�kP��W���>$ޒ`@�D,�
"���^�J��E?�`�ڝ�3|Dشw׾��}��)҅&8�����]���*\�A��Q��&.NA6�� /�,�w�O��7Q-�U�7p���7A��`$^DH��Mg�Mֹ�;6�)<�l�Ύnhj���t.'��app ABױ����W�z�n���{�/��
=9�焼�}����.nZ�/��c�
�������T8Wn�����T8[���1ä�9��W����t�UW�G p�N/0��a�9�:�d&�D�4�U*�0�I�yf���>#���q$�)�8LӨ�%��@��
*Ky۵���z/w
<����P�#Cm'�q\��I
F���f�y�Nd���P�|
�$6��W�\.��?K�ȒZZ���$�!ϸ�yQ �4�	�XS$=����D% &'���*@�W��X(�_���7W_�����Wz��|����j����k��n��m[D��4�f`�ӽp��;���3y�s�\ �\j�įp��ęכy����:~��
�;	�x-�{������������뷧����玺��Ԉ��+W
�.򌟄:���X)�P�M���Ȓ�� ۟�e� 6� �@#�	4�,JW��%x��7��\��J����봪�֧(�uA�A�T�B�Ċ�C�����
��EHQ�#AH$��W���aS��e��l���A4���vX�`D�#���346�FF!�M��L��BeAg۞��|𺥽��O<�R'H�p�s�f.���}��:�Ϭ9��0�0wZ�!O:�Z���4����(�O��l�r}ꩬ�m6p������z�o��oK��Ͻ��S�_��S�cc��i�W�9@�^EС(~�wj���0Ȣ����L�	_�Im�Nmb#�Z��Ɂ-�N��3Ey����B^�\�?L_qq�H����͒��E!1��jԩh���<�s����� _��C���T���h�!�LBKK��(2��&z:�K�0���,vw�Cׂn�$�@?�/©�1HONA�Xpީ����j���nܼ�un�����#	�Jw�=��꣮�-��rn��}-B���C�QCP����\|3�f�|$K3�͸�y� x���Y��!d�	�7�T�`膄�/[���Ս�u%Ϟ |���������-�rR�c�}�J�J �-p�H�9�Tf�}rm�*E�〦�H!�
GX�hC��F'�&6�����x�i/=x���: ���
�2Ș
ZW?�;B-�#��T�,X���~W��l�?lC�B+]���������SCB�=��U]��v(���U+ h��0K9F��/�2Ќ}r�X��%Z[; �H��XT/�Z�,Ӭ�jM�	�����A�)	.�B��iH�M�Z*��ٞH\zɲǯ�j�k���2x��o!\W.�Jo������v�D#�Y����9�g�g�8Gc��9[�`."���X?p��s��H��0SĎq���ߚe���T,3�W��{��޼l��������km���s}닅��"P�;' P�=��5#�ԉ��ڧ{ � �tF6_�J�򒑁��'&�'��\0⁃߳�����鴢=�JT�d�L!��*q��'M����-�6���v�23�W%Y)�~Iw}����"������,��<H>��vnp�V�X,��Ɲ��L�C'��NB��Ate��-9���T̳9��Cs��A3�9P!%�T���1D����Z�Z�w�T������b!��E�\ڻ�śn�ԯ�m�0�y�|jeK��s�k-F`�D�لF����!���-%0��h��+g��W�����^\-����I�@uR����c������R�Bf�{ ��<�$����)���}�����Vz*���������Y4��
4��"�B�r���	Tt*j�����H��Ҵ�P�O��)5>����^�}��Ura�~OB<08�_ߑ�t��2]F9��d2]�i$�K*���Yn3(h�̛� ��8�iAr�k㚴]�'��ٶ����,t�q4N����@�T��b��o�h[I?%���7ѹ��a�T�P.�Y��Ԅ A�u�:�
D�"Q�m C�����Ĩ���м��d,Z���{ 
�ɋP(�܄	���X��"{t�~��M����ī3����6�q&�G4�(�p#��H}̴�s:g)N�����{NZ��{m�;ꛦ� � ���e4'���/[�"���~w�O�=�"� ����o�ɷ��w�@h���㉗������~4M��*G���9�4��:Y����(����NI�x|����>��o�x���\�̅O�x��w,�P�����魌�_ng3�����@[�璢�[m�l]�C��U@ϝc���4��Z�5�S��L�$�	 8MP���y�P�Qഊ
��B*�$���~�v�BZ��D)�<��<�i\3��h��!F9N��X�G�U0Ћ1��P�)���V�\�1�����0�
Y�b5��_����oڰa7����C{�
W������Ռk�J��g;�zڠ�v�8���CfF����BDԗ>�(�x�$�.�]5�����w�����=�af ��n�/��/��B�J��V��ţQ���@���H�� 5(U*�un�e��Ԝ�s�TSG[��G�.?�pE�{>�u!}���#��!�����>x��N*���[$iQ$nA��7
EAW+\��r��k�7&Ʋ�� ��\�B
��~��(l�&8GS9
E�$�")��)Q|�ӯџs�T�۶ E7�A�l�
�,*��ã�ީ���ˠ�K��
>T�,�18��Y���$,Z��1!�x�2�7�����bv
x�2c��ЪK�o��-o5��{u��N��/���W�
�l�c��i�!i�+���Ε��#��랉ifN�_�y��jUAmqɂ�fs�c����; ����m�Y%��ٵ�_��w�^X,��A�	 ��uK*&R-Rc���d�?
�'!��t�4�~v׎=���H�'�X����,�`$�J��~�p����e�f�t�E�:�7�ɂ^*sh�Y'�&H��%��@,r�#�m�I샄8�CgA�e�LW�*��8Q��)�i���s��	Tx����� Z,��ףN"9��v��@$�
�Z�&^��hCU����&����![5 �W��dNUKP@eQ�]��*@( ��n]m��U(��=f�%H��C)_ ь��ڒ�Go��<޵|y<��w(�`pJ0�'+���]�O�\� A`;gE2_t�\x>��¼��\������K3� ��� _�z��o�
��1�sh�)[�jo�s�0������|6�嶎��'�Զ�1��q �}G���C����zQJ!���CGE�|6'u�u�ڶ���ǟT�KݷdI��iO�_����$��0!s���#vmv�r�uI�\>߬�r��2}�؈�݀T�C�!�1��A�R��V��Z����f���B'�"�^���#�2�CbC4�s���}~_�� Cb�^�)퀨?dh"\*����e����I�8ԩSF�4�Q��aq4#����0Z)�`��F��g����牜�Ao��ZEud�϶&b/^��G7�x�0|�}_¨�נN�
*�?��w�-�)�q�]��C�=u���:f�͖���)jl\���!0R'�2��9��&I�5�W��fs���st��-xrtl�S��O�B�&Y�9��ܔF%�؈i�`�N�f��l;%3���>|�x`p``�����<x�|�`>:~��MՓ÷��?���1fb�Su*�&�
�휃�����l&34D�h����.H>ƅsM�r-�t8�uD�w�2��:�)�c���:�Ԓ���7DĀ$'#�/�G�)�(����Ѡ#p�����׈�#�ɘ ��(z 2�~A�1�!��^;��LT58�C�*�CQhW� ��0�ʂ4�'�P)V\0]-��۰vͯo����'|��1�U�;t�uׁs-��ܔzv|���ޠ��N���{�(��L�7]��@}4��i�;_(��������g�2���f�l�xW4|�Wl��ѣ�mjn�mźUS���/�,�l���������d��\,mQ��$��R�y@t�4���
�q@��؆���R�ѱ/��?pr`��#G���s������P�O�x��\|B�����{Go�������Q��Ld'3,4�+W�Vd0�>��t86>
�3iȠ���:t�]N�9��[�S���4LS3����5˲tt*
����\��*�"u$�D�����r\��*Z����k�U5���b,�I�G�a�JID�a�4CS8�|E��Bo D�������D���A;Y-C�A�E-���� 2��TGG@ql*M�jiy��n������V
{]7�ԛV����>]��54���NN���>�����MZA����4��Ն�q�Aם��p."��3z0� q����d8�����!�ce�"��|Q���뚕�����,v֡f��_������l����Z�e�c���P]�(�P
�����Rɦ(cn��c&�MWh�����T��w�|���*xo;��O�x��jO����̾��Z�Z�j_V�
�ǹ��@��n�	�ã0����Y�
"m׽�F�j�z_Sh�'L��>�Ғ��'�m��X"at�uV�[:�D���uI470��ʪˊ\W:�����x�ٴ��ˆ�Ǐ���d4Db8$U�:4� �b���P�t"P�����Bw46�/�0%\��2O�eH�E���8*�	�d�K�`�� ,4+�h���77�~�g���K�lI}���]7�o�|��G_��5�t�&�-�n���x���tg������=���V�y�/���3hԞ/�
�</܍�u#Hrj�Bje�����f���~�/�a��i���3�{�}�-�@��3C&�ֺX/�l��;��,�()��e�vK��cMo��b�T��~��7��yۇ�o�m۶L����˥�%Yh-V����	T0M���(�P���T��ZMB$�rEgsW�UR�1Xڷ�;u�T��g���S/U�ᄊ������|D!`0�}����o��/��격S#r�sA� ͋�+v���b2��VX�tI�'*f�`"���ӽ�Poߢ��}���:{��ŉ
�'��U<��$Yg>cK�t�Ĥ�Գ��P?�i�2��e0��90U�H��Pp�@p�*�������.�B� ��d�ij�a���]������ ��%���XZ���tZ;V�����7n\��*�[1}>�ۮ��O?x�7��I��_�H�`�v�1����|�N��?��s��C���ˁ'��������^��,���V��7�-�q��#a.΄9�a�����:�<������+<j�'p��.Y\t~7;�wں�������*Y���&Ƴ�@��4>�rL����� �HL*R�#�x�|���_x9�h��п�'=�x��>���d^�~9�ܵ��>�fK]'�U�*��+O�����F�Df��\M�ɧ�~�o\ժ��F��%oܲ��S+�-+\r��o�e��;9t�nۋMTS��6��@7������	6T�vs�R$�8��
yہ	W�}#�aqs+����&����!e2�C4� �J�yH��Бl��C]q����p��tho�>I����_�B���/���#�_�}�|4���U�4����aqJ �ߪ������S����m��Nz����z����ﳵ����Ġ��-2+��@r�	���ؘ��5���#�a�󁂙�j��Q��s:ǻD#ݒL�o����_��߽�;�ϡ� ������-��[�q' EuUQd�jEec��e����-d�YF�D���ʍ���B��"������Jv<���T�'@<p�!�Z�Ww\b���P�Bq<�z��q�۞2\((~�}�0�YE.f���A���T<{���7�^w���>��S�^{m��2&T��k���U}E$����,߁X�'�Di��#`(䋀 I��E��۠.K����JT��)8V�CW:}�&	qh��!" �@ �錆	FހD$Dߦ)����j������z�nwhh,(��!E*<��`�����z�p޺�O�,E���͙F��D�4;��?�Oq��%���G�����/���x�xr�H=��^�G��r�iZ�+��&8�W,���٬���5�h�i���ps��L���<3�;�=~ �p�ŷŢ�Ou�v������s�?�łc򄴏�"��\�u%�R2T�H���3p@у`}�#�BF�`���QI��%'��藏?2y�u�^�w>��Bȫ���u���S��eN��V�9��E�H�6�=��8(�ڢ��5�(�w�H�ŵ7�}���ĪU���o�?42��p�E6��B4��� 8�4�U�Ё��k,�`�,j���.��Z�S�0LUr0�V �@р�.H��0��Á\�X�h���fh�x�8�'�b��u�/��I��L�ck�=z�`b�7ZV�|�ݳgZZr��^=�<�m�~���W��������[�|�۟���B�='V���M�J�uq���������K���]���_�ێ�~����>ߤ䃻���Sӛ��]��<.��ʧ��0���I_̪>����5}���MhDj�YSf�`�}�'���`/m����f؃۶m{w�֭�fK�g"���L6}=�h�Rb�X�#zQڀ:��
)z�G�L���B�kaɒ%,�@���q?~~��];�������y��x����+�����wS�t��tb��8>!�ШZ�(Lh:l:	�:o��O.�B9���W����|��o�����Ï����S�����"*-�{UWY��P��M��D�\��D/#�C�����+A	G � ��;�'��&�a�E	x�W�a�d�|���DBvoD1:�>=.ܠ�"����l3( �v�v\s�ĩ���o^�bWSߒ]����ѡ~���(k�,�ߖ���g�>����?�͊�y�����$e`���u�;���S���s�,Ǧ�RȨ�?�,�P����?�o;8����Y�伐z�b.$�_S�k��*�~��g�Noml�>W���ƾsdZ<���>��{����,���j�l�O�.���  JҺ�֦���������\�\-�Ǝ�r��h�� ��d��b���"/Tc�`x%�@��$�Ρt�za�(�a�̪����_����k�y��<���U<pp�����{7*��]f*ݗ>%-��07
�}�$L�ɭJ`(�@�.ko���'�����7n�<έX�;�Q;�+����Tmy ��ɦ҉�X�Jm�҂�^hZ�\f4�===����tr�h��Nq�\�cҙ��!��� Gb��WpT���Vt�p�����%��m*��Ŵ�[$�5�q�0zfA�!��.f�m���uC'�n<Ւx�m��W��_ީ,_���V�\#	�]���D��v��T�����G�ٰc�X`gnl���}_�Z���4.f���x;�FE�sEjW@P ��@%�Z��ج�2n�R���a����<��X�/�p�H�� ����:-�n���8�y�ȏ�ܙ�~3y��l�g\��}3��| d��2�z��Q�Y5��s9��l�hmz�駟����9��;�t�:q*��0tc��V}8�pl8��sRĀ"lH:�c(�P*Ո��G�D�D��P($�?��cOO��]^!�y*88���'��0��br��+<��vux��!H�&p��kf�X)<��[n~��_�➦��*��C����T^����<��!(���c H
踽��>�²K��TU�P)�
���l�$Ƞ
t�����0+2
F� ��@�)	&y����v�
��.:�����}�m�_�ͥ;v\P��IA�
��'
\De�q�R��C�%SS��Gv��\v�W�{��dNB"Q��oEi���u�ᾩb���~_.g��sOr܇�D��`�#�_i�w]]��x�yI@�H2A�9�'Fu��`�f�)x �)�aT����
�}EJ��3�ડ����~� @���0�$�=���CUW_�k�:��\6-0�sg��\DL3S	����f�<�^f�u9q¢X<��j���<����=�ܓ��G���FCO������=�t����C{k[���t]�$p�cC� �x6�$������<1>66�R�oA��w'88�����zK���Zu8t�H���a�z;�' eih\S��a�R���o��C�o�+/95�)��SS�y��`Kd_=�L�Ɇ6�Z-��S$X�d13��ã`p�Kr��� 4���6�а�`��z-�H&����D�/�����m�������Ӿo�����o�z}��;��2�ɭ�f_���bR@�aaS"�j����.��|�w�ܿg��+�_��W$E�P�n�M��e�����K/��VUW)��(��?��܃��S��'���|ĝ�����>;^���R���sL��ī�zxT�:����0��Έ���5�DAϔ!2�q�\~�h˾���m�/+����8���|�w�R������d��/��`8-\��Y��:�.�ɠ��~�(�\��߾��4�9�sL�j��ԂB^���p8��:J�ⱷ���Ŭ1��L���Mu��p0�
e>����M��B}B ��4�:u
t�X
����c)�l<������_y�-jo��y��x����ӫ#��-�щ�a�4�9	�h%��� �LX�l�駾�����a���ǟ���[�jy�O���@T�"�u�J�1�ybXF�g#����fV� �(���&�(.���$l\��x��}p/��9(P8]p����Hi||R�tuw���G�>�-�������Z�^=�{��{�ygga��G�}���T��ɩ����pG�T	E^�q���ȭ��Ė��SK^���l^v�5O��^�:~�A��P��C���t�ftA���>^����x�[t]�A��MN����������N��|��w��{�p��6;��`��W���v�ABԉ�Q1�+0���O�g�e6�ҭW���w�����JI�E���?��G��/�^�y#�l��_Sl_��[qĘ�ȣ%c�0�q�?s�ځ�j��?�������t�!����#�@�u�J�]��]U�*�쳝7�Jّ@x@���,Ӿ²,?�P�"�Z�W���E*I��M��e2�d��i`l����¸~7��������c��@�G⁃y�E�N4����剌@�"o�p�*¾�a�d�Vdq���������7?���[��$��'Ƨ:���B�R�S�3�r�,��
ˣ�a�1P�]v�%
`rlD�ExT"��򈊬@��	Z;; ����Y	C��
�CHe�\�1撅��¥}Rz2��Z�����/�y:_������|�[�����u���:�=?tr���}k�lq}�^�jZ<&ۜ9�
$���H����O����w��{޷l�A��#�	X�����/˂�ϻ��Upm���r[�\�Y�������Ó/;�,Y�A���O�S>i�dI�a��T�M�v "��f�
L\)�������CŇ���9Vg�r�5�4S���do�LV�o�������+-v4������ێ���K1�?�m����Jfe�~�1[8"�6��HA���AM��`J����X����B�t��Xxv4���2>�\�T)�U���,B����	*��j.kf�ZQ7g�TxH���L��wPf�H~���A�����պ�B�dE"=#T�Z{������/o�F��-�'�x�`~���2.Wޘ�ٶ��u����M�����E%ը�Z���m��ڷqK��~�c� �R��xA�@�A"�ި$�\ UXЫX�$-Z}��`�CǊ�X��.qP��8$[[ ��&�e�<3E"�3y�:r�Df��-�{Z����q��CG����_��Yy�=�[�����ԉ��_K����c;w\U��QYuG%)$�ʜ���Um�ˏ5�5���il�ž붼���f���Fx?)l�w��^����*���$b�-�߷h��.:#�o>ֵ�� ��s�N��Ez���h���#�r���B���]r�᧿�$�A�`���j�X�@��ש{����� ,��AF���銠��%cj�����,?� ��!u���i�
�g�������f)"�M;lD>��!�smM�-�����R��'یѭ��qO$h�U���UU@o��tT �k�D|�P,L��d�
��6tM�Ћ�ST����L۩��������G*ޥ��^�u��:|��z��cx��x��x�`>	[c�˝���R&+q� Ղ�,LK�hk3}����}�Ͼ�kɒ%���"�B:1:6q�OQ�iq� ���@� -fT��`��ِ�|�P=*�g���$�!%"�8$�[!��������+~(�(�8�a�ڟ�������_3�M�p���ݭ�2uc����M��W���w����rZ=dH���:��o�f���:�gύ�\e�5K	��b"�o�����C�����������o���3ӓ��A� B`�Hʢ	�"�`9�-�Z���s��1�~k��W�r���-�J$DS")fR ID"��A���9T��{�����1 �S��h��UU����M�]��?N4���nX1�%L�@߅G�������oV�*�NB�͘��8p������L��:rp��у����hy�T�<Q�-0=���B�j��9 (� k]��1��@
���I�A �}��x.
kԔ��7�hWk���鑻���2+��=�ih��>(��U�]�J�	C3�p,eI��ǆ����ٌ� g�η�>ּg?��LdAh ���@Y`�˵Q��k׮=/��W��U�o��oO�>X� J"���H�� �&2$+�7�k�$	���'m��5fX�V)s,���*Si#�%=����w���#������GMp��F�>G,V��d�)��:.��]�# Ɉ���[�e'_�r�G^���۪c���SF�X��LE+h���*�:*q�7����nªuk�F��β�M�4,<��L�������-����d'�0�˱}��ʋ��t���׮���^�'V^�a�_�׿�m۾���.�j@����񞺡������B�_Qн& ���N�o���_��ͽ/<�{t��O΍��Դj�$�I��u�_���_ꪱA��$N�u�A����lI��E�@�18��a9����Z.���&���xz����D���xC����KV�xzj<<Af��r3DQe����I�;�T���[d.g�V�c?�/ro^P��5,U�������/�u?������יm�X?#yQ_-q.~�m���-������¯������<�L��HS�Dߎ[�*��q�뎎�����Q52�k�*�����=%3����� ��;�y�I@�μtoj4�������v��ͯ��w׮]�Y��I��!Mp������K�|e�W�GeE��i8Z��2.���>��ĝ������'/�����Te.'���-��M�֠P.A�V���zڠ�/A+��hi�BCE���<�a?�X��:���7s�Y�0=�'��5��[��#�=����G�u�xl��=����Nly��ϬYs�ꖞ����h_<��[���������ǟl$Bϋ��ao߾�/�|���+;^����+���+�e�Z�xkW��n�z�ˀ:���O����ȑX� UT4�oCm����m;��~�iZ.�o��[�(z�57p��\�o��}�Y8�;v��Tm.��B�/#p |��$H�s\�!�9�B ,�3��*9�)m8?>�x6�[�����[WϞ����?����}? �i��\���YaSM���~��[����NN�e����}�_e�fL�\ߓ@����(W��e�QJb>�uכ�'�N#8(��h'bX��JJ$C�ޣ�&KJ�(�V���T*�r(��mbD	��\����8t����<�ӧ
ccޓ=�bYrs���	�i�RڭV�Њ�����DL�§��fڼ�9��S��>z����o�(q�#G<����+�r��F�a���ێ�6���+ AX�Y5|�4}b$ү$L(ϊ6zk[�Z�8��y�M��s�����1�`޼�/_��W\���ꪕ�^x������7��ŭZ��E�8}�TKgO��<��?���u���׆���g)"��9���:>r�%�ݵ�kk�2)Z(Wd�"�ĀC@cZs�;8qM3 �Q�L�$F�R�b '�\�ZH�S鶎4�{kt��aI7X�I8�m3��;��/|�q�a��("4K�Y�J��g��������3���Z�2�K	|��7e�S�Xh�B�i�D����ޡla�ο��������,qP^~G�Q�Ǧi�CppZ�2):��ϥ�i߸���R�����N#l,I��~��L��*z��[��:g�3����'��Gϋ4L�#�N
<����g�Hj��q�U4Y��'Bp@!K� �{5�*�h.T�@�4�8�a�Dр)�\&�V�5][8zz��m۞;���ϽG���xo�	�1X�¾��v���X�%T:��G�Y��Dh��rt�v*Sv}�k�.�p�D*��bqy,���䊌�@���T́m�,�0��
�V,�{� �+�1n��Ъf=�qҙ$������*�ɩL�N�Q�@�\��c+V.}nن�o+˻���-[>����T�{���/['r���G���Hr���������]e���7b<,;���>O��ǖ����n��u���EI�~�]�%*\ʻ"��|WN�1�)�U�����p��X�h1�t�ph�~^5(����P��C���%���������0d2�P�T��h���dy�c���x^�>\԰��s�7�i�麮�VG)� y�@`���"^��T1���1��_�����=���F����|�U/�m�����r�N^���-�I��3������� a�ѥѷ�C�*u���9�Y�^��3����>^7a��Tp�m�����c �
��f'Ƣ�!˴�i9m�gi-�����w�GF����g;�#ѥb[�ƙ"
~oK
MR)5��,�&�3�0=����j�̺9����C1f��<n �M�ū^zu����9T�4��]�����/ϯ��ФH2�\�Z/C�5�u���M�<�pK�^��E٘m;��D�eG��*A�M$=Z��/f.�*� �s|=D�	E� �JB[W��4(�a�r�"8�RHǲP��y�������N	M6,�l޼����K/+��_���Prdd��s�+��޿��m�(ܞ'.�7zp4]��e8����o���%e�H���)J�%��]��jY�]��@�J]"�\��ST���F-��_u�(<�����I���- 1"��j�|n|��ÿ>�8��Ơ�c.�1�c� uv�E^ Y*V �$^�2 c%a��lN</A&;U- Y���IX�w�k-.^VO���{������6��G���Fs��h�J���t��D��R��vȀk A_�g�g2 ���h�}��9��N%���I�hM�y	D�\\o�C\!��{!��[ \�֋/��B���<��LW���)��u��$Ͱ !GX��r(A�r��+@�<��%)����*d2�Tj�8Y�B1��D*Q�7�����9�#�<�����틞��_4���>���\�P�X��¬k�d�g���?��2]sAR�R�f�p�ڱ�i��rI���U�+H@��@��~����a�ҥ�obG�cHX@�Nj��Vd��4��w���1J���Q9}�(��n�"h٪��Ss;)���{��'lӊ���u��u+�Z���XƲ��~���$-���O=]�u�������x,u�Q�[1���B�f��^��P��A���'eK#0�74 �}LH�F�Y7���K��Dbh��`�0-X=4|�]���<��6�.D{2 ���&��H���� J�E���� )	?�`��'%* 6O��J�u�O��O?~PT~����p��A�x���/�R�gF����-���x~�ip�;(���m뗍�S�+:�$�sR���ڢ�O����x}�<��EQ��b�����A��כ����B����I�r��\��8����2�C%�4���3�����(�J�ӣ�,,QM�_9�o��<��*���um��������~*o<��\���e'��V�V�ţ�5�9bD�����j�Q�%��=�,�hI3����ǻ$Qn��-�)B�𻥑P��J��� ޗ���YJwO�e:AVb05]���4��2���5
��=��_�s�ƍ�)��ᆏ�^}u�C<x�ݻ#+�-](�tF'�F[�[���O+񈔼��+pw{:��4αO�С��,� 3�	@�$	B0�LF�c�0�����T>�D��jLXb���"����$b	�Px��h,	�r^:x*"-�x"VA�I��g�3���%G��Œ0�|�$`B�g��,��3O��-���IJ��?^*~���^=�ǿ}?�{�j�"|�����x	�aTR���.��T�����Ϙ|�P�ab �_�7�>3��cv)�/�;=��g���TH?��Lrl.�D��o�%�x�������S=O�u�ĉ^#�X� E��~�qг!�@{��kĔ�C��g�����7�O�N����b,�@��ǽު���/m~��es'p
��a4��Y�6�yp$�i�@��+�hL\�h��T���M��ܺK����\y�y�1}h:Z���Ȳ�$�@��{
h�UQ�SY"�$��L�z���x�k�L`(�g:�{P���;66�|��8�4y�ٿ|٢W�5w���e�-�l��^7�]�v~y��P8��B>��{��?���}�S�\v�:I�[H���T�'Z� rp�<��fV���p��/~�įe
/ب�5H�#̓@J\�%^&cica��x,��0'���� ���_c�Q�z��mݐ��B���3D�(�d�H��
6��0F= �% ��11P!�|Ay�:8�d��J���xt���_�4]�w�@����˚L�ފ�r]�?2�����ރ39
��:�le/4N�N� <~��g���� $(
��!�S�=<Q\�C��u����r9gӿm:���/M�l!�(���$��Z ���g<��gs �A>?��Rggg Tv�����Q�r9¼�ý)��9S�ӟ��S��J���<����C4u��t������0V.��!��R2aqe��;w��E[�y�Rt��+K��ϊ�1���H!Zo�Ç2�I֡�����zL��L$Si��/�06:5��=<�kjәtj�����_�җ�/���=���Pya��{�+�?��ǿ|ņ+�eVEP�o���e˖�C��d�P���'A2>�B�~����b�1�M�5�"�g�p?A��]����yP(_M�t ��q�zd<~qO|⊵p��)͎�*)�B�#`��P
1��@�N�}PC�����qa?� `���ʖ������C�!��n��V��渨���yRN��l!ۍ_r
_�*av2 �3ig���x��s�&�:�>6�/a�A��� �x�FnQx�`��:}��.��	D�����x�V6l;��8�0�? �j��=h� K*{����Z[[X�p���%��z��(��!A�_�`Ep����=��{��4=jv4����[���^����F�s�2���������(�h�=w���Qo߾��]�Iֲeٱ݌��*�GIX8�M^*�DD������(��2�4���~�dZ�oN/H�(k���z����˰���嫖n�"3���BV��+~
��z���~�w~'y��o�4m+�(Wq&Լ�ի/���tX xļ�'^��~|�0X�4ǳ�/yEt���eR3A�U�2��;Vcm��2ȩ�G%�Yeг\�d>8������� ��R,Z:��ӱs"�JN~,�ߠ��3�8�,�#^2�Hxۖ����z�O�^�rl` ������ǽ�#F�H��}�։J���ܳ�o�9sޮ��)_��ɋ3����}B�?ԡ���zg�>��?I��9�݁��vuw+~���$����+�==G��)v~�e�\C��#�w���&L��}N��Lk
��3��*F��ِ`Tx��a�׽�ҋ�{z�Sh��{��&88�0E16Y����$ص�Pɤ��"�B������M��ȗ7mzp�M�_�8n��.t�y�3U�|�B�F�	 �P�Ş�8�/�Qi3�ݐx�,֗H�ٿK�LMM�����n/���{�,\��_�ڻ
�lܸ�y���Z���~�E�+V,���[o�V�N��謪�n$d���98A�Bx���O�#�B�<���������J,�@M^�0v}!Y)ט�£�6�T�e[�JAe�ǚ(y��d�[���0��b����I0�RJ���G��s��y��^�"k��(�I���<x3�H�;�51�V佋{�L4ݧ��.@�Z��E��q\{��=��s� �i�
�0����Ɉ��A�U?�E�=�3y:n���"�<:�/y.�T~u��ֺ�:� 8(��i�����0��צ�+�,�A	��gi?Ӿ����"(N�T���"~�����g
�aLN�>��Η(9q;�l�|�F �|�R	T��Ŏ�^�u������Zgv�8'OB��\Z4�;z��,p#��ֱ�Wrc���S�;v�r��ct�DZ��4m*bDQ��jV�@��k�e�uJ:�R&?[��v�o
3��*��PIu��YV���,���K����w���F��j�Y��]w�:��縸G�<?�
��ٍ�Ȓ�&��� �VO�(*$^�2Mj�@����P�콙�4~�,Y9�y|���1p�*�Kf�Q�E�p�,�|�|6~�����D.��>�,Gd�x�j��b4j"���$3�#`|J[��X/���눧!Q����NE=�j`�[���4Ǉj� �s���
%�^��&�����\����g{�.��p�3��=�����</6��<�p�����V�(�Z����ӷ�bv��ғ���;��x@�k���<�{�i�̀aB"���q��8��	�@���Eֵт��.8x� ��%E#p��[��� ��V�:	�OÊz��۱m�M/.XJ�F�9.���T:w��?�9�&��Ι��^~����5-z2?ͼ�	�*�(*)9��%W�h����N�T�T�r�����t��I�A�]�}K���ϟ���Y<�����=V"q�Ѣ-U�0>>ʒ/]��j�J���c���o��.��,�oѲ����]�����k"�\��k���������!��B�hp�L��K�*�[R�^e��8.����K�������cɀ�����nZ�CA�E�]�$�_<�.�S�߀�������렊����(�]j��H��ær-*���@�R΃c2*��!"'�(����%C�N-kZE�� B���ż^]�����$ߵ~�2�=·�p68�{�*��{����	���uC���W|�?MS�_FCbUGg�jhZ*�����_�Ahkoˊ7&	�M!;�'��g���>2L?\�@�c3� ]��F����������(�sR�c��Q<tMM�n�����h�<� �	�/����"D�'�WwvGn���jY*%"�--`��wq�-���(�k!����%1��j}zQk���0�ݟULӞ��|��8;mHڀK�,a���D��5�|� Bk*��$Z��{*�Fajr߯�O�tL�����j �v��6m�����ڜ�sow=�����s������z|�x~��� ����c��W$9�<J4�e�JTd� b(߽ʟe���u��|M��P�I<h�r'4�2�����jػ� ����H���"k��H*�bq0)�öX�Kʺ�A^Lg,C��D4�C:*�?�d~�Ei���7�����Q0��/���35���[:�-
��1��3=	���_A����P��{[j�ݘ�s��a> �3����9IܢE""�/�=�R���c����~�cm=mS�X�c{%��_�,���.��aGX�v�_�����gD4J	�T"L����Aͫ�ccz�)Ϊ������W>|��-[vPr��&a�?~���tO��"����Զ�F˱b�Pw|���ȥ=Gc��cOҵjW�6�r�Y�-�ag��S�O��GaB�T˟�eC�7����FN��Q��	h�9�&�jC�L�ZjmK�>o���~+j�M�n����j���N{G�'uCog�P�R�s�uviˮ<t\K�-���'�ì|Aj�x�X�AD0Ѩ�]��1^��H()��%^a�����S�!�o�OÊ�n���>���98���>�[�YR"�u\6g��<0e.�Ikx<(Z�ڐ�&�"�R��yq�7��������^7qm�L������F��� }�]�z f'��j��hx�]����>��	p��~?�������Q�Z���o����q ��szAQq�3��G&&'+��V� �H�(���]Z�W��&V!��(j GN��VѠ� 5D�L�"=cIȲ�k�/o�z��^����@�o<8��jS �^���U%ʒӈ��]�3!O��"
t1�eS��ֲ�UӢ ��EM��p]KB��x^�ի����Ƨ�^H ���FI#mRJD�qOJe��h[h�����遡%/�l[9�n����|G�#��%˖�O�]]��5;���V4�7`�Z�=��Ap����av�xhM�qѨ�Z*d!�J`]��Ae��L�x��\H���L:�BY�E�g@8	t� �	��\҉Z[�p嚅 ET����>��.��2��h5<FA!l{�'�TK���W�xn�/�:�>�!�rq�"��6��
/
�~����xj��x�����?pfE�L���G�B`0��C�%=����U4@��.\�r��s2��xD$\���4�E�?v�\��t�R���{����y�����'�N����%(g��pg��ע}ؚna�a����n`觼)
7��L�K!1je�so._�����ڋ��E�{����xp��rq��DB��ق��m��X�?;�0O�x��[������ާ�<���d�0Ҳ$�̢p=��O�r��u*�L����d2�B
�<Y��P�D�"XF�Ӵb5�J���w�Wo1�k����q[i]�r����U(��p�s��'��b*�*	�����T��0�� ���-����B�yP��#P"!$S. o��M*�������P�g�P�"��C�dѐ�'ׯgA�2�xrӧa�`'|�����R�!��@��p$O���D\Kxm�XId/̪���L��>D��:'�m!�Ns|�G:��t���^�W@ G�U��N���������-���]�0���A��0�r{� }.�8	���c��%ܛh0�r�B����i��5q����d[�mH<�4���{�	(��P�#�R���I�L�1���s/ޏ�0`��Qq��l��j#���/-߽{�G7�8��g��xw�	pģ�.b���%�Bqy�2�IkX&8�`��ENen2R4���W�jU���V�(^7E>z+ ա֬�T�m|��@����m8ڜx�`@=��\s�
�:us�מ���`w�Ȼ͡�F��a�"^W%.ar�g�9V��?w.Z3���Ჸ���rvFP8����a����B<�'A$s���E�\Ф�q��J�*uYD���e/`f�FJV�|	�9�3Jd��ֵ"Dc	(�X�d���;�����>?Q��DP���2P.�D�����6��{�g� �˵Բ�ņ����b���k=]��i\�m���ރ�pf���U3���r����xH�l`�ٌ�a5���a���e�)�p� �MDN�E�������0-�s%!{�ݝE�,�(;�yB�A��iޡ�"FXu�JE���7gDf@�����P
�ʍ�q/�0�4x]3�Q���3�؂��i�~��Mp�kRV�|�V��Z���瘈t�ik�2s9��-8TB2Z����f(o�E������'��M�L����k~�	r!R��6�QY��u�$D�^e���VhmK�A�gB9_�|v��V��,Z��]S�⹬|!7<::�/��(<���#�+ep�<��L&��d=q~��P �oy��g=�b�2ǐ�)����2���Q�!����17&	UV�����*N��l�b��	����)(���5��`�IK�χ��]On����
u�=���" �|�|?��\�Zi>�7G`����ޅ�Ҹ/ws�� .
\s'�1�aͶ:p�ލ/S��� �?�N6<�߮� �E��<|��^�X>�я��l��'��4�)��Ji��Ḑ�8��	��+�P��:墈�=���RI�go[�d,���
~6�88[�g�4G2X%�e���Й��F��U�4I7-<h�7*ޗ+�,Y��!�TK#�!��X�k�>��'�|}74K?���2�Xb���ަn@B� ���Yq��UXEE��~ZP�(K��y�j֔R�x!�
|�Rox)a��Y.���A�N��"y��@��~�0*I�@��soKED���H����T���vݩ9��[���8�v���a|��|Q<| �z��r�Z����l>��娺fz<;_�bRTe�?Ԑ�*��!���g;q���cU'3{�0<Vɠ��'D�SO�ٽS�Z
e�J4���V�Z"�oI%!�����G^���'
'�f���%Z���N���ET _�C������Ci� �2Z�	3� ��Q�������9�,O�Z��R���ZγNs\� �����]��u�&�I��oP#��# 3�0���z�g�L��%�R",�%J�&��Y����C��l�K��:���[X���K�A&�ƈ��b��G��AJ���AC]e)	PQ�F�w��I�H�.�D��}�$Z��Xde%��C��`��D"
����P��CT�｣j"�f�\�8Ν�7��O�,ta����0��ϥX�3�G�Q����Lݼz�k/�p$�{xA[[��}Mp�CV�%p������H��D��pC�N����]�<��ȷ�K�J%r��?��"d��L�a^2,�Z�� �В��Qs!f!����"���Z��RL��M.1	��y��N�����:�0���rʏV��*s��~ڱ͸Y�.�Me?S"I�m)O�8ʡ� ��y;�!�5ʙp� �
1"��<
�x��d��I ��(`|׬̈́S<�d������~.K������	��"�AMC.��H,�<-5G�s��m;a���%�[���@$���P(W@Rc,�󷉈*�@?k�kh�w�hc!�tRU�]����n�I}y���9����sp���f��o��=B�9�ǖ�4xf�*r��dyğ!��\KTD�Hu��'��'��G}-p��������������F��,��y��z� �i�/1|�
W�(f�%�;u�T�������B.?b�4X�눍РN�G!���<�4Si,a�=SB,�Il�i�
��HƤ�b�z�����o��}��un&����7�"{���꣞g�"���a��Ív��0���{�X�h3]�A29"ض���*~��6��n)��7��2�b��մZ�%̓T2�tZ�Q�^5���R������J4߻`ɒ7n|�d<�+Z��/]���𺋿�l_�t�\����׶F����X9a�-2p!��Z~�T�
�l�;�7�Ie?щ��$�hdO�DG<�2�B�>�;e�[����}Xf 	2�o�D��t
�xA׉����g^����a�Z��>�������g�ND��K2�F�$�>���,�@��r-�z��Ȃtbjj��C���Y��04K�~�F�����e;���!�^�if���a��E�]A.PX��7#cBD^�P�����v����Z�RA��(�TZ�`>�F"�Mf(����9��y3|	J�����ͅ������yG�kОi��P�x�@�	a	����е)T�3�Y	�ꐽL�òl��MMF%x��r<�.�|V�ύ�h
C4Gj��C���
��[���a͚�Zhz����h�����X���ʲ(�.�	G�e��|�4�\Gȗ
I�g��[}�"��A�%�� t�Qf=�H @��E�6��h�-m��ni�3�Q�SZ�R�i��3>��o&�y_7����	�M�6�P.�M�I^�GDDDqF*k�h<�#�� 2VP���ą�g��갋��C�$�/�=:O5����,rɛ4yldr�TT� ��o�h��L
�{ބ�7kPvy�ا>�~�i��8F?-q~Y��D@P#��.�f� q˳-0��0��t�{���>�����=�9�l��k28����	�i��"T�7�K!x�Xc���E��ẤP�0��i�2y2�!��R�����g�g?�#3�rdJڣ�#A�}�}��O��q���0yݘ�ޱ�F��;��M@��Dq����=�P�xLyv�`ww��ji�����ڞ_� 5 MX	VG�<IE�S,�.ʙ1<wN�k��z5���`�D��D�X�91�2����+�K��7>1���W_�R{�����h���jp������bD����a"ArL��Y5Ì�N,�j�bܦ��\�˲�����3n4�b�LC�d�v�,cCG���4��8��f �����1W,@�\FeY�V�<�<�b���ǎ���a�ƍU��9+!�|��R<!�̪wYH�~ӽ��?�������Oe���}2+ q�p"�z8�:��.Jiִ�qX��s@qZ�pE�'^�\���fhM��֏��i?�m7��l�Y��c���o�x�!H��A]3�9Q⤆�QTb]�K,����,.W��˾�gϼ�]>�����&��� 0���1\{�z���x��Hp��:�P�e���G<%�o��m^I��,b�dk%�={����?o���R	�ZR���KЍI��;`�ETe�Qt��ĴXx-�\�_��k%4�p�^��ߧ��|��ɉ�ķe����v�ܫۖLWӨ�1��グ��	(86pA����ʒiQ��E��������t!{C�\�����c���	�TF�t!J�T���j�񞢶i�ٽcץ��&n�f���8�� (F-���X\��;�|��ߧ'�h3E�~}���R�Vo��u�B̵Z-#����������R�3!A�$L���g���p���fs,ȱL�V)����\�h�_��bD�U�G6=�;��z�s�A�u����A�E��3��P� �' 8�Z Y��pY����z!ZWp�ʜ�\?�~w�.��Ƚ"vCĒȲ�eT�:�j��i��pǧ~��l�wN�:�=��q�g!_���ų��5���7�t ��٫�� �i���Q�
h���8�/_�}�����o�,�Bs�Z��{@,�/H�T��浆n�GU�jY��9�IUU_����X�.O������k}/H��:v�"-]�5�����c�=�u����*�\�֣�(����_����K.a!��>
^�Y1,�͗��Uf�Ŗ� �߿��X,ފrd}�R{�0�;}��Ŝ9̣��2�;U��&�) `0�sz,@w��A��(zϋD�B&�y5�i�*�R�������A���O.0�_f�Y'����MNM^�c�+;P���O�	p�$Y�F#e���x�%��"%�\�.�%��3��=����.�5_T�"n�R$�J�6#��PP#"p-^�i�5B���QI��Xy_���5�|Œ�?^�P�p����s�R~!��6Y�x�y�,��̈́�ȏ���f
^fﻬ������)	Vb��]�c>��ۨ�&����=��"��f�������,)�\�j���P��_��s O����&�YO�k���_����=������|m�E�$Ƀ�����2ǎT��,p�$����E����o�-�ȱ��\2�r�����O��� �_;~<�V*�����u=�k��>�>����U���Y5�]ύ���)\9�����R�nZ��?��'p�.F��B�/�upm�"c<ǽ����S��CCs?��e���+��`�!W_�>}�g�Y$� �}%�1�xK�b�~�p?A��PHI�h���['�Aމcǎѱ|kkkz"�*����.�{{�<Z[_�:�J%�h|��r��-=��=��/1"3|J�2ꆛJ��}�}�VK��F�އF�Й� �*�ȳ����d]X�Q��U�Q��,C�|Ƕ7�^�z�4��2������qc�q38���#8�c`+�km��E�'A3�Hy�&_��jZ��-㼘OO!�m!8�C�������̒�ǣ,.���5٦�IJ��\������ի���׿��{tw�U�/�B��L&}YowGG{��{��/̈]���:?��!65�a�\�|?��=�gU������}��?FDD�O
�8v�^���zf?���,Y��%HԄ���t��L1�d6\�
��8����1��?�;�}�ݐ�W��7�A����A���
ʹi��
��܅iVґ(�)/"�r\$�Yt�����T��M��={��x"� ����&!�����9�®7��'�ٸX���o?�y[9���u�w���6`��g&��������r���P�.�c�9��{V�E�v���W/�N���57\��-�/,9|��*~��?s��p��K!��Ҡ(��~
;�{!Lt�3���ku�hX���@y9�7���+��	��k_}����|)ߊ�]=S����r��y�aHf�J=��I�Ǹ�[���mo�NL��Z��.Cl(��0-��`�m8C�5?ŭWc�q�/d��NƇ�{�kdd��W��}����@��GMp ��#�EA�㦱Ia�c�����}�(gxhF�W����x������!(qCsZ݃$Z�Ĉ��-��P�$�X��Ss:2mK$!�ja}֫�)Ъ5r�;�z�Йi۵p���k@�`��U�֮��7wm�V���]���])�f��Lv0��t	�2U1P�3�, ��ޗ�-�D�ENd=L�p}�E�W6	$��$��ܰ�X؈	������B� ���Ie�ĔI�I�Z����h�8�ppK��̌,��o톧�����}N櫐=x�mA,��b� �Q��W���`}�<	��= ��@���b��Y���Ǟ|��.Y��E���?��z�%�8�N�Ēf&GF�]G'&��xc���Uj��[���}?iM.[m=�yO���w��� ��\��6�-�����^��T)˻��:�fO����]��	#GJ�B}s�pH�{���q3dal���dT�Rc�I��`H�jl丌O��Goo7��g��!@E�7t�3����聣�����MEʸ�M��a����������G��9aYE��(WJU���עJ<]���:5����^5*�;����1H[{�_I����i��H$�<8����]�w���+�4*��y4�P�M\��7����F�[�ψ߅�=�1�u�a�"�R還�:"�-�~>�_IA��@)._C�O%�Z�����b�D�khuƦ t��%+W�~�u�}�]3���l�|�����}�ͷ>:��1P(�Rm�(c.Ԩͫ���'� ͑�8s[B�<Ga��V�uu�Dg⧡s��f���T��.Da���O ��_�������:��|$�H��]3*�ݭ���� ��
�d���/Y��'G��4�Y�	��A\p!��Y84���Q|&iX�hȊ �� S�@N��@M�Rdلn>�����w�Ge~4W�1����	��t��0�hgM3���X�TU4�*����k�۲�l�����G񞧚 ��3ɜ=٬y8�Ec�$(<o�'���'�Z�
�j��yG_o_������L� VI�@�\f���jf#�O���IAG~����L�Ń�Ld���=m�������]ϣ��E��[t�ȑ�xn'�Jh�T��НR�Y��\��k�0����a�C����.�9.������s?rtxu4%�o�~!���t�9"�q?�A��P�Tɋ�])�oz�7^����xϣ	p�����J��v���Z�_�,�Y�5TȼQ�����u���m���Z~�x��!��M4�~y��Vhҩs� ����Ɉc�uI��\���=�M�6�''k+�����5�"u	�'Y�ɋEݯ�&��
�x"�<F��BC+mr,��84J��� F�L.T�f	�h��4��O�HB��l��ℰ-�O"��\W�B��m�T+�W/[٩l6������X}�e(U-dq�S"��\�K��-W��,��Ǟ�����7m �^����Pr8Zkh]ť/����r��S��WOW��$���B���`���jB,��J�>m/ѤPѬ�Y7������^���a�����_h�7��*~7���RɈ��׆˯�ߵ�(^!���2�#�?�P���H�3W>[b#�p�)��P�\� 0K���CL٪"j���Z-�ѵ��Q2��2 ,r�ɜ,	�"���D
��^uⱘ9aOS��)�P�O�����Qh�d�k�Cp�[-bn��м��}�r�W''&wi�J���V�YȐx�zZ3�l��R���Ճ�L2EB�ǲ#�V��}�ccc'zzz��6�q4��?\9�h5M��"�k~��: L
�6L��F܎$�t<�R(�/�DU*����R�h�9�X|��.	�ꎰ,d;UMGE\f�ױM���wv�m��|����Ad�&���l�R��V-�$�3���>.��BK"
ab���}ܝ��0��Ha��mk}�� �gʵx?��U4��,�Z�=�6ͳy�IOδ����7���tn*��d�
Gd�Q�W�f�S�VX�r%._'&s���xLO�x4��`�ܫ��A�����y�p��ص������5��u�U���/����H��j<G�X�%��T�(�u�3J�~�en�XA�B�ZCA�6�P��MZ㜖�j&���>u~�p���{���9��xu���	3\�����q�*cN�BC�q��ߒ����Ѡ�
�U�o��=�Lf�����lm�ry������T,��b9��4L"��R)o||����W�?�����DItf�/f���`	����~%t��kG��?J9��`�F�[�~k,�nyV��+p^q���{@@�-t��q��v�Q���X�5���T�	^ʓ��o�e��qh��4���."��ӯ1�h�$as�%�jn�.�<G����R+#\��tRk�W#_*�j�ì�g؈�ⓩx��Q)Y)�fH��+���f�y�w��]Uu��ؿ�r����Y�z�����W�-?eKgU�u��2-�DP#3աaX��K@��Zk#x`�ܯ/�8�Ne�ތ�/���% ��>���6@�S���X�5F�X�@k2Z0[��٩	hoo����C��K���	�"�p��$��;Q)�����S���.�/�����*<��S�)�6w��+a��!X��_���pߣO����;�:$P���;t��e -�p�gn�����_���HT�DT@0O�1_�5�.�W�=5��Z��X���{@r������M���t;��U�7-�\���Ћ�����t���	T�5
j�
����ַ�������>���n�K�HШK)�����G� ^I��z�^�G����֬��K��1�(�=3�YA�-�d�$j�,��� �Ȟ�(�h�]������˽��^�T˝�d2](�8����l�QCS��X,2���.P��b֥۶�vj��vtp��7}4��?<܀\������Zᙺ`�����fՒK��|n�FF()�%҈z�8Q����sjmͰ�9u�鬦���sH&bl�4�z]gT��
D�Gd�Ȳ%�G��Ē��w�Ks���o��}��k7?6ܡW+����q�L��B���9=�nia�!4�c�5�B$D]�h�9V7�@�g�`���˒�B
��mI��,����6���f���� B��� A�!�� vF���N��ɓ��S$�B� 2^{�[!=w9l�sߺ꜈ ��T��Cù�������!?��x�@^A�o�a�ͲeK`��^H�g�x�-P�Y���$
�hV� ;��k_���L���'_�����`��S�H�B��,�A�Eϊ:��ӓ-1>���������/{�����q��A�¤���ZPQ�R��ə�X�TV!h��2G��~{�1�쳔��y�f�������F�g�h 1��LO1��9������y�^Z�zu�a�b1�5�3_&����l��#A�����e��X�I�j��t��yjj�#�h4Q�u�����d�0��A�@�hP.�Y����䡦���SW�>�:�tn�ټ���p�X��zn�Cu�aROX��yv�]�<�>x g� �s��R�@�����H1=ڐT�Dɑ>���DsL Ҧ�B�D��6V�Zw]�.���h��� 6н��+zޡ����8p�dv�S���+/]W_��#�pT�BGK���EOD0�+��H��@�� ,o��L(����#Qj" t,�Jxܬ<��6����=��F�k،!Q�b��ʺ
"Χ-��T{t�w�����7���3���h� >�2��yp4���-�;��8�~k;ز>�߂�y����_���NZ���'Ylv@Ea\�������w��!�̃SA��zh��|�o�衝pj�N�3g�1F��=ᛛ6�ީ		V���X��X���`�9�j��w"{���R۝��4zj
����+8U�9C�L�W��n� 4rdVj���ݻ�g��0�ر�g-D0����!�v�&'���[�b��`��YM�f��L��ቋ�ㅾ�~�_��"�
o������9���g�B����c�.8b��6�E�v�T��ַ�c���c����2m��Rmʕ"Bk���m��K��K^�e������U����޷f��� 
�f���Mp�/�˞��j��D�:�Q�.1� �A��;32�� �NF�+R�VNh���?ψ�2Hs&w:�3F�P�<�����]R�xhkka���Ҕ�W����(��-7���}
Z�޷�����_�V奛ͺ����|�X�-_	m��K�"$SQ���M~j��z�k�h�P��A83�d�vA�)�N@��Y����;ҝ=O��C 4B	Lԗ.Q8��I(Q��$%v�ӌx&k��y-p�����ex��0YwQ/'��w(HFDa� T���ptI��O���N(������]&@��x�g`ǖ�೟��(L�K0���]�����`,;	C]m𕍷��m[�Ň7���X�-���0L����ɏß���w���((	-@����xA��x{���������=w���DӃ��cY�Q��u�
�aw���a� ����B�ྲe��ԓ�p�#�B4�ۛK���Q�����O�Sс�~�:�2�X,����1R$"��-��Z��T�SkI�P5	C$A���"�b�X�2�23���LAP?a�k$%2&�Yc�O6:����t2�j�R�VW�����	"��0`�
A���L�1�7��U@�L���j��##��Ǝm�Ӟ��xW�	���=R�D>o�+
QƁC~X��u#��!�ۋ�$n0��C�\�W�Ǉ�z�N��Y�u[��zM�c� 	�[,y���<D�oy��R�#q��W _(�nT@�,I��+/;���}���>�������mG��^4^u���ŋ/#?���+��`��(�x�����e���gO�!*ys���P���k�	\�\��N� ��?@pʳ�6�A������ɥ�i�*���Щ=^c��IH�3��@�t��g@`�.��S9��ӯB��QZ�ʪA�y�N����V��Go�m���T��8��,Z�.�{w�{�d	�[_ۆ�����?{lݻ��Sp���p�՗���^���R���=
�>�4pr�wu�5:���J�5:'�%0��M`�a��t��(�r_Wߢ��J�{�G���l&)~x傔��Q��j��j�s�g�h��.��kٶ,�4���<U~�c�a�Sm�(���Z��c��~�Z�sw}>���'ɪ�jtX(<&7��G���?)�z�yGy\�e��єk�jĄS����y�J�"��A:��r����=�#UE�)�`�5/�H2�,��5K�{"�3P�tB*��m���َ9�&ג��p�v�X��b���mo�^e�E--�x^����~N�����}`Ǌ�;��@�	�	��hYQ2��h),�NbAS�TaS� ��sD�4'�����^Ψ(W�D�jZL�S����
�ȏ\�d	�d=P#�� e�u���lC�u�������ƍ�kb�?����#W�~��O���S��(t�G�a݂x}�v��",_:?ȈF-L$�y=��q��+U�!��<�\����/e�8։6�Y]����߳�3çF6��A腾�H,&
���D�z=qZT_O���<Ԕ�1<=�t!� B`߃mNC*����0,EK����`��.hO��e�R�җ� >�8�:	V�Y�t�f��O~�� $;;�T� _�/���#���O���9�񫮂C;�Bu�4|�w�O?�(ģ*�?|~�OBw&G�O�箻>�����}�9|�@+���jZ�q����Q���K�85����ѣ
|~��M�������9Z�C�V�ɲ�%�.�-i�3>�FݬT��S���-[�?;�����W��)��b�T2;{��k��ƻr�՝CCCh�{\�T|ϛ�
�	]J�Fy��b�$�Bǖ��>�'_I'���h����O���0����h�cM�XY1/�X���
�"܇.+�~Ϛ;#����ֽ��{"�μ^�i�TYY�s(a����=�� @�3����Z�V@�dV2I��Z}ᑃ�W%�A�����MNVuI˨<mO������d�,�D�!뀍L�3U�>�r�x<�!hq��:+3"�1��{4M�������P<��X)�_���¶��=��{���:�߷x�	��o�%Y���N$�=�a��&]�A�E�����_@:y3�Zo������A
7uը07'��M�qlL����T��r��g�=��*�t��:�r��9K$!@B����ܹs����3�޷�]��{g<�1&'��A �(����V�su�t�T:o￪���6s��մ����	���������S�6Q8X�|����	�~�������1�P��(,�d�}T2�6;�{���#�4���zz�6{\տ��k��?N�Ӝ`%=�i\a'�R����T�uk�ŉ�=��Eh.;b���pι�0�����ػw֮^��+������~_��|p��:�S���k�~�!���ek�Ɯ�Ȅ�8�~]|�͙#�F}��mx3�,���|{��Jn��6)O<���A�� R^2��n�f��~���&n�_��π�{�i-��<�[,gS�]�b�YK�B1��g:�v�UMun>gݚA��~�g�stww��~���NS/��R7����x��/����&�I��5�����K��P,�F�rFC�K;;;�E&"%I�y��W�-M���mW�U��S[�+�Gd���W�
��C���\gʩ�����<R��x�>8��lw.x�e~�|�(�
�hh���C����'�����a��jK�|� 焣i<����]!ʶU�����h�#���=Ε�1�X�N�F��
Z������z^�F./�AYo!���і�`�ژ×0���~�p��r�|"vM_8q�X�Pc�й�xφmR��|��x�9�:s��[R1cz\�.$h5�t�̙%A��S����$D%�����^�� @e�:>��*���I�U5a'��y��E$��5����|t��~,�3���ك�E+�x�\t�E!�\0	��(�(f�^�����`_'V.^HF��L��ph��y�^rb� �B�Q>r�d���z�����6�����BV]�%�t5b�qA�[��J�p�U�a��Y�$""�{��gq�W��熕���_�VP�v�ێ���������ڮ�HE���@�˧�맷n�<q�y����}7���"ſ�`gF�☜�c��w�\&��\�X�0ȓc>�v�54�K�����fO;���S�͘>ód���&��#�x�JlTV 첽`�P��q+�B ���8��J��q�h�P-;ٖ�"����x��-Ƨ �E��Y]g�S2x�0�����5�'�����A�׷+c�����f�6L&��@UtA�g�xV`E *ك�%tSt:�y���;s�E�(�VL�/0&�Ae�r޼f��x6�*%�3��Լ�����AWL���{K�M% �"�0k����1� ����<T�.�׷�}B>��XIV$�����]��`d�I
�d3�)P�1����?����y�߰����u�]�1�'.)K�6�?]�P*p!�K�*�N�'��76ឫ.%@�����6ȌY��g�|ˌ2,.$(��轶$[���Y���D�GTS���2�NE��#sE��x�0<�����B�v�#�+���Ɓvtuu�q�b\��L|��C�=�3�(��}�����������F/��Dc1̜1��b	E�Ӛ�t�B��CJs��5��18����W�@45�ǟ݈�����}^��"#����k1�m&2�r�~��C,EGK�|���M�ށ�������ljD`�:\��m��Ϟ���(���i�t��CÉ�������~哓]_�Q�ⰀS,�v�wO��:ٯ�m��;JYdu�O�N��d2�-^��U����t��W�>��s�żh�c�q�d�F@���pNib�A2��ЁZ��&�f2B!��S����Z�3Y��&8jg�Q8T��L�Х��,WE�����"˿?K�G�.Ӱ+����cz"�Q���/�646N�XV)/�k���%[EhM�Q��t����`�t�>L�/4&�Ae�ա��iI��	%K%o��Z���e��ʶG�:K�je�f��`����H���!�������{���3)2E�Xb_��d�5��rk_yϰ|�h_�/:w���jjG[g����)���7�Z��M�R����5�+����9��-��ņ�T��b<DS�,�Ǝ��׷�뗬�Ss���8d���ӧA�3��3B�]�t�_�Z�9q�i/�0p�*���̀e�~f�V�� <�UQ؄lA0_�z�`:r�4�uj�w���>���k@�Ņ#��D�?m��'��E�G��ޜ�x繈(�~豧�t�"�`�b�J�߽��>�͝	�X��y6V_z��8�g_}y����FFW�L�a"�+�7��+p��wb��n�锉�X����\�"@��[?�Y#��kC
�|  ��IDAT��Ȟ��8t 7^}	=��ɴ��֮��K���9�L� c*��c/X���G�o�5����O��Ψ,E�(=�J�fD�ᵴ�O�3K4Ukt�=n�Į�F�#5
�3ӬS�#:�*"5�:��b��݂������!��XDI��6�׊`"e���V�'S�����
~�1�S�T��Z�d<�9�D��?�B�kt]?�Ρ�T�r����i&Q��*]Xh��$c�̻#{ƾ=�f���'�ؘ̾����+I���s^t�e!�����Y��8-Ǽ�e���1��H��-��s�R��3�L���� Y�3r�
^��.{�P�"o�$�I���������j|�?Kh��F�h��d��;��15m�cJ�c"Ev��Cs!�6#�v;2f���tvOF�al���U�-��j���9F�[���UD�E:���\�D�,��B
�%�۠��j�S§ �' �Ӡ�T�:��_�QDUH��Xf[���:Wqw�P,��dt���)2��X��(fOi�Q2°��HDG��{��;n�s�>�=ݝ�	��s���>|�O_�fG<»�o�p2�[�Oxc�lݽ9I��"�l��.��u��Fʲ��#���G�(X��~�u;�;�\��Z��/~���W`��b���ԩ�him���3��6O<�"do3��6b��(���hl��p,�(���w�'����������W�'�WhT\)9��	gb�T�F6������
�r �u;F:�b�H�I��fV�d6Czmdl�=�8>ܾ��9��v��V(��:��T0�Z6+�߹���Yh�\�[:��ߧڇO
U����O��h5���� ��o�&�W�|ŚD2)�D�A^�Css��l�x�$Sq��a�;�۬�dI�:�v,�D�01����$8�d�����R��T�{�YX"�/H������ޗqJ��!��d�`%�b�`�޽�T,V�Ig]�"���*�)�9	�&Z �5�4a4���o�(�5%�s���<,i$���x6�c��9K��>��K%Y'��B:���p�
fQ�D�/{5� y/]��8�#��6�v��g��mPM�>8�t��<�W�@N��#A�6)�f����	�L��� �v�B�;�?�x2.�k����v�"�5H�'<���عg/����>|+�,BWG/��Bc�G���e�t��0��o�N��2��淰��7�|�|�(�Ʈ�� c�A<���	�p���g������$�I����v;]��)�5�K�#�-�ǿzW�9�~��x�_~��� g>�]t.��"��9��~^��D́�c��%0�]Ggo?Zf��u`���8�x?��r��Z���뼋������/�������5:	�Z�3��P����r��)p��.�LpVn��;���]?��fWO��9{�렣�?������;�����f��.�G>W�e;[�v���:�m�d~;3�@���zR��Ԛ���@��~���t�'���|�x0��mG�����,@�;��r6���t-%#��L��`0x^���/b|�1	>��9�IR�&���<�XUw�ީ섍tV��^hQ��༬��T����b��d�-k����������N%G螅�L�7R�jdEm~�j0�B��jcjhC#�?�������7������vݕ�7.����
�J�n�H_jNER
�Q���x�5A6�M�*����u�Xb������
�"N�I�q�ܐ�9ZS�?��F�έ�����)�t7�<�gds"[�U�l��o��oOT�VհU���, EӸh��؊��l���I�8��!k�a��q�iKQ�%)�rB��t^YԶ��N�sj:]��w�}\����=�{�E�� 7��-�C���szq�w���#����n�	�dͼ�W4�5��l�K� 9:����mƾ�^�;���>� >��@sS,],���2�Yh�� M��t��va����'~��p�M����h�ނ_>�N�̩MR�C�ǳɅGz����g_���=7?m��'�Wgp덗��(6���E�V%{�`�k��a��s@ÿs;\�߯�}z�F1_Y� �Ɋ߿���"]��kE=9���Қc �_��T���]�-[������k�:*]%�05���Wv��ƆwG���n�'W�� �息�S�OΤ�����s�.r`��)gt�M���չ��)2Y��9�$8�6~���L[/���� ԭL�R�&��9`�q[�2�n#��f&�
�O8�rg�Q��QU�Z 6�,sŲ�+����92`@�/�3��=:�AfW��j:�vfX������"�Y�54zOVq,�+�ܕ��$$���&A����S�&Wu�u����䈹��C��G��-�\��gLE(��[��Pg����A��g2pV�%�ӥ.��d
�@�0Uy��^��w���V�*���p�L��΋P���h��G�;���1m6'"hv���� Ok�Y!���'�dut�9͍�!B��{�n����d���ñ� j��@�l��|���{u�(qB.�S �Ʀ&���G\t�h�Mk�jב- J����-X�%�ફ��{�ih\o��<��������1<0��&��+�&`�a�p�Wc��7 P���+���`����3	f�[��l���?8w����~��s���y���F09�*�ۘ�MN���JK"�=A�n�;	8[����؆��ó�>�]���/&�2�f.�s��Dss3֜�Z8}^'l�]��� ]U'��m���#��`S~���
�鋂{[!0� 8���?J��{?��=����'o2@୅֖&!=��\We�,Lt:ʚ2Ţ�nh������9����$88e�l^�~,�-�)�f��z�"J����mF�T�2l�-cf}��ц��Ǘ^��(E�3�K:\.3����Y�X���m�H��-r�f6_f��-rٺ���x"���=_�������f�eãw��YO�%��{�#��@�@�6Y2Z*E��S]/:�b.��ӹ4ܞzx�>���W߅��p����8����jk
\=�%���(BW(r!E���H9���l9�ʭ��R�01�e�"9�ё�����Dϱ��Q�&�Zf�`g/����k�#���@�[���c��.289��j�(F�B���8J�-X�Y3�'�>��H�7o�J���[��7�yG&&p�u7�ŏ>�K[wc޼e����CEptSf��U�G<a���(j*&���V�"����C(���m���}V�Vǁ݈1%�F*��4���PdL��|%$���_ހ�N[��k�,��n�h8����Χ��ĕ��C�e��]����wg�����'/jt�cr��2dBP{R��J����%��[��+��� ��\6o%����}��w�}W:v�G�9�
��<��XC<\~����k˚2Ry�XiKZ`/U�Q�|JF��-�S��N�m�޹�l�GT�<��c���vw<_��UG�(H\�%p0mj\NdJ��MCdQYΜ�rrl#�
M,no?ě���s�Ipp���BN�)�t>cؤB�ZDS^(
��m�lB������BYa��@08�
gX�g�}��lz&�����V������|�B�C��s������Q<y+�L�!��B��� ��V�����}e�`9U�	Q� A�O]U�������r���2��.(�E��kQ&���( WB]�4��x��]B�`�6�t-�Z� )�(F4��6���&:8�cV�4�}���Y����#��u̰���->���N�O77R�><���cp4� ����}�49eࢨJr�`�eS��!r��e��l�Tg�q6��c����3�E斛�<���w�����.�dЎ�N��m!cӑ�j��fф���y�1����]�(d,�	�D�|�Sq�<n�Ƈ!:�<MPwo��1��n��2,�ފ7^}	�pC����X��Bq~�Я���Xa>4��kW����~�ܵu>7:���T:�y�a,xW�9�xұ���y�v��p��G,k�B`���+0r9�Ù�6.,�+��V�rE� V���oFf�H�]]]�###�55uw6����C��,���s�=��ʫ��`RYϠZR�6��w�U��AU��Ԃ�j&�*Y�*V<U�d����VH����\R�j��9�t���D�3��)��:�v]l/����A�k����
����c}��cmmҿ�8���c�2�~^��p��KeM�d���t�fX��U����r�{��P�<��D&2_�}�,Ɩ�?t��7-E��f��Ҷ����I��E뼗�+���3�tA�����cMG7���\DH#�}$_�V[W�!iP.���rT�dY����?Op�j�3oA��N�h���ҝn�X�F�����#Y�G��Ǵ	/��B�7��S����Ln�I2I#+�@$Ԫ�dr�l,���92�Pq�0GB1���,[��_�l���㬅�?֍D6�~���uS�3Ǽ0tf2�|�qQxǝ_GK�BD"�tK��p%zF���ko��mx�9̜?W�tŒ�X�l��+�1l-5�8w�B\~�9�esؾ�%��M���pf�qW9��"&8�`"����wc������9{��V~��#�9ډko��x�mz~����[o���ǅ��|��#�_q:���c�118��Ӧ�A�m�� n�t-�@��^����wDC�����?EO5���W4�ә�s�$5*�iܐ��VX�Z���N�Y.��م8�������d��Z�b�ķȩ��b1�y<���3N�m�ގ�˗���DS>���-31C,3KyT����)]�f���z��GHX�~+)r������`ᑅf���N��u@	+s�4�&�g
��\n8�.�%,+ӖmgwUY��׏��.����'�����$8����v=T,����������j��0�?����X�3r�'�"��)�����L���WDO��9ƫh�y��)��,���	�����H�f�7tRe폍�aW{�u,��6o�`,��)�o�H]J�I����P��x�H����&��yk�	JJ��Iӿ�}҈$᠈�Ȳ��ϔ��@�ظm7�\�\��i3I1�n�C���t}��cӦM��[0�hjj�9�� �k2��}��5�`CC��:���^5`���.Y��u">DEL-�Ĺ0���,UӀ���I�/8:8��{7�*�x<��d��$\X�x1�[wa_G/�5u�� �X^<ܵ>�"���<��(�;�"�񵫱�����1:<���a��� G�05ԏ���$�홧���}�'pt����ݷ���pӵWa���?1��n�:"�w�v�˼<G鹸�j�ڦ���r
g������
��7�xN_-�.9R2��.<�@��o�`������?�͆⾤�a�G�L��G�by�i:_��ݙdr�����f�R(�u�h��v�l�~��;L��<��3��=s�x����hL]�l9���Z�'0̒м]ʼ�UY&���*���8���DQ����座�IY{��|
�:��e�U�H�R�Z�������O(J�C�/1`�V__/j�xm'�	Q{�[��MbSʤLd=�hd�p�T:��I΃?>&���GAW	J��eX�\���i�r �T�CY�'%#WEפ\Zv�c��p�`�2Ol�F�b0�B���G��łh�̙e�ϋ��Ud3�1M�*�9�N$���7�oW$�By��H�s���ƃ��k`v3)�jȓ�a=V�؊%:;xKAtP,��QG o0��H3;�`D��\d��Xi�_?v��b��b�h��Ӛ��	�! �%��юx��'1|b�"���nr�hs��"s��I|������m��<��V445c��%p9�).��py*���u #[Hҳ�4ܭ�06Ѕ|2�#�<���`ђE��e���~C�j�-�e�"	�A�g��|��)P�!��%�ľ�b��hin���q��`㫯�{psH��>�v�jd���}�����]((&V]r	^b�]���õ_���8���&�kkk"o%r&�D:W��.�
�dy#����ރ��1Q � @��Q�Ι��֞)�sǞC�K��������Q��ar�ݴ��|w�L��%n�[r���R4"F`48zf&�9GS���_~���ֆ�sg�*5=e*b�(2yY,@'�T�����X�����{N�W7��]Q�O A����ҍ9]�2��?��6�Q�X��t�f��0�*��x,)���:��*�%�������-�6��s���l���69����^l{w��)���E��4�*�ee�%�Η��)Rf���6M��;)_,��D:�Iƾp�����K]���|�ǡ�e����D��K��Ȧ�`�E�����cb���~:��$�K�d2][JE���[sZ�U:R2���L�1_P(�6�V��탤��(�j�����Q�Ί��cYI�Y5��%��d�����E.^r��T�p�z�-�r�eP<5�(2oj���x���)����Ͻ�;o�躡�\.�C�8�r9����T�.���w��G$/c9T���9�ba�yHO���z�Ysf��	�ma	#�4j�g G�*�ڵ��yJ �CEʲ�7^���lE��A���+��qa"Dm���j�����Ĵ:/� �7���"G��a�N��j�x(�w�|816��=CR�y��iz��{D�Ú+��@w/.��zd#!�w��!F��128D��O ֎��n��L�7�=�+�[���Q�܆�X
s������1}J=���r������u�\�D2�����`�^�;��zf�$}� xr�i��7�8�N�Sr4Y?���#[u;!���Ӧ�͟�P+gC˝V��[���5L�Ľ~lO
�by	��H���]�vቧ�!�\{�H�E���w{�����R��#�Vt1G1Nvbb��֯��nw����tfi\�)����Z�/ծ$����BvG�`��/r,W��G"^L��?:&��o�ۑ*)V��J��W�	�Hծ�D���	Oh4����4�v�NNM��vۂ�t ��p���,��x<R�L;����M�;��U�'�s�q�)t���&R�ܩ���i2e56�ǋt6#�t��oͤcu����K�󬺃��ئ�xd��[;�cK' B��d���JBV����ӫ�h)�ŧ�d�ʭ��%E�4òI�t���Y$���q]*d���ݸA�a���x�}x��0J��Ԛ�	�v����p�_G���h���d0�0IC����G2k�s�8v��p\B��cM�^�@������̙���I�%�yZ+�r�-����#�-�Y;�c'��;�p�k0k�l��G^�+[w"h9�nlA��`$#)��udr�H��O�s��3�L���"LN۠�{��M��y1o�6���hA,��p&�mo���ο�\B2Y+� ֑�Q�4��7�E~x/����^�hm¾�;q��A����X$*�V��&�ݬ�h�?����0�e
Κ���}p�68t��}86D�$����]z	��`��@{�7w�3Q��,���� �+9�g���o�lSnVUm���5����My��: A�.i�Y���|���k���ݷ�|G ��C�X�d9�<t�M��)�XKB�� Re��d� ���Dحl��V�zj����� ������pkCKw,���W�0%�q�P��P��O�\��`��k%8�.�S�~v�B��c���
��$����෇�mʒ�H7GP���Kr�̜&{��6g���XT�V.J����ټ7�Ԣ|o�4�G�CJ$�.U��~�W�"�l�L$�x�O�ĹH�@�1v̌�	Lp��C�F���H�ƍ��9�xq�{���sܯ[�C3����&���灷d�@�����]��I�D� ��=L�j�E���!�%�E��*�߳��E����0��ǒظ�Ch?E�v$"<��>6L2�
�����0u�\��,�����z��I����N$KEo��DH��6ŏ���H:*hX��J4ST.ۊX�d�(���
N��
�����Qa�J%i�^c+��AD^�"���`R�bolB�Hї�D:aP�X���1� ����p�ܩH��X������O
q&n�䭫��>�9�΀��c��>�v���0�����`�Gcˎ]�46(�p��/���7b<��Dv��&�OM@�?���]�nX�G7>�ںV\|͍��헐O�qƙg���APT��)u��sˌ8���ph��Zf��2_�{۞K�tt#�@�:�^X�_��@�MUum�jS]l�I��˵S
��
\n������y�q���ۋGϿ���ׇT�6��=�K�
+q6U�6ӱ�ul��L�"��iδ��2_$�*�
�@]�c]���v{+�}�TR|g���/�6��$�$Z�]�_��*Fʘ:0xb�(�:�I��?8&��o��Z=g��Q�2��^��U��꾙X@B��zEU,s�Z0̼gl4���З
��bY����툪y�<)#]�vT
ު���� ���ϓ���}�\�X7i<ͱ�sw,��W������yS�*ML�����כcm�,}��gYޚ�� ,h�@����f�*�PN3ʜ�Pʊ�=���Dw����E��a"��ӯ���W_��w�<�(l�x� g�d�	���z�@39��t�8��� c��tDv��M۱�x��w*6.Z���#x�p;�w߽�V4@(&�himD{o�.���/B��0N�;�=�Е�j�1�l�r,f�Ј�j���X~�5�X�v�c��{�btoE��\�۶mC6�A�@BA��Z�p�5wxx�v|��;��q��o�^D��hkkAM]-�{:�&ÿd�y��SO��+/E���k�>��ga��G���!8=�'���]G)��y�g�B8��'@�_s�e�,̘֊����bř���pѪ�Ec�#�zW��>f>�ʫ9�M��ܐ�N8dY�˄@LDV6I��� �����d�3��49\&>ڳg~�����#���?��Ұ;ݢ��M���iy�BpT���'?Wy* ��(j�e��/r1?�����?�����d�L%�ve�qZ{l�jj������#�I�}������N�,'�Pf09~��5�~�Ii�&TR��F&R���.���s:��
d�9'UѸ�9���`�;��S�?{8EG�P�u�2g�_�����9a�%Uy������RZ���"{#�F�&&�܋�������л��Fr�Xx���K�%�L�?�DV _��j*���hc�NQq+�$�2)�%!\�}�I%���Os���Pt K���������&�v�7��3O�E�L�(H�"U�c����/n����q���GS�J*n�����s�@�bJ��,�c��L������W^�F�.]ÅSVa$Ƃ�F�׿�|�?���z��S�S�R�4Ni���i�����Aъ�I��B<���̚ ��G�T�7�aժE�'�;}�,,�7Kp00\(A"��� �Ӹ�2g��E���O��o|?��N<���O��[gk3>>zSjk�����C�Xr�\~�Uxw�vD���`G���Ώ� �Q|s��&�3N[��{��e�����`󛯠��J�f.�����n�O�������U��9�k��vĲ^\$IL���(�z
�f6J��U�s
�sK�;E�!�I	P�#lW���B��oo¯~���Qw�]HQ��Bjn�rEJ�*�|*�aUG�T1&'�a��O�=�O5�3��0�pxt�b�u��Q[|�|mv�ܵ���.�����1�p�;�-�F[�T��]�L�����RhUŪ/T�m+��e�!���s_|�JV��6G8��/��19���f���x���2��m�� >G�<Α�ep�>�)Um�*TD��EHα��T�ɐb_$��?�ӝ���a�"��m'���q�jS�9y�7H�C�-C�1u��h�&HV����S� 
'�X	�((Dց A����Ru���`,�?����o�o~�<�$l�z:�M�(����1l�u
9B��Ӛ��8�7��C�mE���:6�N�_�l��A|p���n��
̛ۊ�Ӆ&�#}�������=��'���[��\����D�B�,"k��(ߢ���p��aG��L�7]��M��ֻG"<�dt s�N%g������	� u1J&�4�S�y)"Jgrt��x��q����W_��w�D>���"��`������K����/�����p���x(���)b~��!���n4zk���'�����^yg���f�����8���Q��>z��=�2�Z���u
B��p�ek%��G];;W��{/ͩ��+a�0�+M� |祐��v�RُL#1��pԸ���|���eJe���E!x��Є��<��Cؼ����`��	Վl��BV(����\�_� ��|s�@Qlsr��U�[)��9M���}��O��3�nhl��W�o�5G�����=S�Jb{�t�UpP���x=�N�Tj�����+����̚��qL����$�{��0��8#�jA[ d�r���:#G��[��UN�C�H��P҅/��q"�v��o`�fY�h4e�BiZT��햜.,f�'��`O�(��y�Nl�@���جP02e�ƍ� �>����7���?�s�ݕ���_Hg��y��3Hd��Y�P��Ȳ��bD^�2D��HN�Č}�H�r}��p#�R&Q��i�U�q��Af鸁Z?����Q�o�~��|���{��'^�N���l��Z�>p��вr&6����hB�" �t�d��~M����Ǘ5?|-:vw���~��:���q�	���⒋/�O7�
G�$sE��n���$Kt<�KAft�ǻ�b���;�ཷ_��sQX�﾿y#��D.�%Z=�/\�����C���p�=�F�p��Ӝ��sIS��ܣ�ƥ�܎�]�NHB�RI%5u�x��7����\�G�}	G�1}�LLm�xi�n��Z��i,Uý�x��'��2ܦ�ih�6�H{?>$R�M5^����n*�ǡn\�j%�ٔ���ѥ;�+�z���a�$�09�꣩�i�Ɠ�DQ)�LSn����e�LB1��<��'��t����dԞ�.Zz�hg��ۀ懙'`�1����ۇUYIʗi�+���Qne<�\[I�S�NY6��_8j������_�|5]ɴ�T�3n.@�-<��r:tA�$(�S���R*���+&��l&S?26�<1n��gL���~�?EX7��e�d�m�yq�M���[0h��쁙/�Jm�*їK���q����V�l^��8�9�((*-x���+���mB�P&`�șWs�z��tY���hJ���:�石d��?a����M&��<���U���`�	dZ��K�p����eҌ���.Q��E!��J������K����'�p�"�	%��Ko��ǽ��6|�a2�~d�Q��x�Eذ�#��Շ��9�>2l��(t�2�����d:=�z+�B��O�����_?���\�����-$�I�$�F���=��,fm��p���"|'�;[2�m��8�C%�9�D��ƃ�N�0<8����E����j��U�s�	��%tT��4������#xk�S������;xl�st�TD�1!��?8�'7����]oD�vX*sͧ�%0��"[ 4����͈Ҝ���}�z��q�����^44��Q��(91�i���>�}�\
9���ݷoI{���?y����h����$@�+�?��km Ϙ懹Baa�*NU$[�,ɎB._8�7����	r[��?\Bvmnkk����r��H,do昡��[\'�0��O�T>��A�l�L���rJU_8s�C�i��榏���9�YN����d�4�9�.A���@�4`�l�H�B�3246#+���1���c|�P�>����f	�� #Q�6�vF���h���^�I+�]"t��2��`0�I���=������lE�|H���{j�<$����ɼ���6��i���L��A���op4X�j�_�'U���ՙ�~o�K�,}���|�]��Z��ˬ�V�B.���Yl��a�"�'K�
O�	�$������%�26vo���GCx����w�����-<��o�1b8��u�⺫���x~�N8��(� �.�)��54"O�su��k@&���Q����U�B�@V# A�O�y&Jt=g<��+�����F�T.A���,'mSL��:���Nҥ168�|�@��=&�z{Σ�{���HY~�#�b��{��K0;*�
*V�d#�Q�
��,�D�BVܻth�^܈����{�߆{��!��,d��Hx�Բ\��K`�0EZ��r�K��g7oFJ��K�቟��=���w:�T�>k��fHF?ڼdq�2MNW��
v��>p�}������b�[�E����,eh.t&p\�B���bm.��'si�SՊ�u�fO6��iK�-=���]�px����+������+U�Ѻ��z�r֠Z�]�V8�$�b��MQS����l���`����0��]W�d2)E�>����WAI���m$]�=�̜K�aRm���Ip���0].���d8뱻��[6DU�̑�C+�h<9G^�,��^=*�K�L�S`:-NYh�늋�J��!;�b�ʋ��pVks�XМ�����2����9aMc �'+�����|�[���r�]�X��=�:*�����2�y�n�<�� 9<�)�V-������Wʘ�R�$�����-�FЊ"��NR��	`0�c�<�[o���v"�Q\p�Z<��s8�?�9{��K)/�6��g����|�\����E��d.��ƀ�TGF�X�(an��H}�fl>�m�D��D���5���T�HǸx�u���[�D1Ć�^A�Z�a�L,$G�{lP<A��͐���k �$�|����t\E �ݣ�iS�1�R�N��N(b/">6�c�j=>�q��x��{O�q�57��qcb<$x�5�7\l�33�ث@?�M
�G��MoĻ��E��7��x���g�d�bù�B4��� z��M�gs���f�b�r����t�ν��x{W{!�4�N�zu�$%19���wP��S�m�r�R���4�$�g�"d�Zi�M��{J܌Q�m�F&�w�*�j�E�ᦈ���Xd8P�d�uZU`�[��bC.��{���������/mxpCp�Gۏ+�2�&�ޢ̊LnA(�V��Hg�|�(�̔l	�hmݝ]�_6����$8����7�v�1EO�LӬ)V*|K"�UD�/�cX2A΀#j��#A���Bc��Q���m�ly�DF@��H�ܭ�	ǹ"�TىZ�U��Piqd@P�t^�x8-X��x,� 64��ϒ�����K��֖}��ɘtaM]s}4��rd"-N������V�@�ʵ�>�r9�h��Z�>��l�~A�4���8��	lx�E|�֛�p�\<��386<��C�>#S�`7��8@I�[��̏��:�l&��*�2&����-<�y;�\4�(�@�mF$o��:�M��&Ph�s��ȩ[y̨�źų0���������������C���64���%s砉���c��-/SF���l*��+@�ݮ�{ĵ�|^t�t!��9]�k&����qإ�Uk�ݻn���~���4�iA�%vHt�l�횮���^�c$Eƴ���}/����=����"~�^}a�Z�=�X�p:�tb���u�0����k0�����A�p�eMe]G::���=dӟxG�Z��L� |UFe��2�E�C�/���K˽^����;��R��%h�U@���=E��k8�Ϡ�^-J,����(�����k����<�����?���e�In�\�m!��2���98�5��4L�Ś�G�fѯ�b���3�$8��A�|�WƊ�b�d��%<�D�pA�h�����@�(������J6O08�/ƾ�^�b1g�l��:��F�89�ExZEZ���r�@���٫r������2�z��L�9Q�e�#��7l�Y��/~�՗K��.����@y&E���	$d)f
��\��VEڵzP�u����Pv$I2
��89x�t��������ڌ=E}K+9C�"b��
b8��K�ɯh(dM��/��]*�ڄ�)Q'RrvYr��n�-�q�m�ٍ\,I�K7GL,���ջ�\��KW#>x͵���2�����6"<���wq�ʕ�in�ᯩ5\������_�/��e �E�#c���r`Ɯ9�D!C�K#��L��m�ᬋ/�w�y~�Uq]f>E_����$	�E}A��::��M^!�X$���sS�ePdk�)�7��{�p���X�h1"'F�T9�V�� +�0�; ���М^)��G��[�#<�UW'����3���=���vtΤ�bE�6��oQ1���U���=MdpL�XM��+�VS��F�P�M.w2ZI���s���O�M���7���Z�a�
gޤR���*~�Ȉڬ\>+��.��.�q���)�㺃�����������I�IJQ�d��3�s6��؏�IǼ�U�Z��^E�%ݡ��hlzhx��C��H[�f�IM�h���0b�·��R1\�T+���bS����1�|�X���?���a%��g��o�)�����囱�H�-���[��3��ܹ���Zќ/�܇�l&T�'��]  �
J�(��l�����!vd���S_7�� l��&+d�
F��k�%����9]/=�l:AQu�D�7��9��2�ȉ�\&���s�yF�]Q��+0Ƈ)��bzSb������Ai�߽�69��HW�� [�{��� �1���1�G���ƵN2^a:?S��+Mr�y��q��	M�9����9'�bs=-r{k$8��7��3��7�pv�{2��c&�As��
 �!�H�6��	
f��G���q�+0���G�7�X��xc�&t�oǺ�k�͗P�Ԉs�9Ǉ����Δ����002����B��b��17�+><�s�U��Ë�[_�As+vƪ���ƃ+Lè� #�5sR>[���P�%�[!:��Z�>	�9�bP.Z+ň�`YNx��?��G?�����*���i]��N��ϡ�u*�i�r��J��M>g3_��s�YC5��9&���uu�I]ՆL���$���'���I'��,(�b!�q�̤P.��6���%�ˆl�wtR����|�*C*��H��q/��4��W�[猁�[��rK�\�jиFB��y���ӳ�oo�_���w�����;��$��٥d���<�@ ��DN�T|ᬀL�I�%Q�(U��JCE鱌���3h�rTm�l0I�w��G�C��U�M`q'�Da#Oz�bCI���\4��daH�]���X,�چ)�*[�L&aw� ��幐a�E�H�R+�5�na+�x�I��tvw�7�<B������h�r�nnAgo��y���L*U�"Ƶ |�eeM�dL ݡAs���8���4z�{�l�b�h���)����
g���c�ۯ���_Ǣ��pt��d�]^�}^�A�{hjB�>�K ��BOE��e���ѻ�,Y���6�)\s�����!��í*P�H\3�G�����+�i�郏"C� g�s{�������P�f�챬7�HR��+;8�����=�߿)�L-�
�r���/&���.�q\�����Ŝ����6��6g�&i'���/Ď��h=���c.��+�XC��ɤtܝP坩h�`�<�ѨpՔ�%5cd���ar|��g46zS6��[L粲��y���g#�T���0ev.�tN�.9&EL>��C���@ 墟?7s`˗�S��*J/��roqY�H�LvD!��}6��N�fj^��"E�����p4:�D���$�4���i�A a���Y�|������t��P�D�A���d%\h���$��[�$�e-�o�ުV?��,s>�~�b���F��ȶX��PԂ l0�ɴh����\d��.��b8�:���q���ts��T?=g������%����Ȧ�ܡ �ٳp��4����/��Q(�m���,_�5W���#8���aw:�c�,6�I	�nQ,�AH%�P	��oe�X ������ٔ+���3faΌ����[,��9@��d/=�����kQ枠��š9]�R�*�bd2M (��]��B
C��hBl|� gb0y\����W��s`��U��{]c�Xuյ��U���h8�>M>���%˓��r���oH�	 �3	�ڃ�izɲ�{z���S �J��QU��U(뷈�n�u�>\�KAd�*��*u�K5r�����$K)_s͟��_����u�N�%l6)`���'E�$gy��MƩ
��.
9)g����F�A�dJ��1	~Ϙ:ujR��%+c(�/Qs���Ȼ�sJ�@Q���N"V�&+	���F�q��P��j+�����&�_I���EW:�Q�
�?�W�)z�"��bP�+F�E�c5d�"�)Gwq����� aÆ#�VAyk�Ǫ��gz��Q��2)�ru]��VEX��lVy���!� Qf9�r]�r�cy+�b�Lz&�T*]�x�E��.r��e�l*�"�ψ�Wl��v	��&��%��>̾h^{��e�=��:����v�q�'c20� H�A� (fR\QY+�SXYڵ]��]��~v�7��JT�I1' @"D��`r�=�s������4im-�E�氦0�N�����|'}�?�Uy��3�D��'/�Y_#r�H<	®5Aʦ�\���;����j�~�M<����<��˨��`��s/��۷o��m�D޽��v��)��ϧ��rF�.+���f��S�IF"��	�,�hBp���i��8l�s�<S�����	:��X�t6���
a�����i�Z�QE�+Ž۷��5�Hcs+�r���������+�q.�����^D(�A�����Z�����j�PH);���;�Lx��(-�f:Eێ\)��rѯ(�x$i���*l,�HV�Z�N(�Ȥ�n�p�e�Z���:�ua�ޠX�_�NV����RI9B6B�:Ym�|lp34Z5�/_��s��u\$�"
��yR���db>�a4��J
jy�?i�z�mhs~K���^d��<PBܧ�@�ZU*���*I#z|YL�~v��y�L��֛T���<�t�%�=�X� @N]*�e���tj�0x�y
e�"چ�Ҕ �������#Y��=h�C���cY�LGj�%�K����6������_�C��c��?�T�f3�¹��/��n��Q�&K��I�ܨ0O�,�,�yf5�|�y�E�{ B�����/����j�Ե)�)�*W�s�{.����+����� B��ެ���707؇��)�Ժ�~ݱU���퓿D<��uU�'��â�fX�j̎��f��n2����~7�|
[7m���e��O�`|r����	̑�]�P�8y���� ��u����W�p8P�F,G���� r�\����0���������W�I&E:DG
{������&R8w�2��S𴵣�&g⌯d�J�n��n��Z�����{Vu�ÜW/�n1cb��>�	��j�ef�|�Y�������S�B�P��֤� ��kV(+�D�%,$�\��*j͎3�S��vPR����'V���2C���N�2��D,B� �H�p4w.h�k^��܉Ĝ�T���s�h��TT�������ס��G��T��ݜV+���2\�M��Ui�T�j&����L��X���6�R�6 a�8�'� ~�466ĆGF�|�@B��`j5y`j�]�F�ǅƒ�o�Y��t &��d���\0�xxd��a?8�[2*'�TR)�r�{��z����(�3�4�5��2�r�#x��lZ��3[m����ǩ�8�'F;憇������&��o�Щ*��p�bw>"g��d�G��T�d���A�j�T:2R��P*��)�p�e��<��7�B�ԨVQ	-1�d�ИMP�-��j�`Hc�i݂c�hv��>� &{:��[����}�o�����<�ؾC�������~&D��:�E�&Q索��-���2�)N����G�=8�yu�醵�+���ra��p@�hq^�eu�N��,�@��<+����'z�[Z�İ.�rU��ő��G.s���gi�;���1::�I%�[i�nZ	cu;R�w�N �z��U��޴��:�1�,�u]B0A#�����:��d��Y��%M����OE�����[gz���%AW-�_2��&Z��5N��^���j��K��<�f�:��Ԫ��yy�kg�����O�;�>��x��p󅶣�^�&������F��ɝN��-���5E�� ����"$m�cg�,�3��T �F��6;�5:���=����~6W�qOD�&r�dʗ�b@�Yo��h�Io�s�����k��j���I&ӺT<�hvvʄ�'� �7�/';/��I䒫T}���\�LKd�2������tPL�jfd:C&�n����}�k�%�\�'���u5L'�O'���Cv"Ǧ��Ӳ����8N��5�,f�s�Mͳ#�9��G��"�� ��%��ON](�T���p�5�[��jW4)K�djy�^�&�� Z�8*B^�Q�S��Y����1ôѹ��KH$bp��EGC6�+�|ؓ&�Y9�-��@��>�I�^�x��;��}y�q�ٷ�o�8��f��0?��)��I�Z��4�a����p[�x��?���8�����h[Ԅe+�"	c�p,%���Qf<42oAI���J�S&�����"�����8�����`XD���@��{O$	i��=�'ńş�����-XJ��ѱ/<�5˚1��"@^��)%4:����^��=H#8w�������^���[[��u8�Յ+�(�o�N_�3�� 6'4t�V�c�t�l_��a�ed���m��ڥqtd�tmy��[Vl	�yӫ�{x���W��R�L��˗/�����0�ͭZ�Ve"p�U�D�/���AN����LC޹�\�ז�
�XL�Ŝ�n�566~��Ċ8�uq��1S�&2���bA� �3=�ie~K��/&��\�:��,%�/d���W��:�D>[d�:��#o����ϖ�"'�)�������9q�N%�����u��yF�6}��Ii�o7*/1Q�p��Ҳxut����d4��Z����*��2�(��sYM$i��?�l���8}d�ylkS�]s舘�3o���v���̓F)*9h	`iJi؍FE[��l.�.3�x���W�׫�F�Qe0�F�A�[T�|Z��D*E%'�Ij=y��!��E���b�	���c�9y�G�B���g` �y����ơg�Ic���F{5r�9�9�ʭ��,s��O��8t���a��������19I  ��@�ٳg�z�J���bt���c�ںBX%�j��9[n?t�\p�����a�����}"�c4j�\"C������{��=� �D^��NR�c3^��v��~���Q��޵�f	�n�	'.���V�?�	�X ��VXLU8u��7��au��2�`5i��a��u�����#�p��
n��1L%K���o�hb ��b)Xh�qw�60��S�a��Et>R�tၭĹ8x��VOB�X�|���i�n~�{@IhT�E9�.I׭ vA��ttt�./�|���M'������o��z~����ܔ\fG,��T�j�5Z�&k���׫ ���)O�'Lz.Np�����?���sP.�.�LI�sW�;�I�!?3%��G+��I� ~��I��5�����ḅbW)W��R"�%#�H���a���S���S�'��Vƺu�&��9�`vc�g+H�o�2 �D^Ұ'ʿ��Y� ����v�|�<,J0'��Ԧl�
<۵X�]Fn*3��^����֦�)�uR.���cPL��J�[&�b�s�^�$U��_��N{L�^��8����*�F.�K�H:�	�}+���B9F���(*j���ތ݋y�v�%�v5��sShkj�W������w��J���v���E祋P9���s�`��m��<x��wKe��܌d,�"+�F���_~7�[���A4�5b�;q�CH��wz�Hf�AP"WZ�*3.ʄO���{#f�+QG�U\c��/[�L<�wR�Gu���d��"����y�Zl�i.���������h���go\ׁ�d���v�v�ֶ5���R��,�:���@�������c��Ċ�:̒���
fU��/aN���^�Yg�L���[Q����ޛ6�E8��?	��ŰX�{����iQO�i���2��
%�]
�s��V�i��n��j���)l�;;;'/_��n./wО5�V� ��k
� G/����Z�Uf>ک���lS���k��c2�٠Kd��65;@�j�8G\$Mį�>�L1_q�
��=��J�/�\#��w��TW��~�B��yi*-�Q����h<&�Ag%pPf��p��R���g"4���7��(�w��k�����:6OT6>�kH�X�~R�ԨիDa"�TD�ߜ�33�>�����5|g����Q���ҏ^۟���l&�oME�I��ܳ��f�1�^�7�u�b����Q�hj%�dM(ɚ�H�i4��O$o�I��zZ�l&9�,���ҦX�t5.|��݈���{��Te�5R�D����8���)��ڈ��؃�_~��־р.�����(�8u�mx����ݻp�ͽذanٶ'�{��J����^X-&53P4�L
#�����5ԋ���Q[[���Q��#�sp������B�/���n-�X�=�i�&��񜏑�i��� �at|F�w��}v��}j7����
ED�6O�S�u\�p�o�L�}dVܰ#]K�1�`�c�A����{sᴘ�!s���ă�n��߁K����7��Ƴ�=�����w��� ������_��UHdNg�r��qI����>���!�W��R�<ٸqc��{]g������!=c�Dx?W�J�K@u�M��Ʉ�������nm��E��گ7#�TZ��\W :)L�TL��D�A�Z��q��(�,�d�)�rO�8�F��������Q�N+%eM�أ2P�;���SLck.	�`�Z�i��L���3���l,�h�S����$4��p����kۉޟ�V~�P�	�~�ĳ4�𐥔JEI
[�FF�k�<��GY�J�Q�cf�%��k�mz���V��}��Ku�u�OlY����߮�����ǧ��Yڸ�b�\�P���������U�ܗ˃�d�����琝����󸅼��ΣH����Z�He�X�~������z�;�પA4��OcQ���c�]8s����zz�e�&dSIQ8�[1=Y�L�+_��ɦ˼�~o�E/�����tw]gt���=�װ�Q��{5,�]����,Ak�����h������u�E�j4��J2��{������$�nX��>uzfB]B��K}�
kZ\G�7���������o~�;
'����_�v���-�5ȡ֪Gj�Z�	��|�N���	K�-É�����è��E>�G{�b�����Ybsa$�F0��m���[\<�)Ii�����@���>���uN����e2���}_�
}4�T���:���D�������+�O����Ϟ�0�Ӥۊj٠�r1��T�"j�u=�v�R�P���bQO���Z,�o�8��Rj����՚�'�c�;��5<��v��$b��Y�2�zdt��ZC�YU���eh�GZ��#�����Z����"Y~�IT~�7���	�e �F���Uf=�Z�U��eԩl��J_�����y\��Q�Kn�$��\���G�٤�}Ն����)VD����������i�����=�5o:�K�����sJ���{?R�q�����]2�]��#�42 kc-b�(�Wu��G��_}�G&�Y[� ��ӱ��_���av�
:vm�������QSӌ�ߏ��l�z�XÖ�z��Ί��8�)���[Yq�Gw4�+�����`JkVZ\��```�_P$��A�_C����E�dA �L0�x2��?�"�!x�6l\�db0)9xg���Ʊ��!ٝ�]�z�]��t�bR̔ȕ������qad�g/ᶻ�=����ٯ_A�-�r�D8O��W��l��:nܲ��5�����pW�zx�h�,B]M-B�i4�ߦ">�X\&����K�$E��Ng��޼xES �D a�@�d���=T__�=<8�)Nc2�e��1h����<�c,����r��w�8:9��D�f7�Sf�9�ȥ�1#�'�=)I�2�q��UX!j"�m��|NW�,�Xd���,,��6Bcc��V��M�B�6a�U���2<؆.{y��z+Lz�<���b��\:��p��ǩ�U8gW�a������D�C�S�����L��+(��M�3Cc,�e6l��F]RJ����eS3!}F�_b��|a�G�����'����wI�l�S���L���.�����i%��
v����<������MFj睻Q:k����b��ر�<��+����bu*�\��jB>F`vUv3|��ع�xg�14:%���.\D��������rWG�0��z_ʑ�2��V��V���䤸Ov�]����d�i�����2��7�.���W������%rJ�P'N����$:V�a��[�"<�I��HU��k��`� �9݉��)H�,v+����M{� 4�Hț'�a"�D��'ϜC�h!��:V�2aȤ������	�$�8zx�-��T�=0���U�PP��lHă���@/���0a<�#�'C�tXgs�����h�b�_Q�/��C>{Ӏa�k:1d�Sux��ƔY��[���{�\�(;l��uW�р���J�@v�������A���of2ޫ.^��h�u�jc�m���ZM���#ǄG�vE��O�e5�Ӫ<�U�O+0�S4��K�9��� �!����1W ������Vk��YP_쑕�dps���Ecs�R�.{�q��Fo�y���q����PzI���٬""�_`d,fd��p�ü 8��in'*�W�s�|N�	��k*�i::�+��V�8;;�dxb�e=�����a�/)��݉���{A�h^~��������L���	�p���KW�GϾ��6�EC����Zl�r�Ϳ�s���6�/u��C���h���`zz�?�wm߂��]��m�`z	><ީq��AO�bb^|!��Z1tFSn)%e��砯и��d���Qv�S�q����Y(Z���hA� �\��!���`�����K��8�-]��KW��7�R.A(2��kV���?����xq�QLu����|�CPV�6�&(Z�v���(��J�BO �|��g������O�\:�m%O������b�r\s��E�K�G>[��b/����\
��{�\�^���"�i?���t&��n�3[^;�S�F�ʝ[o8}f:�N�3��f�g�ON�	F#�ð����*��������ӗlh�.T��~Ģ�t�H�A뫫7��|�F9��^S��tf�Ď����k��P�m``��GQ&V]��%��+H%2E��H\(��ax��y�dj���ya����-���tF_�/�~[��?#555�w��z؟�ZAf��3)2��B���3ssj��$�M�M�H�a���g���\��
�����狀*s��"T�$�_����ee~�y��b9O�)��MD0?C2�&��澡����a�?p�����?[�Yrf��ek^�ت6���ɔt��Yܳ�F��Q<�� ��}+~���Ѳ|1���ƹ'p������8p�|y�5�$���1c�+4����c7c���b���!03��(R6�r��~=�|�������*��d�9Y(�
-7���t�0k"��ۇ�е�E����<�ƍ��݅��+c8v�;�paݍ�/Z���/1� �2�hu��\,�6!�3�%m !K�G�3�T��怺������FE�=�P*	)�����,A2S�\0�U��GO\�ADGP��H�i@��2S�B�#�E��v����s�868
2�p:��[�b����W��˚���I����d��贴��M����ِ?zyp`��+o�w�|��{b!�p�%�����X#�Y�M|�����eB6�Õ)�AG���u�d���됻'��:�/	xlKT��d%�L�u1�m��j���Ȭi�ĜN�1{�(|(��B>�`K䟗B��nZ��M��H�A'�jZ���hh㕘m�hnW5y��.2�<�РNgS����%�^�����D�5�G��Z]*Ѽ?T��N��A��jޯ�XCTf5�=kʹl����^](�=�����Z��K���0[�/t�n[�q�|_ﶈZ��)�z.����]صv5d2NϽ�:vlـ�����ygprrO<�B��tAo��H��.��$)��c^49�X�ny��^fE�ˎ_~i~���$T�)pe���ϊ�RU�rarN0�%�&W�cp�B��l�[�i��X,!F�S��ƬׇGy��U���N���0���1��D� �
k��ڡw�J�Vڟ�!�1A��$����䶣�}��n�t��p�v7��DA�
^���9���}������{��|5;yezA��7�`w�@^>�N�v��9DSi��fTW׈v�/���7�^����x�R[հ�;�\~�dWخըKyT����F���J�T�$9�Qb�H�t0��F�t]�T�7>Ok6�0L��J07�S�Z/&�23'�J{tE'i�jQ������2�y��I�L&뜝�i�M~�h굲r�ʂ�f	��z%�V���ވ4ׇ����Ot�P@��+�M&]0,`�MY ���f�������T&�.�J�r݁J䕙���+��Y8D}m�� �ȁF�4�b!��h,E�y�ǇUUrQ��$�R!/_%ҩx�֫�����٨\[��* ��	�0@�)���Qh�:)�.��ލ���-k�l���8`���5�/z{W�7����m oW����#�w��i�ټ��zڪ]x��gᴛpݷW�{�������9�?~E�N��8y!Z�Uu��9�����h���wj�j�U5���a�ޛ�Xm�P{%���Vڼ8��%C�yYA]*	��J;؆M����{'`��D���<�7nF��Oݍd�$�en\��a܏����㧐6ؠ��P��=b�4d�~UH�G/*�V��n��k�&324��ZAuM���ːtF�D��2���Nl�D�+!0l"���#gN�^��<7�3[���ъ_�~�T;7� �"���(�:�v�t�xV���ɬA��lZ]ݪ����FEZ�T�� S(��S2�Ԫ-Yc��d���(^;r(�����+�� �M2��R��Օ�˵�+��+g���P�/�YQ�t�X|����Ҟe�;�>�u1 ����͜N����+s-�I�*�ef�r��$�{<'����s�4ׄ]�!y���8� R[kM�쎉@ &4���v����t1/��$bq1v�lw8p�F��|��^h����ǽ	)��(ju�B!����|Ep%}mԀ�Q;R�]e����e�Ģ n�1����dJ�F�G�[���;�{$D���J��@<���m����=d�g&a6�08؏[Wߋ���_�ʅ�X�ڈ�j��L�y���B����N����*�dU�#šR�'o�D�E��� �G�.�M�[��v�id|�Ĩe]����N&X,�rjg��rOxP�N�'����S���&����E0�H'ϞC�݊�t�lݎ�~��x��8��M���=�4�٨J=�
��t��w�Ey�%���S1�z���I2��r���Y�5�����cP�h�𼊂$�t��!�*8��0�y���l�bVP0�Mf	�LԶ�B<S�L�.LbۺM�x�nێ];��x�f�j��4�q�F�UWB�ݎE�(�� �E�Rh���-�B&�����;뫫'���ZIJaA��$Rq�'N��A 4ψX�r/J�Ue�~b}U��K���z-�6�N�,Q��gp���L���J�S� 8K{�� -�y}�R)f*g�(0{I.�ټmPcA��8� RUU�sV9�ԣ*/m�6�Q�����K��H �N�M��Q��U�9�AJ�%]8n��l��[0�!�?�ƿOgH���<"fGO.���HYIU��Ҩ�9%��f�	�+���*�F'�Zu6�u���/�Ə�:�q�}��jM׺�=z�6���<�����.3�#����Sd�Ԉ�"�J#�j�/Ʈ��ƙG��Uxx�N�d��{�8�L.����gP�XK��Z�������7%֗ #O`,h��\���ث��rQ"�eYx?��_�tHg3���KX�bZ��^U�p<����cfro>�[�E�\8���7�[�z���/��d��(�S�	f��"����tNpa���ކX4��=)nN�X	 �
i�iiƽ[7 ���q��98]m�rd��L�H��i���VD��(�V��d�����}509�(�K����RՈ��={�r��e�u�֭]�w��qnh
Y�n��:RNZ��<�V[Q��a���H��S���R��X��:��͡X|����q[�ctmW�PRc�da^��g5�\�a1�U�G+Ɵ�/�J�S���Z�JT���*��:�漍�Ь�[�"N�>��i8Z��!�x�J�T�-Һ�k�ey~�N��h��r����TX��� >�0!�;��M=U(�ܛ/Ȑ*��9���=`yj�C���%
�Z�Z.$�{z�Z������C��*UF��4�t�*����O@����o)J$˅qPʇ�Ċ8T5��H��P��^�&MS�k�Fk�F됫�q���H�7��;V.�C۷����ؾa%�;�&Ot� �E��p�V\�x5u�����|�ڵ�bNw�E^,�8�W��K�b蛘���K����\4(�D�絑�,���W��5�pw�P0��V�X<"�-B����S�����I�y�=Xޱ
k7l�����I1�;N��.���\��f��A������,��Ȑ�̦Q pXJ%Q��	�h�\�2��<����������wގ�����}7,��}��ՆS��h"���o�Q3^���HX�n��;-b5{lp[\bz���(Z�l���o;��LF2콙<R� ���bh&��AL6��S����n3�\�F��p ڒ��U�\dy%��J�E&���F�lI{����7�z��ћn���Ha�'Yz{{��X������@�
*D]�(��Í���R�����5�[	XH�l��g���ao+�ot:9�����)���(��Y�k�|��$�AJ)���"�N��ŒE��rU���&GC�d4N'ҩmv��pH�@�_��!$�S)$�Q�s)�6�[�`4Co���d�jbbrQrv�s[��M����\֝�t��n�NU�`t�r��O�1�W�l�ԕ�z�h���lN)�1���t6���N,Q��nIZr]&��KH/}�5NKZѪ���$�7�.^���*�D������lĢ�Ka0�q��۱�Wp��q477��_�"��� ٪�k�m��RɴX#.$ܳg��{�S�m������7֙��V'<��	����m�&}>"��<�S!N��g&��1���gh��@(É���'���i�Z��5�P�&D	Xtv��}E.�y�. g���a`u �ʉ��@��Q�ۍH(J���5=F�Š�{Oך���"�F�C?��S���VF(���t�b��/��n�YZ��x��	T�4b�-;qd輸��mAS�m~�rI�{�",U���5tn�H�0�;H 6�=����cr ������)��^����g6�	r���k���Ԍ��nj]�0jt:���I$"�t��S� >��B9c.�i�j���$�j��-�e�#n�e�TﳱV�-��l�� ����Q���N&���g�����8`��hJ�.'q0�$����L��)�AU"{����1Y�+JɜL���5� >�8�em˸/L�$�S��s����M�¢pnvK�/�AoT�lwAep�r���ox|���`3�ȇE�z��`I!�E�-�N����I�g,1%h����UА�h��kԑ��h1p�4���`F^X��B��"z癷�)��n ��!2 ����]C#[��	����DV�~2�T��F$R9����Z|����_�����Y��X�;�ڌc�bxp�o`ld��������_ác#�E&Z`^5$ST�-�׿�g����Y���t"��!O�LTE�
�W5zT;�d����za�T���)y�z|A�� 3[��u���{0���'	��|A��C��@�ʗ<�w�	�ކ_�}F�Ƣ����{��$B��*���>��)�#G�HE¨��F��u-�"��I��:���'b&��y�*��	��L#�����C�б۶n���:a\�ƱL'����!I��� \u�x��ql��Fl��S8{�5�Ş{w�`R�B�];�~�,Ώɋ�B�7��l����i."2=��3�VD�aT{�Hɥ�0�	
}wE%f���A��Lz?���a�k��`F>��VcP嫱�R���\���r����l �E{3�L�Gק`�B��b��#����Xl��V�F�Q������M�W��X��X]�X�֜�D���C��9�6--s��HC��D�.O�Ϭ��������K���8�F��ҩ)���3<:9G�I�a��F���h�K�����ʚ�:�j�1==#�8�G���Pz{��C�h5�lI��VW$C�c�k"�OD�:
r�l�<�4��y�Z[�i���/�Ew�h�Zd9�0O/*���y:��|�:7�41�m���Ci�k��:W*���dfN�O�3|���O?���hiY�lK��DCM-��
[��&�zޗ�-%}��GQSS�'�z��^��?�i|�ч��|?��ߠ�,�6#����D�K�G2�wmjjB(���}8�'�]ʕɍT�_�d�z�{�/>Aל�C>@:�˽���׏�g΢H�~+�;w���v�z�>t]�Aߤ��	�F?V��g��V����l��diڼ:�sr���Vҩut_{�Q���\Sd���\�L���W�v����PR>��Q�HY��d�<7T��gϠc�RX[1���w����7����W�$��ĥ��x>�]մOuF���X�����0�	�vU9Ds�'ɨ�	��H����#~�g�T����4q�}>O�����E�^�։xق|\��b�B�PK���٢\&˅ߨ��K,���˔��2)OsT�ԹB�埛[��8���
GMCI�Qe���pZ�`��Z�bq�l�DN�C��_�,+:�:�Psp�,��(\���=��K]��q�#Ť�MF~%L\�愞c��hI�i]B��v2&:��7��()��.��x�;�>80ͅ�"��ɤ\C��LjT�ڦ����!��a�C�}N>~q�.*Jg#W�Vn3*�ZHr�9��n��ʦ��[�q��N��r-֟:ӹT��U��t
*�LS��ڇo}�3�e�*�}e?9?
n�uy@q,��Bg5��c%^9| u	O<��ye/�ѽ\�҈���%/�M�ɗ��W�x_��7����=4�l��6R���!ef��R�I>8n�''�p0G�5#��䵇�ȥ�q�t���?|
�[Z�ڲ-�61�+C�Q��ct: �ۋ��,$��W�c��F􌑱-j��I�4�� �w=��3�茴�$TQғ1.d0�s�n��,����*<�e47R�ۑ
L�?g��~�~�/_N��ӓ��'C��
;�n�['ϡ��L�3<;�5KZ�JGq��
�w��ͣE��~l�q-�k7�y�R�.�����v߁��[��O�Co���>)�̠qq#�c��\�� �*�@6�Z��G�#�-Be�"�-���ɡ|>��]=G[b��cJO��;���_\:�V�z�u
;B\?ÄCRi��kY�1�a��)�TF=��9�?X��D+u9�S��d�V�!W���R�(jP���-&B҈�m��.U�kZ�d|�����Ͷ�\&�K�*n���hIi�u�R�ʤ���NFIm�¨��l5!a4�Ky�}dlt����)�,�LIV��d\�v3f��ۓT�U"�
��
pE8��e ���dJ����1c�F�c�����z������������%��͞��Lb�ۂ;6��C�o��MB&c�R_��c��#�U�Ł%k:���A�������0fK����v��|�x���|
��*|��?ß��g��羀��,,t��l6���*��Z��:�%�{v�U�rV ����FG�RVc.���]����]�����r=�o�L�g��A��7:ǅ��l�{�/���$��:d#)��S�辫��z^vojiC$���\0FF�\"ŝ$M����� wlY���>4���q�\�ҏ$�щY��^=W�AC�F�V�������o����e��ڌ;Y2ZɈ'�`��AK�at:��|:,fP�U����7��Ka��aQt���[�͆�9<EcB4����%eۗ-�oz��}At��1YK߳�f��>�c�|:��ܲi���"��I�:��F�H�X�q�]^�0���g���r�teJc�n��ǝB�~�X"��es��P���`��#Gy�fsI��]����ʿ���Vd�&�+gK"r��H��Y B�ڜɪ*�P �M�&|
��%�d6Y��r:�Z-F�6yzRh�2���W��7�3�}`��(�}�����:��T�q+�C)��F�| +�Q*у
��DF��x���kT�2�;r�4�]��ճ���K�D&QMOw��l�Cm4�P#�c��ڃ[0�7�W�~w޺����5�O�
�--�}�}x���a�q��{����q�ݣ�k�-X۶'N�FӲ�����
���Ļ.q4/�����z�����(��0���&�*�-V2dȲ�,)G�<8В��b˦l޲�O�F���t_��b8x����H7޸���!X��$�V��b UB�?���t5M����Aͩ#0%%��C�Tь�R����i3#�A�I�&���Ix�&ql��`��/��_��X�h$�`,5��9_%f�ӗ���p:17>{c��~^;~B�$i�vVD��qe6ՑN�z�V~����dxKZ�5�aL"�aӦuH�&��Tx���1��g��0=�CkF:GQ��ʆ:��q���F�:��*DgC8�?�h"�q-��Z��H�w[�RA��&�H]y����yQ�T�1��ʼ�J'T�GEG �A-��29LrvS��m�v�c��*�C�W�
~����L+Q��c_fF,1��8�F����'x�w&�G�hK5��ר�ka�ۖ�2)N��A,��Y���w,P�;��:u�T�{��x�y�?0R��Y�A�Kg�{]�ڎ(:�$��(�R��d��ˇ�Jb��<��K%�:̠(r�j��6w�to�28��ϟhp`�����M�dv��ڡN�Chq�p�m[0>����o�q�2�ho�p�t�n��Ͽ�P<���B��W��?p=g��Dkt��Q�>H�ܪ��0.�s�A��^W��"1�藿�W>�%|�+�������e���]9��y�����R��L��J���[�j
�IP� ���u��h�C#���Л4ؽk��KO���ϼ��d�'gB(�=%���W���C�,t߸@_+r��K�مl������>�@����O��wppż��w�J�ü��Gy��͛���gM���}e�K�����kpe`��c��6ܷ�V�x�4��nw�ۗcvh�f19�D2��NFS�w߸���s�X�j9�� ��X�_��*���nZ����X�18=�E���La`Ƌ*�'�" �dN�h���D��P[�Z��umMCu�?�h�']�榍����R���2������7<�¼C��=�/#ͷ�!f�+��5����}�@��~�s^�+���.�GNU�%�VE��!SIT�*+�.�[�� )� �!��4�}Y R���D:�\I���LΦ���rI!3��Z+E ���Q�A��Y�6����O;GFo~w?��>�'�r�>�����RQ�B�k7����2����4�[\9(�>t������d���N ]��OП��J&�G��6�>�s%F��lcJ�gO��_��ݠ��,�T1�
2#��+ob�����a�J/��5�܅.��$~��t��x���p�,y��o@� �飇��[�����|g�/��+g���=��g>�_���8��F�꥽x��=��׿�_=��bM��*�[�f
�"�&"� ��(���ػ� \UNQHw��q��)^=��
{���Q56�ƾn�z�mص��x#�љ98�0��FS���b�A)���m�q�Bas�JoP�睁B{ĥU�m�Z��/=]!��.�do&F'��5;w�.^�C�ߏ��)R�Qh�5%�d�Hkzo&O��a	�͊��.�j��~���5�k�a_�
� F�F�FU;w܈B�����Ջ�W1_���o���	�X
t�N�_�	�{�e�G�����S�Q���:d��y��ń$G�\պ��&�]^TS��-#^���P� =3{��H�~1�5_�-RIe��
�1��S����cD���� ��nL�uFc�ɐ>��#h�R�8R$�qU����f���6G'�K�ߒp�!��n�l��Xr{>��������,��
�b		R��T�<5�(@c��d4"B%��X3=8[��zOI#i�I,M�C��̚�s�*�_*��J�A����Q.�l�9�S?�lc�ȑ�2��Z�gr�D"�>�׷,���'�g���S��.	Gc�zO�&�͉"<I�:�Eâ%��]��(�����#&�&�i��׾�8��������\�cIKy�4�ў ���ݻ���&�E�A��?�}��j�]�E�(�Ͻ�����?��~��$SXT�!@��� b$��i���2Y��4]!���?�>��?B��ǽw���l�a`Ā�
g.���}
'/b��x�wQ����������9b��TjR��rm�Ak@��4�I���΅�P���}���0j�8{�]�~�V����Ak6>:��y��1h�s�W��W}s$Ġ�CK8�ˋƛe˗���Lq�#d���_����_� ���gQ\�"ɻ�w���]w!�b��;�݉��:�MbhxV�[�n��)�W_�қn���������0<�1�� �s��zg�hSK�y��8Y@0��j�%�����@��\�/0$~t�bċg�k�e���^��)�haQ�B�X��}�eFd Z���#�`@D�\��c��|���S�G?�Z�4��R�������F��a+�kӲ�b\�'��8��Bz,���2����������#�)�P�2�r*�������Ay<���̆H�_�����i{>(��ҥ	��Y}z��弢R��vpQa��� ����u:�"zP"EZ��T �G��#��GD��*Lg��ƫ2�\���1�O�(+WBn�����D��5�M���R���>�>{��d���)lZ��}��d�����˗�Ʈ���g���Ģ	���с�'O�w�Fu��l��H?��w����o����~�v��~�n|�k_��?�	F�14�kb`����m���V���0Ʀ�`�7Û������m[����;�։�2��%�����c0ND�李rԢ@�=S(BG ������+�P>ϴ�*�`s�eh�qb.M)Kϗ��I�O��������p�,�����u�q��b==M��ب"���@���Ӫ�רD�;��0	��0=1���Ehk��Ha��{�jY�/?p/�>x�4�n7���N�.[�g��HG�v!�����ԷcŒ�~3x��AӒv����xu�s�&��޴��b^L�+Ĺ]́�]���j%���l%�~��GO�6޿�%�:q,�G.F���l�鰗	�*��<lN#�5bБ� OB4M�m�[�+��S
b��<p0u"�����'kӑ���^�T*�������� ����I5�����g��E���*��CJ���o�S�٧��:��,��	^A=�ː�,"�N!	�E��$�a2��x8L�Tj��>95���C{�-C�s��b4ڳ�\L�Q��o��^�앹�l�9�<�c^�7(����|�ε�����"��Ub�E� �����F�PK��?�l�	�k�Q.����=si����A.�.C�x$���9�����@؏7�#�ib���O��+�m�Z<����OBFT��w߅����F�@ߊ�9L�ԃ��ځ���_a��w`��u�=��T@���K���O?���'x��_b.��NqN*b���a�1H��'0K����h������7���>���Kx�ͣ(jB�2@lx��F����WyH	�g�>�o*��"&�ifE�{h�{����é��7�Æ�Kq��א��czx�|�~�n�U�~x��������! ��&A����T�2�vg2D�D@!�!���%����B�C=���ٍ_8��/wu�V����q�8��^�N ���[w@[���a<�˧�y�*ܳ�V�階t�a��{q���0��(���'��8�W�Eg���q��Ȓq:�]�9>��s�\�)ʡVI�� �I��dX�N��H�X�!��Tj>���!�+�8���F��|TZ����Y���!�� �gҪ4*O80]������N�^۾�OGً��hO���8�F��G��U5>�1��D,�;�J�dUyJ#�|2��J&O(�H4J�[
�v�U��Cs~�c`���]�}��>8���U�vcZV�h&���y>�jgA�eq�0�a�k��,d���,\��+#�5�CĆ������K��[:�ob��O8`�؆�W�s�tV����Vk\���kr��_H���ؼ|����GN�MF^�-������A�)X�i#��/����:
'yK;�u�t��^�V���'	{�Z���A]U-���G���C�����\Օ.�W�:u*��A�V�9!������x��s�̛7L���<��IƀA���Y9����9T��
w�]]2��̀�z�O�U�uN���Z�Z{���C���͟܇����s_�?�T1�]�x,-
�b����b�>z
�ь��G�
2�CGN
����Z��w~���%�)����Z�\D�i�Py���sZ��iB��sgJ8�:�W�]�-W\H�h��C����9s0�Ƕ�O��փ�.������L�Zg01��4��hv��\�d:w�Ã��q���͛��jr��z:P�7������}Ȅ�DBx䑭��uƇo����O�r�:�^�ǏƎ�cւx�V�:yC�Z��1�?�=���|���M \��%ȕ
uIA2_�wL��hjo"S2f�J�7�t��M[�A\���s��3�d5+g"9�`E�2�AjN*I6���mR�9�<�.��5���b�t6E��zM�br�]I������w$�ET��-e����ee[Z-z}�T�N��7�)p�F�۝���2��?�/�R}�Dޠ�	`����4�$�yY�N��𸽢�+��J"n<y�cm___wKK�[F5��O�T���^D��!B��J{b����|	Z���VY��W�,T��4fhq3�� |��+�\��g��rf"���L:�����z��AF��]l-����r�/	��v=�ou}S2_4p�Z����_;�;(�_:o!���#t"���E����M��khn�GF�{_ߋi��X�d]#�����s���װ�y�.^�����G�`ޜ��;>�o��s����[�G)�q�-p͘��G�"J�4��(�U�qֲ�p��8�5ȦTd"I$�Qcؽ��f�F�0�_:�HR�B@��]'v�vr�Г��S��r=�b3�]�������!���\�v+��}���$K���s������p���D�WM�#hd����m�I ���a$�iV�"�K��(��E��nv:�F�8��-@�m���s�0Z����\�{6���C����o�g>�7��:t��c��Ch�97|�J{�{����k����|�q���d�ї��p�@'X?1	�h���.U�\������syc��E a�_x;�_�8t�!�LՓ=�%bt:�:�3r�I��A��J#g
*bLlx��L���)��l���iy͞Le\F�q}��RI��_�qUlb��Lp�L.:I�L���(bd2���[c
��Q�1�y�%Iћ��EM���x�d%#�:Z�D12Ѝ��dTM���NQV*��d����w�hg'��%8�I���7j0�h�b�O�;ӢXI�U��Ş�-�3펕m���/m��d-BEB�ۓ�t��V������o����"}v�/��k�N�$(���.٦��������8-�>���pxq��;��7}�ο����O��Y��j����������-���ۿ�?����� �͟���V��as��lG;������ي�x2#�d�J�h����^�#۷CcZ3�9#�(J*�����f�����Qr�/��@,}��?��A��i���0�b��H�C0���y��˼5@NSM =�$M�� ��n,�=3Z�V���hh$��b�ldE��b3.<,�uZ�4o½9�,,��kz#"�$�6�VT� ���Ż�U�'ػ�V�Z�i�� ��ю�p�Gqɚx��ݢcal܏����Ⱦ|��+q��^=.ZfWݰ��p5��u�J<��QtMDQ���d�F^:?r LN�B-�Z(%3����
FY�,��0X6?~���3���Ri���m��~PG}}�|�h�4-��U��do�f��е��B6�;��5	� b{�[
l� T�+Λ�x�T���k�Νt�a�!���VT��l*�J�v�M�����i���S5oS�������z}���j�`6��:#M4V�˩�P�l��pj��AmBx�#��H��1:>:�tGGˤv�[NL�i�(�1�J%���&�E�t$T��0-�r;c�а���5�$C�,p�3-ˌfz��
����c`iS��ˤ��p(4�����y+W��_,-�$�����Ѓ�|Q}����M��-o(���D�|hn��l��'0�v��(jx�W{�ѥ���~l<{��+��O<��?�i<��SX�z-j�.t�ߏݯ�u�U�i;���a��s�+.A�D
'G08\��p����0��	���������og�\��>u3��!���G�d���m$��ۼ�	F��_�L�Ձ` ,�XL��d�� �����\,
}:C̏��n��Fl���&��<-��n��ǰ뙝�5s���#���	Vm�����9^&���2����p8-� �bޤJ*�	��hW"�B^H�"�?����C�2�L,�DΏ�ӛ�7�c�����bɆ0��f<��q\y�&�k���ߴ�J�x� ^��������ʻ4�eh��U�.���;#��Tv�bBz�*.��W��d*��Nm1��  �#�Zr�^�˩7*�3���$U�H2�N��~]h0�t"sP�(T�4y�Tj������7��d��w���TS�X�~�Sl8������&�+Z�j�<���;��=���rz �)�
E������(Z�糈�C���p�"U�"#o�;PPÆt<�r������m�otX,Uy����"IZ`E٤H��ʄ�W�"V�H�'{�+=���_~/���� �s ��,�˟+�Y��1�Lշ��\2�ٹ��㒙�Q�+��(Z�sz��Ju��$���fݸߏ����j��N;���p4H 
p{<8|� ��܎��x�6n��훨kjF�@_��8^<z-K��Ʊ�'p��u}S[԰jn+��i�w��f)⯭F4��b��"�PU�Bl(���x��¼�̩�������'�Ķ�v!�*!洞���a:��5H��MVr�I�z�
�)�\�N�c�(���ji�s�r�|�yh�����W^A�����Ӹ����|��-2�(/���$4g96�P�sX�ز�FN=A?��^D"!�\�K�v]�%��D�q{��&p���gτ�N�b<LQ=9�,�_9�p��0���'�ō����������O|��x���x�D7,u��`�$6�1�,t������<#�k6�D��h*�@ �@@K�ta5��y�.x��獩x�H �)���G(2�M���m�x]:��h�L�se��#��b�Q�3ଥ�ՐIe�8��V�Π��Z.ȘΩ�BV~��7�9M�^D��9V�¨l-�p1T�)~�~.(���JS��7�)p�Gc#�i��v�;S���7���1�P���[x����IS�U��*
s�E�����雙p���@�d�F���i
9U����7�,) 9xn9��,�ڸ�d��$���>o/��B�L��\H%�*���k�l��ҩ�cphh�p ����#:����W=���W�C�����f'��k@O&����/���OLM���g����*�~��1<4��'�b�ri?�z�����UK0o��<rUU5HD���x���`�p�����D�]"�Bov0�5J�9r�ӠPD����{�;��9�,9A/����G�*<U�<T%���L(����b�i��%�(E0�$\��4W����ݢ}2� hC����7� �#:�}�C��I���L���L�;�L��E��dGV�K�Y�vLL�9��MN�V�%��y[M���Revu�G�p�B�^�;^|i�_�<���Z����~����7�r��"���<�����!��CWWd�Jd;��f�Ԕ��\�^��e�u%,�&(Z�Adĸ�N3���dM�Ѹ����<�]��kS5�0��KϽ�Kg2u:��ج�dqr���1\����
�1e2�L&u�����C.�3��+I:Y�f��E���T6+i͈�^2p�Ak�p6I�=�dw+5
��
��T��e-��M!�iL��w8xk��k̿w��'i&B����[_"��]\O����(��E��_W�:M�XG�s�92�t���n�ʷ"*����\i���
��G��EN&�U���_M'���&G��O�<E�\t�ؐO��0qL:N?�P̥�v�#jN"K`���Ψc�gty�k0��P��`df��#3J]]ݺY���+ߧ��t㵏��۴�}C�nl�cFO}:�����᪫/E 0�mO>
��ǖ����E���CB_(�K� �d���w�(�k?qs�/$?����<����z����J��L״s	�F=�-M�e9~=ܾ:�3��ދ�#�طgwvCr�'�ftZ����c ��� #S��C�N�`��K�� ��8�������������t�L�v����{{���p,ݍ\Q�F�& �l�%2�i:���Ȩ�i�-&3�h�U��٥�0�F�!�~rc�\�R��5� �$GA��\����b`l:W�輭	L��vDJ<���p�J�F����0k.����	��R�
�N�N\V:GrN%]�����ɑ8:�뭱�wl`Ȑ��5B��f��w�=�����7tS ��0����d2Ӥ(f��*׹�>�X��>;_
�E	��ת��&������z"ea7�;���M�I����P*X���;�GR&�Ϥ��ʒ�l�
p`����se ��5t�Dl�r��X�+�����1Œ��1���t�f���FFF�	We�I1�*d�t)pD8E$��=��x�iS���E�X<0���#�Oo��Zlٲ��;�����l^S,:��LPS�BP��hJ'�4�Uѣnw�`&G¤9��'�U���ip�з�V6#0C�Iς�yM���W'
�D4^540��;�؃�E��o���巖JC_�܍�~�d�u����aZkA_Tܵ�����S�Q�Dȩȸ�ӷcFC-�~��M��[n����+
���}�`{�Up�HE	Pѵ<q��}>j��7>��=Gq��-�ډh���l�Z� ]O��B��FD"Aܳ�y����̘���~Xk����`1�����fȉɠ9,4�����l
V-[�g��z{��cú�X�n��ك�/>�Nu��WEs@A���$��t�tȕɰn	4�+�ʅ]!�>�7.���~
8��#�Y12�&�Y��x<&�UH�\�Ja:����^|�֛�`�\̙��:��d�3m���I�	x����׬�g�O��F'F�'�a�����">��2�B��W���yD���<)���xKL��D\g�Eo)����9X0r2��� �o�1���?�Usj��甘؈[������;[�	F��L�s:����,�$1�W�*���l��F�a@�T��J����UU��f	%\���\�z�I�dnL�:��}c�XI2f�S<�5����0�֧[fN;�v����eSII����ȉ��D"��P�06�>2�n��Y_Peoǩ�%===u4��oU�X���i!��t��q��
�tߙ�C�\��eE#�x�/�A'��5r2��X� ��b(J,q&=�&�d��Q�J�#z�c``hI��O�`�?9&�&7^�ݶsW�cm_P��s�6��fua���F�cW_����o�'�z�5�`\�>47m���D ����zp��~\���ii�t��zp�Л��t�R�yA"#g��)Œ��VQ4����k�h8�$1.��z���B�[�ƒ��y ��E2�H��j��="�2�U��q�A24���7s�d{�p�K,D5oWԤD1k��Ğl�0�+���X��u�0���%Z=�3l�����u1g�tcF��)� X���)�Uf�T�"K���Ͻ��|�zr�N\�E8�=�*A[w>����Dk�����W\���a�Ͽ��v׽q��L8�324���tv:g �n�A/E�%r8L���kSy+���ȑ1GB���rY߉���L*��m.�bxm���7#5��F#�i�b�K�Pb­t:qFO�"��e}�yur���<q1(sq;��K1��-M=�X(�T�vKW��p&��3��w+H��E�J �X,�)L�tlU�#J�l~AU9M7�9xӘ��=���Fk|U��F��gS�&V���r�M_����#�̒��� ���E���z�?Yv��E�������Qe�T���C	��^��eF�@��b���OW�30����Em��S���\���g����d	��2���JdZ��dV���b$�T�+�`dF�@��`�4�x��I 3��xi{,u�v�t�_�u��ż����m�`#6/_���v!�,��L��$�ޱ�׭@��V|�_�\pn������0�u�\�QAGG'v=��7o��y��T�����.��͉��QrTE�Y(LĬ�V,^�`��a:M+�=�`���(Edv��v��͊���H��Q,h�����;�Ŋ��^~��ء��A�0<<���~�>Q2�ĩS����Hy�k-���5�L��0��Y��)jf����	aX�A��%�bΉ��@���̔^��KQDi��G_F6W��C'Q�CmC5�Ο�����GF�
kh�т9M��e2�`�1szb]���C��Gl/8l$r�I*�<m_��Xk����s�|�t�	4�`�Q���/������QFK���u��4���{}.��G��J QW鄪���h�X��
"��B��Q�Q``)D����8�� ������˼cO�\NUX)�����*�;p{v�&�,�j�t�4N�s��KF�9c4�L�_$����1��!-jN5�l����3�R�LV�F�Ӯ2�]iE1Ipz�js������W��z&��?p����+�fb�?��w�3y��3�R�<wJ�$*�X4����]��>wX�:�\tH��4�"3$�{���38p:�E�H�4��ǁ?t�� Rq�D���;�,0�܅�8���kL~��������Ou����枳v�y㚕�_=� �[���q��.Dba̜;��ux��;p����<�p�]p1�?���F�>|������˻�CӴj,X�m����m��g�Ñ���uTQ ��Oep��5X�d!�>���8p�0���a*P��:6�ǎ�>r�64�4���8�,��4E��}ݨ��������Z��G���������#(x6`�?�ӧ����#�_&�9���uB7��-|>�	0ɵl�+�_c�b�x���^E����	��ఛ	E��#�|l��r��ES}��Nx����q���uǑ� ���D���9{��jl" �Fkk+~|Ϗq�UWb�E����?M��5AA�Q(�!�?�H9��4G0m)��9B��$��U�=f�'�P�"'��\����3��W��J�]S]�EC~_6�6�v��b��|���(�n����L���3�2(��!{'�#9���I�J/�$7�h+$@�
^�w6����U5��d��|�`)�L�����q�+� 5��0��� G2HY�����1�4����88�{�!���e4��JR��U�:Z04Q̗�i�Y������	��)dn�	�>�M�O�����v��R����y��>�^ԍ�͛�\bg��3��\j�1G}�(E~��P���Nͦ'[yd���=�-��
��#"E/e�����eŲ�q�'��F�����6Mr4��r��1��0a��'�Ƿ�_��s��b�Q�G��H_/�Oo}���݀���?��5t�j����'����Wq�E�q�Go�/݊��.�/� �΅Z��sG�!���������`��
��=�86Ψ��/^x�5lܼ	7n���0��2d>�+�oA�Q�U�bl�.���(l��/$�Brb�~�1t|g�['��|N͛/�c�0�V�\H��Ң��
�ВVNTq��W8�����AG�<(�Css3��0�Ir��8�k�128�b٩��	��h;uJt>\��"�`p$,�N����G0k�,����ç0}�d�9z� �5����Ͻ�&�^��t�>3��q��A�-Nr0�\^`jzD���V�X�b�ymxKO/���&7)ӫ�4*��bN#0g�u��|s\��zy)�����.�x��СC����*��U���sCd����8ً$َ♀���P�u���N���  |�ɮ��z�߈!��c�P�IyI�N�9���.�u,1m<�i�K+��L�� ����u�A�5�\h5�4����0�\�������h��L�jQs�蹖�UY_�?�gxO�W]-��jj�0A�]�%��69z|���As��ǝw�Y��W���OdԴ�Q4�����Zn�N��#{�v�}�D<*�:��@S3���1Z���dr>v�E\ e�}�������ˁ`����g~ h�_�R�� a�x�U;Ju�����l_��/���~��oc�+/����Ɗ�K���8|��0f=��5�a���ןÝ�H��p��H%���x�՗0c�J�>{9~l;�:��u�1�ۍ�^'���k����|r�O�������cl` {�3K��K�ri
�tJ����QE���/Ƭ�ٿo�@�b@04���n���h����5�` ���U�B���I�梗�C� (�ܨ��q���ĬY��L�k	�.GG�D��χX<� =�PD��˕�F��������-ق˗b��xm�1��	��854��?���>t�5X����g��=��?�֯Z����|�j�w������ŵK���g^B$�f�AK���!� T&�"�b-k2�9�b�m�+�
9�reQp�
����bK"�7��r%_�sv�ț&���H�9	M+�J���(Ŭ��&����s�QM�:�.$UĖ�1W�ar�����+���+����O�{Ǚ�h$a'`�X&F�^qadNtE��T�:Ud�ҋ�Z�.4�K4'�6���$O��c
�c�_��������H:��
�\��T6�������9��F��^�6'���P<�9z��ٯn��,�bk�bqe��2�N��<R����\����3G��H���u�[A2p�A��*
-T�E�&N�qϺ D*���7J�cn0�(����pf|l���s����\�8j��O=������'?��'o��Ӎ��'����$3<<��Ͽ�"�,���"��6�_��n؂]�=���'�X�C�}2�D�(!+��|�9��b�?�
F�ؙ�3h����+7by�����6#,�<��~�����͟�>�����U<���p�֐öA�JB1�F�X{�Zܰi�XN��>2�y����}=������"���aQC�`Jm�^�p6��qd�^���`c�u`9C����O%2 �^�cp$ɿ粚�q�h�ϙ=S\���	T�T���^߇:�U�6�s6�cit���Ğ�>l��rl�h3���BV.Y���!��g/��K�CQM��t6�]��'1m�|�C��?~z�UMtO"P8
��%焂E�]�^pt������+���D{��H(fUȴ&�yU�To��?�s��(b{���A�{�E㳋���kJ8���Z����I��*V�x�ߪ�5x;Kl;�~�TXv�e%�:�,0��}���_��j-����ȒV%�Ӵ�27��L��0�9��D�����>�՘��`Ĺ�D���'h�͖$�Qd�BIdr�2m(��b��H��2������:�����׿��}���-��$�dj�Ntt��c:K�29L�5Zhbah��/��j����h��ٸ�	�V�/�9� �.XH�s���l!�!�ϭG���lfe-�F����=mR��=��P� aX��;~�����߽��?�|�E�o|�{Hø��+0w����lni§?�?��	������<��='��k�;�U73����y���qLol@jd��	l��,���Fv���	�K6�9X2�
�\
���[����+6����1�8Չ��*r�Y������ݯ�hS+l��v�م��Z-�W�f��C8y�$�Lh�/�'I�L��H0�!/
�\4��5v�###�����u��e�Qrlp9�E�]�Upׯ�CQ,]�[��CC���GD����}�^<����K`�>��z�.�z���r,[�/�|+�,�mDNoFdt5���n8�F\�e��5m��<z�C5o5r�̠�C�9�L:8gT#ɭ�t�jD�\`��d��h������1S$���+�u%Q[#�5I��:��-�c��Y���������skj~5
g7��R鄰l�x0�&oJϋ��!38୥�*��a����t�Y���H�� C1s�k�m+�7�≚��Y}f��A��N�8�C7�0+��Mf�2��L�-6k�b��'�ןsL��wi�Z8c|Wm�s��z���z��ad���­X��0�j�@]]�xN�GZV'N���m������/|��ܭw��I&r4���e�Qq��d��\F��9�����F��ș�hT��h�D�p8F��Y1��E;�P��#������Bo��	iMS���������]\�5������{~���?��Z��[o����o|Sw����j@��9��'n�����Q|������ Zq�g>�{}�6��u�������? GdG��?�ڊ�^|.Κ偔臤��m��^�Y����1�Bn|�kwb٦��j�\�?����j\���%�O~�S4��P=�h��x�>"���>w;dU��i9sd3ٸiQ�\�^���y�g�Q�Z���!��� �l��Ћ��F^G�]%d��084���	хsÖkp����o>��@/>	Ϣ��ַ~���~4�^���qt��\�|.��&X�!�%_��-8�;��/��a�y��-�($h;r�^~	�]s��u�u���Mߑ�#_�.�<&�E:��y=LF$�a0oGIg '��ROs�Y�
\Y�u""� �$6�cZ��}4�I}� Ah���T��A�b`e�{~��U���^١2��4U(1VT\�{u�i�����y���DF����^_b�ْ�Vb���2����;j�& ,'i��d&?��ğY9�<iܩ�-߼���Gt>�MB�%'ˆ� �;c
�{#�:sFoW��)�����fa�V�X,l�6B�?>��gd��T�0h�!B?e���ջb���u�y]�`v�+eT�1Z�Y�Y�K�ѡ���β���0<�5�v9D�a<��+����,������N�D�?(^�峂�#I6�+,K�t����kVxx���Sx�������>��������k�6ϜO��WL���wu3V,Ų%0����V2�k��>�Z�-3[q���W����n���_ɱ�`��*�E�ψ�[�KV�ª�A��p��Ɂ�(��ֺ�d>2��>�����l�EüذtV,��o�����g¸`v-�'?���]v�-���?Μţ�֥��pM�e��'��d�I�557 H�0�c��G�|�9�bm6�~:G�LZ����֨ӛ�vK��#Py\}��X<.�����`f�]����`?���� j��[�p2����}�c�Es��H����u�s�Ƞ�tۯp���1�y_y�^z�Y0��Al�V����C��f�`��gw�k�N�RLH�����rKf<%��d�Z6' +Zr5}6���%Y��M���yr�����svi�!����n����JE��j��x5�*oQ��g�ފ��)T�+m��*�s��"Z7���[�z��Y\,�?K8Ï`2*Z�H��50��1�d0�6�cp�$ ��-ݦ3�,���g>���X�4���;c
�K��϶����틄"�S��� (�˕���gR��8jsz"�˵c�d�2J0��o߾�}�w��w��rv}��R����m��iL%���]W,�!����%�逋P<k;LL�D�A/@��9{���"
9��v{	]3g?����}F��J�:]^�����ή���b���I��;n�u����~翮���_�������/���ɏ�z�|��W�C[>����{��+�����F4͜���3�Bx)�	Oc�ׄ�]�kZ�h�bC��Y[�Of�[ڹTS-�� ���]3�	F�Q4~�ea�����O?��	s۟~
3gLìi306<"���`S�p"&���f����L�7�ֈz�@8$  ���wv���Uhpd�#`2��d�+���S"��վ*�CqA@��X[Zg4
q1+��M�a8p������3�����$d��t��^z��Vl>����2iH55j��r�b:�o}�h�7^���A�k/���Vc��V���Z�h^6�6��w��c'�wzQ��J��[�	��c#�s:0CG��2�8����a��dVE�l���|$uA�=���K�?�s��16���3�VY6����=�|����Pd�����a�Wa��$�d�9\~��8�H^�MF�|r��[-�E�1�r4�ˊQ�c��F^˞yb�`�ʓ���(�<d!	��2J��~owL��wq�O���L;66>�KF����"
^���0j�C�����jF}mF�ǹ���ek�;v�ᶶ����Xuu����<�=�Ne�^�b40�x�ذX�(��"b��f3�f�,65�B"�l�J��
G��X]d��昐�6R�,	��P� N�|��L$[:N�l^���ᭅ�`�e2=�ⱻ�{(�����'6]sբ��S�.�p�f'΋�����������������߿�-�V8�r�1���O]{.5Z�d&������b��9�Ӂ��C&�c%���O�­�ݎ�d�{L �{�`^m5"��Чb����6�tvvb��FMB2;����謭!Z[i.��0674��<6�ӦM��Аh?dc.�G��M�A4���؄�4�=>D��rK(��K�b�E�ɧ����s��@�ϓ;^��R�y��bչ��l�F<��M�����x�k<������B������p���;��c�?�x���VȺ�\y�r��h>����.��i�r���F����4-@�ZWa~]�;p}���a���:̓EP����sy�p'w=0��L��zR���)6��_��q͍��3@�M�j.�L�H�d���V�DݑRQT�N\��[�z��>��p�
�S�Z� 
?��P�Ken�͛BL�S�����6ȣw�̖ɪ.�ͥ��e��l��k��Ѐ�sa-Z�]�m��Ť����Θ��I�fp��S�N�8l�Z�5ը�:���r،�������h���lƘ��9r(��ة��mmmc,������o���΁�'����f�h5��r��XU��� o#��@s{/X�_��XTQ�ɂ4Ei�by��������DT6(t�/	T��F_�D-������|$b������Ҙ,R�}�'�����=���-�,Սr�p ߼�A|���в��/���1
�Gw?��Pf9�b6��&�t��j��Q�!�U��^��P����6y���ۉp�@c2����á����Ǒ���2Kxe�!�v�a.���B1��t
W+׈(6��i���!o�O�0�/�	��7��G��]v�P�.w�
]-נ��[!�K�qVf��s|������at�{��M^��SϾ��V�D� ��cd�:1M�������*��REs�-X�~=���v�JE�'͆�e"ǔ+A��㦫.���8��KX�dj�n	�pׅ�i�k`b-Rd1�e	˧��dN+�k}���F`���V�&�0Y�3C(�s�A(�&�����#�|��[�h�&���ϸ��mOeQ��>17އ �����5�l��ֿ���� ���g���íl+0FE��'�<�ʝ-
}v�WJ�?�������k6����N��?�/���tu-<��0�'���P�s��.eC�d����6�1���]�sSs[��$SΌ��
��`L��/�l���bW̂@�9�d�cل\(�Ou�\��>ƌ��xM._�f5w�r�Rr4V���Xk2]�N����C��EQ���+h�3�g��柘@��^�?��9aJ��Ġ	�Io�!��u�V�����G��}/i-�՘c�'>�dJ-Z���|����I3����>��7��i�uB*�`��躰m	U^�rV��@��#G��PDA�%8v����)\)�Quv2��u��1��}�>���A�DV��n�p`��^,�֌�G���/��a�o+Z[g"�L
�ƺ�F���:Ud�U�uFCЛY�QC2C��Z�&0X��D6�|�Y8�A%���*�<W��U�e��o|����X�f9n��r;Չh,	�х��!�b�p4��գ�!׷"U*�*�����D]N�-��N��:�μ���1���M��J��\��⋱vVbCX�`!�j(*L���
(v�hΫZ��ݡ+��J^�s��j��|��׻���c�a��`�s�T�.3�*�7:��]>��d:&��v\&��p�{xF*�]�؎�c���<7�/s�2�_j�����ݪh��E��e�m`�� �������f���Q.�XMV�%��
�Z�BDi����^��I�|��1<<l��;�3	�N�QV��E�� Zx�
�%�PV��4����{���wcL��wy���2��[�v��j�M��L:aΩ�N���MD+�Q��3�@mm=�F����x}�#�.{Ou��:x������H9�Ju�a���G6�yW���X(����r�(Ōf�$��:]6��gR83�A�����C�?�t*��Ez���8��w�#�m�DF8!l�F^ 2�jɜΨ�;:Z�:�>�Z��������;?N���꬚�5��H\70J�5W���K>�v}�])ֵ�aJ3�a�R_�=X�"�jy�=O �`��
t"�$窅��}��m=~��f�J���r���h���0�yp+n��*(�,Z��G`qXE{����0"3ę$�`��w��&`b&2b� .4U	|8�>;]L�a�XQ���ŉ,�[�K��޾X�N��w[a41���/��^?�α�Qh�̾&��y�^� �78�y��?ϲ%X�j#2!���`����p7E�z:f.0��.لKV-á]�c����� B��X,�b.��h�-3�J&r����|�����p�?ց�}cP���{(�<6�5́��4̜-`�NCӽ�ϰX����N��J��;��x��?}�W�Z�Ƕё�x��@�-�-"P�X�iem��������ʛd�*<)<��̞�Θ�z��2Dف�|�1YDM��4k4}�o;C�����z�LS֡�n,ޮ�r��/�`�1>��(�K!M�D+Y�f��q�'yZ��c
�˃���چz�sJ�ck�Q��`0�،Z���P6��YN�C��m�	��oUlU���A���38�lբ���cC��Xw޹E�ħ�n���_z�����Jz2�攧LW�!�1�k�l&��a$@�7Xɠ:�Q�(J4��xh:-E���E���C�)��k9�0/gA���A��j�ztt|a��=\'��l\P�@���߽�W��Ӄ�T\Us#:�b�Xt��(�w�a*f�������8s�T��dS*0r��E4Y2�F��fBN��}�Q�<
9	�o�Q��Y.�˖4wt�;�K����)��IFȱSl������BV B� (j� �Y�39��EĊ�f�q����`o/|�tOe����G��b4`��٘9g!�}q7�F�h{����6\�K�"�1w�R��?{�T���*ͯP8Y����8g���/���x}C'��箘��/���+Vc�9���vԐ�^<�Z*	E��a�B�:W~����
`j�Ds��3��B6O��j�2,A��/I�J-e����	���"�d���T�R>M`�
)�hBtBd���Rm�q��w֣�^�C�2�~a���m=��$������9�DX�M%nafFU�1�ɭFv�L��s��B����ذ(M�rG�LD��#���Q�LjQ0�Vk�ju���"����;�����t�"T&���r�3/��d-�"�d���gL&�G��t-��;����a̟ߘl��r`db��j�Ւ15X�8h��3�"�,M�X$L�P �u�d����AU-�Ʉ^��ݽC+�{{_,m��m��{Q��SS�(��yv�b���Lh9-;F�1�N���DF�5\N;N�]!���e��ba�C~x�^#�6+L��yߐ�C�Џ�˪jd/�I�l�pha���Cp0I��Ǉ�{�;�\>9����yv(69�N$�t��z��������\5;`v�b�D�۟�%�,-=���A�����'�w�&\��!��đ!�o��p3�7r����?N�X��t\���g0�³\���y&��vE��*�e/��rʘ����=e2�i����*2�Q�"~���O�w�a��������у	b糯���V��'���� c��,�0k¡2y���D�l���F�şL�P(`�� �y
�+,n)�8<r�,�	�H��bf�k�-C&E*!�$����N�#�J��Y�<>�	p� �(��Q��Պs�77O��j���#C�Bʹ�#���E�;B�A�s!9>7��|.��gir(V��\J���k��Nx_�������|F.���z��9�9�&p�Jf��H��56r�@��	���t��I��eGD����CYcA/��8��$�B����$�h�MYs����6gry�Dюl�uBSC�ŕ&Ϸ�	�����y=pF-M�� N�@z�ј��+q��1��)W_�����ԱT:�8�+ҥE� ��8�'#9����A��C�׃��E�J�����y}�Y+V������|��},]k����Й@Y��".���n܉P�T����PS������J�l=�|>ܲ�k�Q��ǙD�D4�"�D�/w~��)������H$:�����J���X����Ri��w��ط�/w�{�j��Y�H�4c~+>���8���a���`3�ۥ��Z�H�ƃ�g~r��k���oN��q�C��ߏ�k�E>����\{����/�F8L�-�E���դGJ��a���K�t�ăA��ݼ��`-��%pȎ_����oH�P����7�X*t.z��煦���qr7K��?D&�}�݃M�\��j7ο�_�G�V���(:bx�C�O��7��R׌��Dߝŏ4�Ę�D�3����>��_�qﶧ0ͨ����PE`��΁u$\�u8�� 75��5�˂Q):G��u^�~�Ȁ�"���jo��Np�*��8�$9u9�D^{�׸q��%�� O4�uf2yH����7&]��J��,m�p"�f`���d,��&�7�g<�5M�Zł�d*�V�xU:J(�V�8*[
�;����N勺��bE~��tˢ͐kt(��R)]�m-.������Ρ���Q�OO�'k!
����L˔�:~S�T�d��<��*����)p�g�/�4ֿ�r$9�f����P6���8��w.�1���UOQ�n�n���Š���G�:֟��ľ�wE���k�;FG�iU�H62��"&��H ����'cqXl(��}d��� C&��PI�ztl�h�"�r1���*�\4��`�4)*U�V��H����X�o߾#tZq�ǖr���K���_���{t��R�a���Vf�<z�7�?�#��xo?�ͮ��%c|�Odj�SW�����t�����y��+o��kףm(���|����9�Arr�׬C$���_��e���R� e{w/�x6�?��LO�L�\o�F�$�tAT�Wl��վ�頑��y��@��i�\�-|N���(���)<��e�'~뭟E�׬��̂P��@V��C(���ֵB3[E���ea�9���wѹ	T��!�BY�Y�=n�@�:њ�ŬR=j�sr��@X:���aR�pҼS��� ���1��n�eg�u;F�yVCu8��B�2��܆z�^\�f���w��]��J�&�ۢ��B9�^0E�z�v�F뗀�NM곩=W_un�����_|<`�'Ͳ$;�JYU��k�B=#~si���3 �;�3aȶ�{8�����:(�
��l���keE�r׀��N�$��\���`u�X���-|���W�0���փb��.	@S�k6�-�pXc��wL��?Ө�Bj��%�{���8����D�*HBXV�S��QN�0::���0��Îx���uZ�b	�+�ߵk�dD��U���&���N�T���22�HQ ��e��X2!����9z��Pp:t��͈E�uy! �-��n��\dHMh���s�^��2�	���&E��g�#��[�><*[�/��Ŀ}���ᱛ_x��ւ޼r�y����6��k��P��Q�jfPD�ENo+���kq�c��d�0.���ܫ����g^yW�p#�>�R=]ؼd6S�>�@��4��n��6��P��瞃ݒ�����JgR���X�V'_����+w2C\�R��a�fr
fB��������_F����������;�:m:6n܄�?�ކY��Cې3ۑ��Hq��Z>�����b@>��t��_s��hÃ���X�5�c1����
c0վ��.���-���~+W�G$�$K%�BZv4L�\9}������n4�6��������j���	 11��
sI��������z��P�w���Xk�����~	��ixk�p@.���rɂY_1����wn>g�����`�֭R(���ff��l�기U%�ǀ� s��3�&[�+ʋ�x3���L��6�dDf��#O�VE�jP�
9޳ &���Ga���/���V�$}`�,U�	 pAbnR��� Wt���D���Z�]6�sjK��)p�g��������{*���1SS�:��t\�d��a,p�@�hV2D5>'9f/-$�QKF�7��g�-;�m;@;���ٲeK��;�������յ��,�)���!�[�_�t\�u.��9�{G/@��b�(�R�j��.�*��=/��n�s�nn^V���&m�����Y�v�Df0�ϙ>o�0��+[�ߍ�'�_�D;s0����v�>5ECtF���6-Md\�nX-e2��]ȦT���E`2��3H�a՛����&m�l�2�$;Y΂��P���d�gtl�����~̈́�Ga�e5��W>�Ԗ���<ߵ�魽_��Mf�^���+�bq�?9ы S�+�=�	'���ѱ`{�)���a|폿��ݽ�o��n��n'���3۱l�R��������^K��d ���!l��*\{�����Q����"��?g1��H��	��̳$�7��[��⨨$h	 ��u�V�ի�	�O�Ε0<9)��_}�]�t�Kc)�jx��K�}��L�le���R:��� �4��q�B2a|��k��v��?ݎ"+*�Ϟ���^��H)0L͠����"���ݻ�r�:,6�����|7�,�ZUƩsH�"�(I�k.��A�"RɑpT�N�Y�v�	:rV'��ᠯ�*a�	LK�h��Rc�d�P\�D`چN��2vnx�봽tӆ�?{����}�����t�_��]���:���7�S��~��x�ad��Z� �)fM�˹si�>�ȋ�A}t�^v����u�r�9�Vɴ}��tjp��D�5j��^K��;$��dke��VR�=�����Lg�*��N�?�vS�[�����jnn�>��;g|��3f��%���J��ei̗D�vzj\4
Z	 x�vxD���ʖ�Xb�;��^B?t�{4&655g[��B�P���SC��6��"�D!k(0�o"��� �D>�ˎt""T3t��P�F��m�٤��dbL|�3ٴ�q��-St*�j�<cLơqb|r�a�$��G:]W��n�?=�CS��|���{����KՒtx�;��o�5P���y��05��_��C�`�:;E@ъQr�+/ۈ	�4h��k�r�􌆇Σ�q�M�p�}w�����ϼ�X��Oܼ	+7����'�	��"eU�(�����pnU�
j���������	 �z�!4:L>����t-F�a4�w`�â4�����^���l��ðhr
]YOƿB ���r�6>w�f�ȏ�h�cC_�7\�'��Í� 9�t!��o&�\��������Gp���"��"@���;{�W�9'��i�t4wu�L��f�#RL��D�����M]�xg�^��s 9��*9,9*M��j���4&ud��L���-P����/���^�n`�GL�)>7��VN�۳#eG��w�$KdfE��_�Bz�Re�xlp��@˄Cz��g��X��`�k���b0��[�\���
<]���J1�g�8���q�߯h8� @��d��S���(y�2JE��������o.s�k�8�^+��ٹk�>%�\��E̘�,l�2#n>h��g�}`y��A8dO�3��_]YI7��a�LQ���9��J���2�'�Ѯ�J�V�H� �C��C7)j�1B�
Td<�v�NBA��z�r"{��Fəit���	p`��j�*n1+	�6
����t��������g�0[�G��b������i��ơ���g��<p��+9��G�ѳU!��Wm�h4�W�z��l���<�g�M������;1<<��_}-�-�GP^��֯�?̆��Ù��:�a(8��/��n�&���}g�?Zh�X�&Ak[�ȘS"��f����BC���3=�P�/��$>�E�<xܝX�f5�^?B�4����?�2f"�d�� �j�)�`�	̒�r����;�yr�F-�a��W���ۮ^�v�CNo@٠����?~�<��6D"�����u��j��H$c�e�-�af%E�e�{�L*A�ƆT:F�1o[� l�X�Œ���!Q��Ż;��Q�@��	�g"0Z\t2eA��zL�t��d���#�_��՗?����?j���������P�G���(�V�s���|�4)����W��� @4ʚ�zIa���� ��f�W��)d[>,׀415�TU�z�Qs�|A{�GqyT�š��3b=[���~�f��M� >"�&�k���^K|ٲ�v�^k4�=�TB�T��LZ�n%m�����F��腑�5��q8s�mxll���G�oݺu��w��o�k�������7d�����ۛ�rV2ku6��V��^(F�1��y�y^�Ƅg C����K�kr�y��џ�r91���b� ��,�!K����`���x�kbb�����߅�>�b-�����g������g���=��sMw�t�v�U�pt����g����*���14@Py��OCEf����_�Ξ=�W^{]�RjZT�E�Sl�9i]Xy�F<��+x��W&�Q��!W�832�m�?�O��p�F�wPd��<N�4z _F������k��E'?� hbi�<$(��g�ln�L&�g_�sCL�8��`�M7�lk�o�o&�<��u2��w�g�U�z�d��f-&����G�@�C��67�'���U�V.��O��{�V ��X]���;,�6�[���\U�
&�F^y%�Ĉ 3p� F&�%�ZE:Gy�6�A�"`˒���t�3'0o�<x�]H�u�r-�xi����?Ad�R���˾���_��z��>�࿺N�:���l#�٩�M Tb��}G�
؎�3���O�G�Z<:�
�K��l�����h߱�f����h�	��d�:-i�*�߱c�j|x�E-kd��4�X/�5����uh�G��kr{C�\.h��1���cF��k�/v�{��9s���=��c��dt��"�z�H�&:��bA���傣�Y�2�=S���YMUIv8t������������N�g"3�����|�(�x���ȺXA2]S೓!Ցq�&/�ۅp`FD)Q�C��ҩ�14���0��z�;�%2Un��$�=U�șt����/$�å���yl�j��_�����3O���?b�O����o�\s��/�����C���ϟ�tP���'G|��|���v�:�y�<��Yt���3�o6��Q�x2�S��!E�m���g��9�K���e��>L�?���?��>~V�]����9��ɂ�
E��TU�v	���TAw�<�t���DF;��^�Q���O~��qR:�{���GNK�ی\2��y͂3�{:^�����a6�	�f�2�pjʇ��4F�L�|�rA�m��Xg��8�-������羀������/�?}�A���I����%� P����c����ʉi�*9�t�rAt��闵:3�n3�.�/E*6��N�l���!^|���m/`��QH�r�N�ߢ)���C�=�����G�*i��Hs6�m"��f�^s��\����6#�R�X�@�\_�3i
@��ʈ�_id[�?O�/�u���`�P�@��Xb��Y���Lf5g����.wps)b�L*J%JA��W*՜�`om��0�~���uي���=ǒ��H�`�+٬�L�]��Q֐1K!
#DN�J �nv�����A�"1B�r�=2:�n����_~��7n�����<��y=�����r��:O����B�D�E!�*�)�p7{av:)J2��!�r�!��g����Q̟?-�z����:��PmbB'���
 s���/���o�Ex���"������3������oE%��M�/jQ47"��`�-8|�<��?|��p�H?::�@o���=N1��͌)n����f+\�����45c~�2�v;��.3:���=����$=o=���A�3E�\��T��S�2@f�N�΄౹KeD���;o��{�BF�B�,�"@�6�l���=�`l邽��Shj���]����ba�r�~��رg?��4 ��qI� 06������נ�aM�Vu�[���W]�	iO6�=�o�Y��i5�{��y(�b
]�(������#s7���ׄ�@ ��B���nT)�\���Èc����p.�]."������C�o�]��|l��h��z���n|b󥗜��^�Ą=�Pt�Z����ld_s�*�BS!˶8k��Zpp ����d'�B�����K�>J�h��P�m�W>W(��6�V��P���S�D&����L���=��2�12��	VF4v ���-�T�JA�B_���~d���w�9p�Y�+W�E��KQ̞B� ������5$�/DT� �`S[߽��D� B1�V���=��%����6��)1n���~�g�;��J*Q,�M��z �!�ɡW�%!�ÍF,�dv�D6��t�h2!�NA�Ո�a0A �����D�MD
ܼ%R���,�N���TUk�t�>��H7�c�b(-�����L"��T:%���|8�^�YdIo��h����XI:����������C�;�� zBx�%W��iw	#�����s���L��4�����@7l�
��/�sϾ�G~�|�a,�H��>�y�tA��"dQ�g& Z �#c���݈�s�����؄�n�Ͽ����
��O���!�~�:��D����$,L�E�iz���	�̇*��7��9|���ǎ��PYК�(W�0�qn���lX��n+�z�'�&�/_���T�1�	�,^ЅӃ'���@Q�F៚�s���ϊ�����w*�h��5��J��<W"��*�&��ܞ&�����XF����y��=��AR�8y<�-7������>����o��ڳe`�����w;r���"i#�ꍆ)z�G�.w\�*"3�\�ʙ^l'���z��	�l3"_��G}��ސȶcV�3���d���57#~���ԤV���Z���ɤX�Z��~=�T`.�%�\��3�&�5kj�hl�o�����`�����3=���7蕼]Q"Z�-���	�2�}4���3E�M��"z���Te�욘�]v�ԉ�;�m�f���].�2�����cG��Ҡe^:$����H��e�����(�Y�V�7���XL�!�ry1��`!��Z�����l����aVfG�0+��2Ωd�mdr�����GH��,~��T�C�O��oӜ�+7,��TA�k�(�҈���y���Qd$g�r���
�A�D��a�?0��L`f���� ,N7���82�9e̿d	��Ե��<�����/_�'�_�D)���f@F)�sԣ��Y4�MNL��5`���v4ѽ��:�������z�#�q�$z�	ir�XDt��fX�ف�=�PSD_�G=�o~�a$�Ə�S�B��UŲ
FG3��$F&|P��_��}]�[͢P��(a	��-MN��t���=ܓS)q�@#�
r �4g�U�Q��|��5ƽ�G2B�B{��};�9h��f&��7\��#����E���r6��܋��s��/�r��sma`��W^�g|Y%�i4�u�ԋ�Z�?����.��Lu�"~ok%�������>acxB�@��#uvj2��0��7�R�j�Rɚ̖@�������w�^�������0��3�B��R�+|O�ɕ�3�&3[���)j$�p���Es͈�q́���jjBn��KN�9u�(E֋I;*��T�hF���m��x$��IQ��6�.�mmm��O#<�hJ�J���G�Z��{l˖-��qa����s==�>q�L:��Y�fQ�#� ώO�X[�"!��t��b)@��C��42��`T,�k ��v"���)Rt��B�5A��M�*����seV�UɅb���cc1.<^t�Bܤ8X����r�㏾�+{z:t����Q"ɦ�����Չ,9�bI��Ͽ�/m�7��	<�ݿG���H_�FWJ�7z��f���*��jh��p��aǡ�h&��u�)v@"�8D �y_�җ`!�}t�n$8�C���X�z%��G�,!�/(L��w��n��W�CsK;d���F���벢l4!G��/�{��`s�ڵ��	L�P,�����.]ډh"��Lz�tF����~��6��k�f��z)�k����BK@�L����E!�:����˪��t"�S�3�fDfEIB�Rc�˱��d0 �~G�2��\�YgBCs�]Kb��b(	��k�k�N�S�����Gl*�V:]u$ҩ��|�M�@����z�6��A��A�Z�{��Q��ɋD-�3gt�>0 ������c��ߗ.dxR�R�R��0�����s��i��0��&~=i6�%�j2���k��*� <�r9��'��s�
�����hqDV�z�C���=��Hj�&���p8��D��a�8D��N�=G{�H�l�2==�����u߼y�22�@a˖'g���wL��_n(�����ғ㖵z�3@r��(���=��=]���B�@�WQ:(�q�mGcYdL&,6��[�w2ƒ�,�ƻD6��F�#S^���G�I�ìŒT���m��?��+�����U��w�CN�{�VQ�k��"�D���q�����C���M��)�ew�;����Z��Nap�W�	�^�B	�����w�%���"	���u;n�r#9�r�:�v!n5[����Ǎgq��	�%l��۴�X�T�'�o�T @Qz���G���b�,�:؁DI�hOME�8x��Z� V�����s��`�b}_����{á�	U�j!�VW^�	v�);F�V�Z�Ls�
��<��#�d�D5g٘Z�y��	R%�f���4\' ��erB�2RRUW�8>8����tva&���nA� ��d.��3��ǎ�4ڌ�7]���� x��]�Tv=O���d�jA������VAݹ��ujb�<]œM��4>�� ��z#"g���ϓ
*Y6�1`��\
��/�Q�n�^o�������c�&1��0�{}*����h����bnnn_�v�ì9p�;\d��<}��a%��ţf�l�M֩a4X�TRH�ፅ#�64	�"�.0YQ<��t:�.�-GN��q��e,�|�߾��tw����SC�rI�Q�j���c����+�'�(:0I�d�4���&����Hf��'�J�H��V;,��!	�}bD�9D�5�̳��%]4�虞�l��E��/�
\bx�t��?��v[�R���ӵ�u"��@�x9S������1,h��_�2bScx�{�z�����p�݂�H��;���ܵ]�qp`�8��ƈgl.�Ke�	4��O������DR����!`�|I�-Y ٮi�q}�`o�=��H'ǦuV�㇚W��!��|yA���ir���}�-�:r�Z<h�����?�a�V�(�!�3��~n�������H&B�L�!�`�	�Ԧ�q�B^�2�i?qt�dr����`0�tj09=#�U���&��E���Kd��4:Z��$�)�^��z��z/+�V��#{�ކ'֯_����h2]3>_C:�mרuZ�q�Ι�d2.��-by�j��H-k��2g��}��gΜNX��	%W�*�4ÅkhĴ����(o�bD2�NLݨ�`
}�[R���}�y�޽���y�*5ʲA�A����i3O�B6�{���Z���6Q�f����6ό�f�X0G~�>k�#ՙ�����G_Ng�c�xo1��XMN��K�Ҧ�4##�pz\�W�j֑1mC(�#�b��25[�{��+��Γ�?��O]h�����m���ָ/��u�&��/K*�b,�Ќ�˕<re�g��q���L�|��V�]��H�J�P��w����l�a�&s��9���u޹<BF]��	�k5�R�ub|�yjj���G�J���<�wZ�}��?y�|&8q����5S-��YVZԡL�k��%��?�2<r��t|�/��?�����'�id��8WK��*-J��F85<��5W�{��;���wӳ #�4)V�4A�&�6p'����dC������6n�a�y91�	r�i	�)n<c�D�.$��ΐ����X,2scb�z���聓����X���ڀ��v�� �{01:����4�HĦň���4�CB��`d2%r��H�@��pZ���4�����$�,�����W����N�"W�vi�r3��ާ�6x�͂�d��IVW+�J�ر�o���ww/�O�࢙�y��L�����Jn�5z�<�A�U[��j�xչ��s�
��^1�@��f�/,�V{�)5��%��i�T&Q��2
=c�-�A��N���;��fkq�ɠ�ӳ�g��e��Y9r�
fx�*�d�'2%����֡���9%��Ys��w���k�<4<2����l��dl<v#�ِYb��t+�k'&Ǡ3��6PĮCs[�@�c㪬��>s��uKO��u��ÿJ��5YR���w���}��֚�&�6G�\����"�=�3�8r�$�8z���Ņtn*[�k���`|�Lb�"L,Tó�*���(���ɸrC#�r1�wFC���䤓ni�O1$��'�~����ăVwKK�,sI�����n������������h�#-��Xv%Y��V������/��P�l7]{5V�^���v�W�lē/�����9E��ңq��>����>v�*e_{�h�\����C4�}���Ĩ�����>PECش�:\�z���&��m�D�P��i�H3�<Do�<r$9�y���c�ؕ�bå����E.������?��AԳe1�I��3�'r��'7رT���Q,dɷk���c�Z#��݅:97*��F4:<�9=�:hې�(�T�J��N�Z������z���*�����1W2�Z�N+��v�D�H8nN�s!�����?��M�Wx��P�/H��B����#gu�p��Z*�4���U��Bp.��n���l�1�>P��������hy�TZ���-��X�j-���~�hk@D�\ӫ�R�IW鵳z�~����1MQ��k��ҥk"�{)�ɮ�C�X��e����������hhl��&q�(�A,Ì�O�bE�����wӽ=�|u��Ɍ(ݽ��9|�o�V���E���F�g~+U��,���x�F�n������K��O�He�$[9��7	�1۽̅~u��N�N��LO4����D� ��Z�|��mO<��f"�ˠ6t�t9����|#��X��E���4�-��������x|4�/�����_���?�D|w|�ftw6�_<���L�:��+�#AQ�ַ"_���bF$��J���܃���m?:?������~]��U�(s��w�ь�
���u���MP�y�x�yGaq8�f�)�{���9�y���,��Coo/�<Pq�,�a��,v<���Eq
J&�l*-"N���A]���Zx?��Kg�5*_��T/t�3 �n��pV�N7k�J�5Oc#�ѦϜ;�V0�ފ+����]T��UO=9OVI���*��}�P~���s"�/d�UbYd�}n&pp���]�,���$��>�qG=E�&���?+�v"�.�*u�iw�y�I_��~��S�H���쐤�i�~L�R+�
~	6��^�(F��vk8�>m�n�+)|�5~��Yʾ�扣��{lG+4g6���tഌvKQ3���4��/8<2ɔp�Vr�ұ1�  ��IDATg�}����C�'�ti1TkL|d���{���ck3��Y��5<}��h&&�qwoUbD�o
o�t��&�Y�2�$�w�"���� ����G�0X-���k�m̡�EU�ե2�����&����F�k1Q�`�zFg0>��S�UGB�{T6GgQ�J����i�x[������=��;�z�p`�.��g���X��
�{l C�Ӹu�ͰPd�¶�x��{�r�J���Yl��R����t�̌Nr�X����s)����W����/�x�ŗp|�<*"y?�n����}ظj)2*� �z�Z�lw��(�C�p��Hs�H�8�
�P�(}���X�b	�N� 9RE`d��FT�"�e�lN8���ħ�kڙ�`?�� ������W&���v]��x�Ke�a� �������*3e/9/������g�F�(y�����.s$YI�v�a1�PoR�gPg>���B%]�P�lb�����L���S
���T;d@WSz��U�w<�.�4�q��5ɲ��w��m��G���,4�MN<�PEi��)/�88a�6���d���Ȃ���tccù>��#=���ḱ���Z�h�����;�ĥ�BђW��P��G��W��F"!LOM���&��ys:/K�7�7h��B���Gonln!P0D��3�3���C�Nf�I��������4_.����5��!8��6��dFLh�(JS�䈎�8e'�/P)����5�̆[�C��}"ԅ|�qrzb���җ�[b������ǟ�������&&�MT�ض�6�z#^?;��م��Z�����)N>��7\��{�b�у���k��ra�K���u���S����� *7T� ��i�K�2����"�<�Q4���]hp8p�'�B�t�%8=z�����۸��p%FN@IDp��WѶp���>�]��Ǝ��AU��-��f+.�l#F�(%HܶZfv�
��I�os#k��7��^��A�R��,}���jxw��>�5S��[-�ck5�`�/�n9n�-N�T윜�g�屩�?|�T�<�jժ�t�.F`��dښ�d{�l���Z�)~L��ɦ��ag�#��Ě6A�=���E�p3��dο65PN�*��B0���,�đ~*��R��5Y��v�g潔f���;zb1��^
`�h$�\��tN/d�D�b1q3"�ʨ��}��xod�z����f&��h{�>̚����岍kO�>sf:�����t*&R�ܱ�Z0�qd��D�:�$�-V467#�#�W���,c>�e'O�|ݕ~�:�o}��_�ű�oþ)��r���J]&��I��42ǔD��`�9)d�%d
�������H���̃�4+�D��k�2�b�$f-�X���J�r��%�H.��Fl�7)@8�@�'���������MM�D6�fB���%�uh��z�$�����c?yG��7nB��C/��/}����>z�8��vx:��j�
<���(��7kL(���⚀'7�p�����8�/]&X�v�|w�}l^7�$N���dD���Ko��Y}M�q���ѵf=����;���3"=���&�s�R�UCM��+NZ-;��`kTr�Y�Y�F���s�>��P���0��gy��Y5S�,�^�AY�� {Y.'6r^��RUc�t��W_�9�������z������;���߯y�W;��R�,��<���f����U���sJ���
���b��ǫ��8�����^B��RwdWc�
�1�x�R,T�V���t�>P�l`�|����1�:�I��i�ehO�^P
y��%�����j3צ&(hQrQn ��=~���3����8�=-���|Չ�˖��O9�"�M�dQ&�a62�j����}Le��l��h"�(?����l�������{�oݲ���[�.���l��Yط7�Ig3����0l�S䦣���i����2�6x�[�v9ŁO�H��Lg��M65�d�͜���,X��Κ���,�R��T�sr���ܺ�f�Θ��}�OgO��<�l�lHi�l�*y�Fpj
n�9����ޓh�Z�OG�p�
�yߝxm��q��wd��^ďVѱ|�-Z��~�*�GDު%�b�kjb�1tr���B�J �ׂ-��h/axr_��g1��c�3�)�L#BN�[�����+q��
2���f���.���j��<���æ�E����g��]����aD��yYE{D]A�%��Y��\*�&\�J��޻�! �=π����h2o��W��/WY`IK��7Z]Bo�b�V��G�Oo�Ş��槯��w=�E3�����Ȉ1�L�ӝ��U,ύ��Pt��S��2˒(1�x�_�荂 5�!�oR#"�\���G]29��ɁDY��'�.�Y����h�y�e�@�R��l�j��JÄnEA����X����k��Fje��VD�5'3L�dk{��U�V�0�>К���كK7n84t~dG&��(�XX�sČ|՜�Ss��B޴вohl��P3f�J�R,4c������c�,���֭[�9U�R���3�'����KJm�\�d&��i�B���>;u�g�S��%����su*�L�@Dd*8�12�%������r:Q�V����";U^��[f��%���g/^|���Z�)�|����O��O�=-�<SH�%��3DI����&�*�����E#x�� :�[����X�v#�����O=�C�G��݅[n���=b�|�э��>�L�����s���x���/���r��+�! �W�_��?�3�Z�O<�<6T^|c'�� �Y����n��ϡ�g1�����w��/��=����+��K�P�u�C���hj+��缯Q�U�dQt��.EF^�(UK"�ōe\�{��2��b�$,�I�5e1�`uz�nh��^�3(�*���c���>�jKk��{���t��A.+��>�Ng2K�Œ���J�&�\��H��^�O*p �.�0 `�@��2��^{����h���FѦ(��Ne3Y���}�k7����|��\N����9��ko��d�F����	�֩5i�=3`��{�{"h��@CC�o��胯9p�{\�ONVC˗/ߓJ�WǢa�Uz��$��Ü����>���h��fw��t�6;fȡgSF9��z��n~缓�)����#�E{�w&��an��zc^.R$)��/�[����A0���i#�a���M�#(���œ�19S������I���ϖDR�LIN���%۔Ͽ"8|�J�]��hMʟ~�ɿ{zkv 0���3_�q��tz�e54f#R�tU#���l��%�qx�=3���ڈ�v���S���܂�7��݄�~�C�d�[7c�Cw�ǟ�5�]�L܇��q��˰�.r�V,]��<�s�a�������_��8��d���pbhL�b�^<Z2�,�4z��{�O݃@$�]o����zqɒ^���q5jj�<m�Y�2�2�uY���B�V�.��"91���#S%�uZQ��^��$�y��D�������H_7�!Iryj�}����i��x������J��۱c�nrr�/������В�5UQr�)!>U�x�,@�9G�bz�X��g�7�fC��p!�P�Ff[��Qb����4*�qw�X�降5ڭ�2�tlx�����U
��|eV[�=Q�I�Y�%$l3Y�{��tϜ餿�L��]��˖�̩0~�5~ϫ���V<���v�UJŶBN�d*�͌��"���#�"�	IT��1�1�0�G�\Х��ǎ���vOnٲ�H�9q������ht�V�t�t!�u�2\U-�[d�f:�|�y�yr|B��02g�bM|/�hf2Ԣ
.+08�d}q�xE%�j�����}�z�E88����%�Jc�g�������3�O�6u��J���sUbAN�ڠ��1���=�p��x�����ILLN��=���N8,f|�S��@F�o��u��vXqh�;p���o|�1I��q��ص�m\{�8<x#�����0I C`���oA<����/�?���	���N�����ى��B	�O��ی����֛���.	�O&T�s�a>-D�8�̲�:5ϣ��gԋ�D���1��t�.UU���c��\ږ��F��<8��q�L� F�6t��z��7tvw?��͟���P���݉D��θ�M��=�k)�fyx���#��Y\c�3�C֨U����w�Ur���:�U3�4b�x�T�L;�����}��.�/��ݙ���l���-���lT:������V��`��;S�z*6��L��e`ٲes#�b́����kά~+0�_�t{�~�./�*"�Z���f���	T�%#�u��"'�J&f݅|�6p���-�'�-_3D�����$/^����^��f��ds9� $A�[.U.�3>���F�IЎ攂 �H�"�4c�0�����D(�UTr��\�(�$�����E���Q`�����l�����ޭ������s��1���D�(E�Z�h&����ю�SQ$�~T6��p��1FX��/���8��v��[�����8޿��]�d�&�6�P���x��K����x��ǰz�Ft�wa�����/a||���	��&t5,�e+aǋ�S�hD��Ũ�XM�f��"& �ƥ+!�|�V]EJ�@,�_���=GN� ���T���E3�D���P�p�!��˂�Jeޯh��	8\A���8Y�+�R�!��g6m��MgO�q�kpI�?��7�H�����v�q��\&�$��8�u��Q�G�� �������x�ω��h�\+-�sb@`�`t<vJ ���Ȏ$I5�mn9��o=�߲�ӿ�w����p���tB����.�\��E_���Ą�٢�N�hf�%1.I�G�2m2�u/똾عV>� �6mah(u���c{'''�S�b^��UYH��� ��~Qǳ����"���4 �r�VVr����7�vt����}�O��O�-[����7��9oc�A%�YBک�U�V2���P�W�Ղь�qّ8�~��"��X�W��T"&�4��T٨g�)1�\)�Ƃ$<G�B$�]����2_������]<�MF|8����@���S��M:�U���ŀ��ӸZ��^�CUD")<���б*!�m�?���!|�(�W��L����_�E���Bgo/��:о�tG���с��.��'��M��c�"0>!��>�8V-]���lD5���V�����2�F���a^W;�'G��)p7x�q�?ҴG
y��X���H����
���-;���Oo�#T"/��f`P��"V��,(�-������H4~.�+�����Y��5z��(�����}S��Bq�wFsGģqQ6`�z�G�b,�Z�ЌX�T�����g�I�C����#��̆Zo@*��/���l<��l�~g�����?x���*q0Saif�`A�"�;&�2YL�{Ed;r^R<��*Z�&��d�jh�`n}�5�@VO�9|ŕW>�m���6�ݞ�)�����z��	,�%$�$a�E7wsc�PS�l��L��+��<��jÚ�w�����O)o6oɮ\��W^~�*��n��Z59p�S�����xM=8��̩�5�"E�|ii�=-(�q�h��zcmT�5ԪMp�Y�"����xt��?�&��C�~1@�VG��^��ȞC�K�r�٠��޲|lZp	��� ��V�T�	<��;a�}rzdk�.���3�%E�,l'O���U+15t�xN����Dsg���J���[�_�*+h!<>���w7������y-�|��xu�Sh4�p��BU* d/�CN=s-�� �1�H�}{S���e�ș)5��)��E9e�IQ���c2�R��c 3�J(WJ��s����:��������q)�HJ���hr>ks������u9)���N�+mF�Q���<�"z@��FE!Įp� �/
�u��}<9U�5g]h&��~}j�j5���ΜEޒ�x��n�z�u:��N������-ש��2[��J�{c���aSuV�(�Cyզ��B��ht�����V���I�>� �>�x���g�;��`4�(ٴ,W%֚��W�F5	#�Z��Rhu�T���I��ɘ��i�Ǐ�_�q���-ݶe�_$�,�4���o&���jY�h5�T!�JΆz�X�M�3�Aq�� �I�h��tt}pVC����եX�Z=Jd��Y��̸߀1@�,q�&��vMO�-���,3=�=�+G~3�Td�,W��jIUL��F��wʆv�K#WTH%s�
E���B�ΡScݚ%��C��8}nS�b�o�ʕb����+hkkò��� �yw�� n�|���ٺf�	*2����cO"�I`eo7��6;��+6�[M���`( ��$w��,�S�h���`��n8�$;��DQ�$�F�JU���<^���0Yd)

�2��R^��2��oa a&``�: i�,�S��b��a�K�yϑ��q����¿|���x"��>u9��;�1�o���\�����3�Y�E~�������^$�8�2�Q�`�m��M�ߩ��7U+U�G�f�Ȗ-w���﵍��_J��A&D�eulTk���l���,�e=��U�l&�T���RGW/_�H>��@�i�_�yj �I�ߙͤ��\��y��.:g��75-�^*�hN�44
Ω�b6)��l;y����)�޴��F|>��,��}{v-��W늲Q��KLQ�5���0�%��r3E�QiF�d,�8�4>Vo4jL����<G��,c]�Bsݻ(-���Ο��d��9p�ֹ��gx·� �ZY�l�X��o4i��sٞ�I$��fɑ��$�W����/?�����ޝoC�*�c�_=��_~	�D��0�ۊ��;' �$�(k���g�w�^x�y|�ڤ�C/��݋��@Q��\��3)j㚵���R��2�a�6Y��#J^ZrJ"!Z�d�RK�<R�T�ALb�.��%GS����!Kjq�:��媷�c�F.cqO��j�F��JZ���F�O���s��߮m۶�F�G���\D���L����2�x��z
�}�F����3�u�Y�`��� /(���;r��I������h���d2:��dk�7�~�|��˞wv^N��g0��D6���P�#Z�а1P�q/�<��b�̑�lW׼�ޫV�M)�k���K�N�-]�R`z���r���z�T��1����FdK�G6�h�u�i�Aii"I�C)�,6�����3�Nݴf�z(�=�ic���΍45��_X��:�jU�/�`b��QH���Y�$ H>u<2�
�1�T��X��D�o���`d_��t.jөh�IE)��������L�K�����^�ժ��~���T6�ؤ3F�5�޺�c_k�U����&z0��Ƙ�'�V�X�l�դƑ�'q��Q<F�����S"b*�I��ΟE�%�W_}��t+*��O����聗"�y=}䜁뮿��}��w����uY��W]�R.+��fr��������I�F2�LMM�A��j�|�Z������TX�ZOѩ"�^��4��>`�QIP꬈��'2,v
�j�T�d���v������Cf��{.Cx&ܫ�XhI�e��BW���� �S.4"��r�����dSlg���uev����Jd
�se��F�Y�5�D�H�S�c%%��]΃�����	���x���١�tZs��ёY�BoЈ�&�lZYO ����6�1W΢%3�
��4��Ǘ/_~~�E,��é�?�ţ��]��t�̛��Z��������F��J.��ቱQ��2\.��}������w��QI��,�N^�3�����%�%I�Y:���7:O=S�B�ĽX��h� H#K @?�x���'s�BaA��d�0�l���ͰYPҙ��k�BF��7���U"��O)���#绮>~��ԹF��X�ь���3��lZ�Ӣ?tӦ�,�i�'㦜Ƽ3�ɮ���n��D�A�@:���MH�:1�a��д���w!09�}�p���X�~��(�y��~'� �Μ�'�r����%r�Z|�3��_� "�ͷ݌}ߡ���Kנ��"O��a0��5He�z��eVMlnpC+�n�$�'�/2�l����1�N:�~�y���H;�3R�}泂����*&-�i���ݍ�;=,,�REJ*��a���^o}��4�� �{��O��_��WOw�́���{2E*��B�G��C-�[��r�l@F�8%�\sF���:Kl˵��$p����ieF T���L0��R�*�jmh����^��~�����BeqSS����ɤ̇̚-T#	s@��r¤ӊ����o8���-Ij�xSKˉK.Y0���[�9p��fGC�W\��盾���EK�P��t�|Y����tX
�I4�6�����E��>E��4TQR�D:�t����:��5}2�f�h׼�ώ-�TJ=�j�f#�Uk/��N����B�Py��C$�N��F'��z��WE��Qa�R�ϲV%:�E�5!�����1́��Xg>g���jQ�5o����=��!�(!��l>�1e��gs�F�E���V� j�-���>�J�8pF�wݲ	����8;�b�����$fؽ�]��`�=��=�@XL�����(�]�{v��I��+/AU�3��;�M���&m���a�L ��x,,<���\�΀y58��h/���&7��*���,�T�Do�8���Z�D��m4Z�1�(`VG��P)GQ��5MOZ��]t?�9`�ދk�����r���T��V�H�gq�l�j,�����J:�,�l��Ch%��"�%TjY!�U.�8��̅��K�J�L6d�9�ں:���~y�g�Ξ_�Q�ڌ�̽:�v���@�\cC4��v:P*V��'�N5�(Y�����]��\�)0��k�.����}�P,u&���xDSb�zB�:�����N�t~�e�	VW<B�L��N"�W��V�c��'O}~~w���-2�]���}3���iЪv�yr:�n6e(��(^h2�
���0;�&�6X�fe�$2:1I-Dt
�6�ј�U&�x��K�|�z���A����7_���I�Rk�k��4$滤<}�x���OO�`E��TcA�T�24:2���QPcE���3� K����>��O����?�idb	$L�dlUF#^۹�s#��S���7w㡇 �^�):[�t9Lb�$����-*(�3����3g�x�FDr8w��TW�p�9�	�^=]�"�d���Zt���!�[g�+�j��*��f6O�v���JzMo0?jW��Hfi���֣�>o�f��&:�~���qI�ވ�ٝ: ���A�u�ӳfgϣ�\6Ш~�/��?��g�p?�M0��:q�H$Rù��;�5�3����~O�8e:v��eS>�:��a�~�:��esyd�<z��G<F��<Q��Xf�Jve�j��۷�wb�1��_s��tuu9�W^}ݎ)_`i2�l)�r��xR2he!K[(�!����ES"���W@Q��
�ˎtl"�j����ў<�g�9>�����ar����k�kW��j-�-hE�,�l0����I�d�}Η�cLf<O�/���q/�����&��$B���z߻����[w�s~U�/I#�{x�i�]]u����޳�oK�4����N̙ٹ�����JY]�̝ZY��(�1X�����J���r����a6��\�`�T/Sjt�^������t�cќ�Ba�D,6��� `�����x����ܲ�����ER�H:t�b�FZ=nJ�L^(r�wS�X)&_�,/��Rv�{o6�q/\�f-}w��@��λ������oC��6�s/�r%ضc'd
e����Ѓ�b�*D,&���B����=��j��"�{x��xX��qhm�1u��^ ~�|!�VʈĈz��0"	rjU�x0���p�^b��Z"t��/��\?�Ta��W}.��=�P/���NJ.�2�i(����G�Q�2{��ja�\�+[��Y���/���:%$��YmC��'5�#J蹵V�	�x���
9���~K���k_����c���k%p��[�O�>���t���Zb���*�� n�"�Ц��D B Bx=�ӧ��]k�,�
f����1�ˊ/9s��|���R*�J���J���'igѹ�N�&�����c�~�͘!si6F��/+b��`���}���.I<8kVG_"1rftbl�S�zi5���J�V���0�jt�%D�|���5���u���P<q�����Q�I
@�T*����f��w�s`�%���+���l��4dS���*���̠t��Qs��U4(㿹Wr������U7�tJ����?
U�/��6Z���;������]{@�x�b6?�ʫ����A?���A��A������Ͼ ��~x�>�&�I�>�f�$|d) 	8:x�8
����U���-֖�T�jx��ߺ$��!��GbBbD4j�5����p��^���3��g9��i���C�a`ۿk{��_y��.�]�,D.E�999^'5+�$�8�U̑ϓ��7~'�k��L��s�\6��'fJ���E�"L4hp�^,ƚ��ε��L�{����u�����Dre ��%�#�zL���4�L:��>�+1��&C�s�/_oW~%���G�:03��92<2�R�T�BT<����,G�b| ��$�f;�^4F�P��2�X,���`�'�Y�r���tC?9s欞T&���^"�����1~�jUfH�1�I�%*U�S&�� ܴg����LA�&k�������������������0
��G�1~��!���3�H͟H�[1��I(�YE��6�bA�9ك�g9�004�4M����d@�.���x\�	w�~�5~���;w.���a$�'����P['�5��;�σ���n��ӛ`���L9�(��x6����aU/BS$
�|ښ[`Ŋ��inne����b6i�v1�-�X�X�`�9:�ɆX	�����h�[|xL��U�{�-60���p�p ��-��D/L�,%LH�����F::�ozU�m�L�L=�l��@�5U�*
�$�y�;�PE�Z�M��^�9���֛��<y��:|����2��4z��a�q��1!�]��b��w��O����l��M�����#n���֯[�'�ͬӴjTS� 	$i�A���cU�)&��pM��~mlC��
��E*74<��ֺ�1�U��p8��>}F�|�Y�� �:#�ᢩ�bga����^fՃl&�l��9
�S������TUY�ț\�:_;f1n�"z���1��ؓ����ܬi�'��^;��\�޹�g��Y�:��q	�,Z��}�"�����UL��?~�#V���B-ˁ?f�T]*	���Y��{@BD�l�*�8< ��y+�hW����y���j��O��{����	h�!�Ia�Y�����N��t�~�F8{�,~���5�?��L�XjUc32�} &S�`�	/�Z�M�;�^p���6C8ڊ�[j�,X<�_���<j���9۲e�p���6Kx�Q5� ��=�
�~X��#�$�TRd��G<S��z�u�"���*Slhhh`�L�=�N'	��\.���Owv��<���_���ر���s���f�W���s��X�uҀd���}�ɏ�ǀ�jkP��Z
&X�@�`ٲŃ,��_�lp�7�{,k�����K&s�^߂��4,$�:����ʹ4�K��x�� :�!6D#J0`P���8�X���>_���Z���3���~�"��D`}j�"Pɑ��b� G%�fz/Rt,���PS!�"x�$�
�O�*u=�:Q�""�Q,����\�p�0���O�|��Ev�;�&[RV�;���.�K��ӎ���?'rE������2^�m'zB/�����Iٝ��)����င��K{��	�'���;Ol~�x@K!���/�d�sĂ���,���-/�W�h(f�M���J2��h���QNgg':ܷoI��~"*��&W�!� 8����ج�^g�{�2?�[v�Y���ˋY��i%�z�p?� 5��\	l�Ϛ+]L/�l�v�Jұ�"��E&h�6��߶C� "��:t��OU	8F�<ŊXKP�9�������%��RU�����'���7���r-�I��v��dFH�ժ�/��Lp�{Ȳ��8�ڲ�'>Gs8䡆��+W.�I�l�����q��c��gYᾞR�(;�fbYb�99.MN���R�0&���f���a�J��L<��3gN	+W������xX�x1�>}
ʥ���W:U�.tH<p�,�� ���Uё���"ԓt{jBĎV�C4�L�@Z��� Nӌ�������0<<bY�3���m~�OGs��������k�E��E��U�~3S3#��gpp�J�˜)�� �aV\ω�`q8����;o����'a��{h���`�2~VT�
p��0(�sC�.�gN����0|�s���7
�!X#��p��;*fx�x�MV��=�����c#�����	���T+&>��Qhn�&f�*�L:w$��B���2�/a���\&������6��)�*S-A�_�:\e�4<:ExD�kdTi����ź�� pu�$���ц
���?��d<a�&Y��8>m��ӏ=��/\)�޳���o~o}��\��y4�L�';D�j�%�#N ��a�`��g��Yھ)�-�{�B���ŋ�������cbK�Fbo���m/�G#w��g�4v *f�&Q����k6c��3v���$�\��Fc$S�>{��b�RPTvSûx!ɪ��N�K�*�����~M0W�u
�V���P�X;� [}��4Rr�C��X	�J߆Uu������i���+��W���_��o�x��b�܊b�{�Y�w���� ���Id��)s�3�S���D��\��&V���b�U���2�B��!�`������d� +������>0d��,�I��̚��pȜȪ?�D�Υ!�L@��L2�2E��9W���8�8q�Ɂ�v���႖��
�ө�x?(�=n�ё���*'X�\a�����x1{�~�2F%�C{��/��ٖBmYaC�$�Ĉ����
3�SbF�S%`��?U5��P���t.#Q6kD��n��{L�&�uL|��pS������/�VbC����W݅/��t�yں�;U�À!��#�3��"�B+���@���q��h������>&F텑�����K����4U�&/{D�p1�iOÉ�y�qpx���Y{���J�<�D��c�W�@O_?xhii#���ӹ,$?t�K��ќ4�����L�[*����E�T*4�.�l�L���Z��B�
-�=��O�>}9�}��76�X�wՑ;u�boO_���d�I�jN�׬H�W@Hyxk��������������l����S\��ik����x�|$�Y<ԝ.���_�v�y���<�(��Sd�6�` E�3<�_n|HPȕ ����u"U:�}�� hs�4�j3`���np�3On�r�R8��~��%(�=����I�醦�v�{A�J��.�~}�M����KZv$뛈�i��L��+R���Q�SU�0eé� qЁ��U��S!��!. r{�/�L?�g� ��Xb@��ā���#���x9�`ޕ'�PKe���C���uC<�X�py�DlD����:��G���e��~/�v��j��gj���x���e��׬Yc�}Hf������׮;�?8�fE�v`�>G-�EQ@tO�S�� �]*9��!h@.F#�Uj� ��V�?�;��4�TG�ws�́Ç��+�Ź�>;eĹO�����|����g ��B0 �����*L�DC�g���e��}��Df��ac�ز��緁~���2�c�,�j��H��X|�)]��9��|�J��HD=|��k�r��_�����M+����|��X���PK���@��wP����{��z2cÓp��+����&��H�4Q�` ��ðe�N��W�����a476A��\:.���c��tu͘ɪK�x���=G�8�f�e����`�bE�fs;��Q	.�Uϝ?}~xtrW���BvU�1Z_<���R>��6��6O����r?�}�&�J��V����:#~�>;�Ι�B}��U�DD�&���N��=Ϗ	�l����#Ŝ����l.��ؼw֬���/���Z�o��g�ŋֺ��f/�l��#U����J:蚦b��!����J���^�W|�[}�C4|��N�_7x��Tf6���5�11\�	�2�@��?�#�vcF'����(���U�2���3p��iX�x	s~b8���=A� N�'H��%ȗvՉ+��;�.j�*�J�t:X�A�B��V��Z`H�	�Z�Vue2�����y���7c����Q��P�4����[��.�:���@����QA��˵���߅'~Ѝ�9� S%���./@5��h?L��Ц�`x��(��L՟r�3e�0߱����,������t�D�C�E0f�������ZU�|��1��x�mj�
��Z;�I��?.z�X�Od��x�'���I�~Ys$Ro��<ES硟9���8�m���d��xUM
˪���B&h�Ǝ*����g	ގ>��Z�]���!���sL�>�t:�h�޻���G+���;DJ��O������*maKs�ˍ@�$�YA�Ș�Z���$���mN�C�<$�qĜf�!9�/Y���5s��j�����cfD:>n������B��,�969)sB�U�ڨ�F�u�?NDE^���s�
����f�����ܹW�ـ��vH�2��f��� A*m4�D����&��U�(*�y��b<Ԇ%)�2�1���@�9VݰL]�m�CC��Ǖ��f�����@��?c!HӲr[�<r��%&~���㱛
�������,���翃o��^y%�����7��n��Y���z�jC��C3�pc3SG<12��'a�.@l	z�ķ�l�*:�4��U����.%K���p��h>���B����$����R���d�C�N�~y�uk_�;w���Kۅԅ&̶�k����Hl �>K@����S�Df���O�K�0�K�*��5��8�V�k�lӬ�~<��ѓ�t"���
~�㿨jpj�N��]�]�_�p:�$�&`�]N��Qe�K�]�Ωag��bt�T)� z{��.X6V��>$�����Z[��c=����сڪ�>��Uy:쩴O�� � �#sY���0ȷ0k�6#8���^,�A���� �aaV��@^:K�
F�f��!rm8�K_�2��Cd������(:� Q� S�|M�������u7c�����X(T���nt��s�rz,{�%9��ep��n\n8u�<�&�`��O��U�  ���7����O_Kv�U���@�J޽p3?�A�<xo�aB�e:������9���OC&�b��i���.lܸx<���;��&��������s�6/]��y<TΓ���Kq;pj�e��Q 0���b0�o��c��P@Wu(�Xј
U�a��dk�|��O����E�dbGnFx�����*DzT(��������"0���H4�����������q\�w���(3�j2��J%�`��$3�E��}/�O雅�J���|��C�\3�^s���S[�lv⥗�=�����.<h#�P<i.�L9��}>$��Q{�࢕��B�2f(i2h�:cw�YX�p1�
�>�z�z�h���*U 08$�I���J��|��2x}8<nƝ�u;Y	�T.@٨����3/0�C6�TLg:��;>:�<y!9�Z�j��s��#G����}���'����}�v��R�m*�������[���k b�?w����:x�NXw�Z�<�~����@����	E�4_�{V���+���Hetft���D����߂뮻>��G�t|Ũ���%K����($�1V9 @��=JbJc�����g׬Y�y���$��,�bD�*_��l����$R1����R����#��|YU��,��@4�^���lmU��@6u�&����Y�A@��Z4ѿ��&(��Bi��mګ�f���E�IC�Om��-UúJ�>���9���2mP��{��f�=H̉��t1�xR�B5�\h�D�-^�6fo<}�f�����y�u��ɱ����?��/_]�OU'2��Y�~&;yP+E%Ȧ�P��w��[�\ɂ�)�1`��������=�	C�!�J3Bs����r�D�V��I���K�
bt�&��H�2�r Ql$�Î(�'
|�\n\0;����h}��bŊ�q�ė���-�w��N���֛�B�,q�}�/@ULx��Wছ׳� CL��3�u7��Y��7@�h8<�K1�/��/��sp��٘Q��38c�q�͂k6�	9��X-����� ?�H4��1Y�~�%f:�}a����#0����b���Ry&�A��+��4���M�����#)�(@�#�%�� ���v�h(Ѭ�LU��'�5�L2�'
�����>ƃB�`#cc�/�L�\0y�����N͘�����n<vpѹ�����h�~����ID��3k:	ĞI�� i�����d6���%:|	$��EsϭY�n�$/����clD%{��������ڨT�+2��l��i|@�́����%	$�fdh�C��������J
��ip������tBkk3�R�$��M�� JN�kbJiD�L���2%?Z7��L>�fj2�:���.�:TUU����d����g]���l��V�r��q�=ǭ7�B�und��^����+�?���da"������	�!7�	�|�a�ޏ����1��}�U��/d�o���,�~�28����_��?��j!-���<�8vOP����������ϟ9�M�Ŏ��[�̙A�l�/q�ضg����8�s���\2�$�cP�^=�z�D��P����t�)�պ��V �H��� @������L��\���39]U���3g�5�c^�}���sA�Q4Z�|c睆eu!q�x����V�k��ȚLtmqJӁ��@YQT_ p����^�vŤ�P\�������iI���O�����;��C�7mFU��<DB>�z'�>j�;�΂3���pKC������)0<1�B��il�Mì��/��ar�>GR���l�(K
nj�!~�kJΚ 	���L�\b���0�2
u��8S�ʓ��{��g'�\8
68�,Fs*=)�З���Ϳ��o�G��k_���*���%xy������m7o��o���8	?z�YXy�F��_�����'x���4�a�ϳ��l���*�:��FI���} �4�s  Plp� >T �G�Ӧ�*d��!"���wr|b�7nxb�¹ݶf¯f}�'���ZUU��pXhmme�A�⊦�FdG��TV��Psc����TĘ!��2��<�Y;s� ��6Q�nb��c�/�09��X�Jery^��^�b�Um�����۶���ԋ���6�C�F��'����s]�S�$�6�<Nk_Ѓ~N����	��v��^�5W��`�!^>���������׾����f��4�<88�$W�^1��_C�S���i2����c��h#�>(e�-I�>gd|�M/Ϝ="0������!���VF��`�K����Ě�B ;E��4�Hzj]k�MES&���*JI� �<1:6�/��Ē�?�<��B
���O����������ܱ�u'&���9�g�'V.��砫�������'�'���Cl����^��D(��FC3�� Q2*8��x�(&���;���?	C�(�L�ÇK)���F٦q��&�'^��S��kWW�~E������-04e� ������iH�2m�1(�+U6HL��"Ɔ��hkkʻ�����SʫtP3ĺ`�6S]Dߗ��%3���bI5T�^�t����Ρ����
,Q;�w����C��}���-�	mQ�Mi;�Wz?�d���uA(�[0~����ֶ�w?�ٻ�?�]&���o�Q96����ǟ���[�htm!�sQ)��CZ�u$��S�i�$�j��Ⴆ��NC2��`)
��P��H�(!�DjM�z��Șq�j#�!566�ﹽ�n���UtB�T�F�&���c�J��R)y�����V]w��Ճ�b��k�x�:�������_�pq嫻v��i�{7�+��A�����{�Uˮ�e��7��]س}3���w����7!�Y��rܽ�> ���AQW =���'��ff��:�Ag:�-Њ��çN���=w���k�E{+�W���T8>_�(�t��'��Ȕ�:S`,��*f?'�sҴ������T<���h��M��,�i�0�O���H���"�K���i��T'���UˮޫL���U%�L��曟.U*+�a7�:[\�gU|S����h�"n�@(��A��A��������/�Z�條D\^���o�56rŁ��ޡ��Ȁ �С���i{��(cp�y��'�B6�����G��c���D��/���9s.\�h���bA�(R� l$�c�U5��R���8���[�d;���i
��["@IF0��7�7g��q����fKC\�B�:����Fe�S��7�f�����o���F��G��N�]��?�C��?.9 �]o;�	:�u�(D��A�Hl,K�FܨB
�!��?��Am��ç����Ͽ��K�g�����W�-[��3G��_��W���g5sS+DxF��)�u�2�?u(�v�����G��*c7���5DR>��)N�t�0I 7��B��ܙe����.N<��c?s`��������h����`���vq��B�Ez/��P��r9����Ḥ9::��cf]N׻]s����l���l68�-��Ӄ�O�y��������<1��rAC$�#��~B�=69f�!��I��H��4LE�x:���0��`$���Y��<xDа!��#��CA@D��l:�M=S��鼫�J���dj�$C�y��YO�����s��\v�ヴ>�c�}�a�����Ǐ�Z�7�M�׾�U�0-x����}�{���L������m���o�� ��7�y�L���6 
��E��<������DK?��b&��r��~��~��+&���h061�Fմ.�Rks[5fe�& ��\���"��N𠿓�ފH��"��@UE����!( �E�`&˦3���T
_R��5��5K��x䑟U^����{޾���6���F���:�0��}	0��E����J��b>�677�kooݽv�u����7�������E�WQ�[K�B�n�\�PX��%�9=����"�xp{�Ah�6�Û�Ĵ�N"9f�<8J B�¹��i�,#!+�
D�T*�j�-���q�{�����;e-D�B�֢��LǝL$�9}f�����6��e5*����z���o���������?~����(X�	[��W�d�+�̂J�kV^Oo�3V\�X�O���a�8��o��ъ+�Y���j.1ڷtF�3_���O�i����9rDzk�;����2Mբ-�-���l�A"����܊�>3-��@>�V�3#��Z��T����	.7kQ=2Ur��������}�V�z=���������S��ڵ�^��_ij�y�~&%.¥DaJ���	Sj��Πd� N,30L"��{�UK�ڄG����o��r�e��O&�*��!M��K&�~���Ke�| �(��5)�
c��R���&j���I�Ɂ�x�tpxZ�ή��l`����\'N�|�%�D��q91��L�����,����k�^7S	e��XR��ѱ������iC`�e�:@�h3Z�y�ᇕ����]��y����}�)u����WRU�ɉt̘�Y����`�2tp�C�d����A�,�"��t]-���G6���<yO[����q���������x�����9$��8[?&�� ��0"�7���8/�gjS"g��k��[u!
��FLx�&�F`��A�U$����}��t�6��<��c_��v����5��w6oH%�O#���D�D��T5 ���8Y;������.���FS%rt|ܒ�β K':fL߷q��I{���c68�-���v���l�0�&�G�O��C�L�Þ[��$"H�HZ�Rۣ��b�F��������ys�����-���i�=~(��ð8V)��.�Zp�W�X��(S����s��@�M��(��ѱkN�=����v�ƫ�`�e5*��瑰ϻ�_���{?����X�٤��) y����(�-���7o�S#��n���(��py��|e<XL�bY�X�����<��{6�p����?<�����;��^ZՌ�p8$D�5N ᵖB�U�nln��i��h��|�tX8���?���~W$VI�y\	�6��s�,;�c�$��j:[]�d�s]]��~���i?����ض�����eM�l�E��"&���8���U'h�ޛ��|ll�@����p{k���n��t{�Mx��2��ڂ���;�N�*�S'�J���T2�Ъ*G��^ '5�������"W�ܲ��)Ï+1�������U`td�͝0}�t�xTF:#C*��#�����Ä�8vhP/���֖�ߝv��^d�����Jf:��_Q4��]ｲjê��m^^�ڙ������g���֭r����y��}����pC ����޳z��������$8|aPKxa��W�4�3�8�02x�f?����¦fo��?\���x{ཥ�bi� �R_����Hi5�M1�*U �[���y�~���H"hP+�UF�g"la~������wF�'�����d*mj{c�ޘ>ݓ��k#�����v��g�%EY�t��n��%���b�Z��66�L*���I�
T�g�~���e��kٲ�o��ڔ}����ŶvѢ\yBٝN�У���t�i	��Uxf,���07��;1(@��@+��M� xRG�B�R���^P0�L���*��INb�J�t�I>S ���,�r��P�5N=���ZN7���T�8
�g��;��!���W����:/�-����}���V��=s���ǃ����՛Gᝃ�����$���xPJ
F"���hz1;՜i�?���m`p������rMYQ�54��hS#�<9i��X�����zK{������V ��TAMi�`�ʔ����-͍�ߣ���'ѿ)�/�*V&W(r��5k^�7��慄�ڶ>�D�۶�X)_��.���d�@�a2ߧX���m7�<�*J0FGG�����?g��;�X7fǀ_������=��T��ʶ�ۢ��{�{�x��[��@�U�j �+4�(;����@��%@7t���'*���8p��3�f��$�Lc ���D�Ě�1��Zd��z������)8��Q���AJ�Ԗд��	w$Y���}f�֧�t&��}Ğp���d:�Z������i�O;�~$��~?wnh�:�j�����&8A��p��@�{�-ZZ:52�|Vۏ��{6��d��a���+�;n��*+���D�� ��"ʥIΘU�M�ZgN"����p����W+D����S��IAsS}��u��gF���#pW�RY={��׼0{ƕG>����Gy��u0x饗[�yi����.�+*H�*ę@3N�~H�O�E"��Q$7
X<c]��4��|��`(�ʺu�OaR�~�f���r�]��n��R�<��s/������9C�BxEcÂS<�$�J?ڌ�4`jm����"
�(�*��V 6:��H�i��.a�N�P���ࠡF�Ϥߣ�emk��=(Z-H`��dc]N�2i�����K�?��gS6���3h��ku@�s%[~��;L�����F�w}�� �	�m�Ұ
���e�}dr���X��i�����ŧn�qq��Xb�@$On(�J�=>�LU��e,�NfҬJ������� _,�����B�>O[�L�"&�c��C4m3)(#���O@:�#?6��llV���k��歮W����ޭ{={�ܵ�����1��v�"�[k�-|K�ZՀ��>�/t]�P��Zn��8�Y�|��M���g�~f���[��� �}�̩�F�㯛����@TT����C�z�J�J�
�.���:�!&ρ�?�Tox݄��v�75F@A @�iԛ$ ��yYi��9?�3���^���&����s�[[[}����ݧeU)y�R�����1�O��Z}%��3~������ҰZ]_���Y����> �)��!��Kjyt�o��9O�كl��I���/>��K�*Jq%��?�pS�A��/������;tٖ >L|��[��|�1@Ў��>��^�� ��D?��l�h
�|4����k�n����t;a˖-����޵�~|�U��>���8h��K��NY�����Sr�8P(f`b@q�
OΜ9��믿����f��#V�'&��#��y+��U����+E�j`���  �mA�Fj�C�����A�����(�H��Ʀ����6�\C[�@аd�2�	A ���P&As�=�wN�)�0/�y�j�Jh�,���x�&b�dy����;�U�W>5>>ޏ���]6�g���z�������3�|�x��+52qɅ��hr �rU�TY=g��_��֭7�����v���P,��P��>�O�C��!���v�4F��o�;��&���)"( �NU?�Rr��k�CT5�a&V��'Ґ����bQ��^��ߝ?ca�}���p��c���Ĵ��_��ɵ�P0h���(���uB��.��w=Qp���4&I�~�t����6�|���^ye���!����@8r���?�EЪ���*K1�+%���. �@�βKb�@%�|��[gy`V�P4򠐂�a1Zf�jBυ^���BGkU�2�R��$�B�J�"7N���7:t�)F���/�*F=�0f��rEF9o"�'3]��<�+ՎT,���s���K�=��k38N����������:y������7߂���J���[���<r�om�Y��3�ly��E���qs���sM�y�a�2nk��YN�*���(7�3*b��3'���������9�D���eV�������!�b��ɛo��]��ڃ�>z��֋f�j����-��6;�~A5L@� ^m%�3%.�'&�p��9��JY�T*mz|�ɆhӫKV,z��[�%l��͙~�l���\n���I�tW��ͯHEg6��HV��w���A�%(�x�;���c�<�|�Z&��!���L�b:��ln�V�B� b����;u6�H��S�Ū��@�~�"���K������T� �����(�Q4�u`���J���w:#�W*o�����Z}�?�۟l޽o���7�2�9V�h�u�m��4�����ڹ��"�Lz���E�4�E��'���(�k?�(�aCb%ų�U8��c��B�B���ύ _C��B9��f
��T�d�зhѲ��f��4��w�V�w�z����=��z;N�L\���AR�¨*P�M6 I	ĝ@��ĐJ3u�E��p�{ﶷ��z�����o�lp�;f�~�d��ّ�d=�R"Q��$�\� A��e~�Z��h���>,�Y�T�*�+	X� �	���Q�t�Iё�;��J��j�m�*e4���͂�xƌ����6)]d�dl�����v����X,x֩�+�c����z� ~��^���G=:�4U��UW]�tWqQ�`�e��=��w���B)�JQ���jL�U(�j�G��U�L>ǸdAB� ���l�@ ZkQ /�q�녆�x>�&`���\�\M�c���_�q���K����#y��w�Ͻ���<�{�,��3�V	�j�[��@sE���v�x��<$)�=����s��77�s�M��0�Z�o����>/59�?S��f�jEr�N�g� !���P6ʠY:�4�'B#��/:'�68�m !�
�8& @LG�|�X#X���)����%{ͨ�6���%�R(~�^k���I��>��תj`b2�l�;�=�\!tm&��50������G+e��0�z{�M]]U{���e�O�����d�z]7f#(��������&&&0�>$����@�<�,Jl�����
x�)��x8Wal"�l�e���x��m�ƍ�m����c���>��۷�w����7�x�U7G�Q��v�˪��� "% ��$����$`���ѿ�T�0��x0|e�uW��a��,��7��ez��R�]o�.�������h+W5Ī���v�5�X u=T�Ztdxf�n#F����A�G�	'@Q-���(Hxh
� V��E@���0�Xղr�z@�h`��4�)� 
X�ݦ�f��g��9Pt������'O���I_�ƍ[����ڃ��[�q��ȯ�����8�}vI&�^�~A`�y�nV1dպX"���Ln��i�Z]e�g�|���<
@���Bp_5�R.���t*U&Ӆ�?}w�M�l������ =r��-�+�7��W������%��$'����fd��|����Lm�#(a��HġPf+��Ϟ5��/>t����1�[ ��+����5}rrp�I���A6f$�D�F$�=��i�@�)�Ap�|&�d35��NX��ܹs�����@��|�*�L-\�k ����HTd��+_`k�4m=�Ag�4�Q(U��v�"O�c|b|� r����ͱ��-��wfΜ���l�m0�O��o?ޚN�ע/�C��h�h�ȿb�	e��B�c��m*�68��c"1`�CP�鑪��\Q:�Gp�M`"�+�����^����8��/���!���������m�]劲��6�./OUC�?���Z*�H��cm$�9$��ڲ��C*�`|�!���"����_��S����Շ�z����?K�D�7�����Mp���� ��S@:4�@ˏ/��E$"N���������S3�ho�Vcp�C�����Zą@}J�}����_fDJ������v��� ��(�F7�8:2�Y�悅|�3�Lw�z��;��4l�!��q���u^�xqU�\X��B^������� ����j�� �k�ff��$���,���u΁�d��,T4�*�F���^�ꚿY�����?y-~�tl}��������V���~?k/�+*�+ڊ�D �!��@���f����'5
v���>��z�lN�>2f�ۦ�{�����c��O��nת�D5B�\�����<��%�b�9F����1XQ�@��d|~.�c=љ3��{Q0���j#)
Z�Jx��jE4�P�V�@�L��e�m�`xt�4�<~p�e0�"8D��`[�kz�Xȷ��j�����vŮ"��q��'f���T*�f477�n��''`bb�U�h(��$�I@���aƎ`���KL��+ҒXc;-c�O��b	2E��u��-*'V����7�q��?z�����wZ�����g/\����nE��͈��Ir�O��鶰�G$$�D���`T�i�q�t�/�
��[u��o�[�<�}���1�>_w�u�y��O?rZh�����i�JN�d�϶$���i
ـ*:���T4�Ob���v�+i������+���q�gs����Q�L��`A�2�J�i<�r165M�@:���N�����L`f"��k)W��D�4-w"��[QU!_���|f���1�%�r�m7۳g�w˓ϭ�l|Y��9�N.����k��7T�B�~G�7�.@�c�91 �v����/ɿ�'s���4�\$�j��\�rf٪՛7���ݯ<tK�����o;����>q����aI��"�|O�w���B�/�+$�	���	�ؗJ�X ڹr͊����8f�������KF$Iݪ�?=�?,��uWlr�Y�*)��;-J߁�
pU&�d�x�^�!�ʚzM��q����+�RV��U<>/x��s����T[y�~%��5(S
��09c:���Y�(<)MR����ric�Rj�羲.}��{���Q�}�����s�м)�L�4U"b#�-)"�uD:��:�(��Z��g�^?���M ۋ��2��d
ʥ�Je�!�J�l���U���u�ݯe'��~���p~{{���[n?�s�a��cp�+m��ŁC��J"�2��|�(���NgmΠ�B"�d�	�ae��M�v��x�֛��g��>�f��>`t���X'��o<QԊ��o�,�arlD,�!�\jIe��Z�V�8�qh�e6I`E4�rè��P �e˖��A�S��lu�� ��K�*l`�T�,Y�{1��>4e;���Cat|�8��q���\ID�r9�]��dS��̥K�l;��hѢ�����Q�;v�wn߹�řl�761��v��$;j�$$u.�uzr�H�j���a�����l�*��H%�hW�\���,_�̦������?{��K+��Jx�'BOo~�SǏ�x���������1P�&SY%1%2��f:�.v=�L�U���Kb%m<mj|�3��t��Hl�H�l����=='�ͯ~��bUJ��7;dw��B*S �$���d�9���\m�yJC����K�
>���)ŵh��e��l���i@ ����@ߧ�: xj�He�MB�ϩLJ}Wzm0T�,�bׂ'/q�aZ��7������&���c�/�]x�c`�mQC`�x��\��}���pG"�@�˰�੊��4Ee��������o� 	5�UjC  pP��Z5,L�����]�ܵmF�1��bJ/���+;޸���{�BK���@�=��U#ǰ434EbFk�le��e�롡!py=�$9z#��'n��η�/�����G�lp`�ϵ[f�V�9r�I���YU����E�ڂɀP��h�3x/���ٺU;�1��P`��(��ѡ_���F�DU�t*N��>
5A&F��ϫ����߳>p{���LD��*�d�m-P�!�H �� ����D�W-�VE����*�6���
�bW*�Y���?ڼtު޹��-��ɶ���<y�s���}}��Ig�.�!`k��c�UopP��yj]����N���C�g.�UP�?H�����aqV"�-�ta�ʕ߾��۷��W>�������-��>sۛo�~��.uy}�8�u����N��T����I�ɞ�w�k2�T$�O� ��J��w��]��=�\� �>�f��~��X�����}���z�P5���ܚ�O���.
N��WjbILͱ��h5�V�$h^��	i�����2���S��Bh�ZQ��]���Â��T���0�"��Pⓓ`Z��60�
Xx���E��z!�9I�=Z�\8>41>�<�7�����G���	��f�oШ�`��kϿ���B�'�����$Z��!��&��EI�T=�j�@�u��2y�f ?$#��B�Ęs$Ů��V���8~Ţ��zǭ/��ܛ�߿��ky��ǃ۷?s�[��}O�+������)��O:��t,�B���)U-���Z@`�����:��pkG�����+_�����m��-X�@���9�������Ǫ��ܙNŦ�i���`Ǵ����M�Qd��頧��n��@o,]���8�q�y�P�� �R.1&�J�ɞO��*$�7v4��Dd!�N]ڟ�*�f j}Y*�蠎l�T����b�ڦÇޛ9���V�իw:t�{�ʕ�ض߄! ��~��m�O�����R�pe�T	�x6�C�Ԫ�D��@*���.w�/�:GBJD�L��e�l{���lV'�΂��5EI�����7����Oܴ�/~)�o��|�n�~�;{�~Av:�^������d3�1Q������)����2�%��Ɇ�ש�AIA��74L6D��/Xx������`�_}l��l�m6f��Ns��G�蚮ݧsF��)br�����H|m8qj��HZ(�!�E����NEU�@"���Z)�ߡ̃�z\n(;+����]:���9s@Ȥ�����hU�Q6����k ��d�k���/�*�������������:}񭁁�Q{���_��߶����ۖ\��s�D,v�]����/xb!%�RV�Û���ZS3=��CY;�k%߁	�}�G`M�S*+ �N3�L%M���p�M���z塿��;> wN��1xi��7����/:��E�(�U|����G͗�kc��I��>��5�`!?-����\>��^�}���⏏������Qa�eu��:�,Y0�?�s�D̈Z��5�4|��I�,�ěh��
�Pe ���X,��b��l-хA�Q,���WI �\,�� �}�/�R���t-��� +�Z�΂����2fVN&S+P�e�~nq��DX�s%s�i�b!�Ng�$'SW��n��®�Br�z;��v��ȑ#RϡS͛_z��T��d2��X)G˔"+@@���-`��׬?�A���BL�&eE�L6*�c��"���T*���u�'o��uK��Ƀ~�����'�<}�޽o?���{���y}`4�`0����{/k'�^p��
��
UJ*�f��#7������=w<pt������1�����5-��_�~�}��i��}�oK��r3|�WP*��� �,���k�n������L��	���N��C�eQ6�`�*�5bD�4u�pyX��2!�x% A�M ������D�J�4�X����XU�dd9��s���'V-�J����JS"��?�۳����޳�w��u%{`Ѷ۶m��۵�����#w�O�?Q�(sKJŭ�)l�3s���Hw5������&s��3w�F�kbF��*��9H���k%�O�⑦�W6m����f�<���nQ���C��������g�wϩ��/E�^���I�y�F�dUu��$�. �w��#=#�-��P�Ԓ�b�X�1c�ᖦ��z�W�΃m+���m��Mi1|���lT��[��Ei��Ȩ��ts�^U��`�<`��ZmG[`bb��	�F���E@�,����J�f4�d���;J������U�e��}����R������	7�㍘���Ǟ����ǜ���=�����,�,,�@� /�@B�eZ�m�)_�>3����j`�b�V\)�LfFDFD}�w����m"�J��Bm� �� �Y��p���:r �	֯�J�U-�2�"���K�bԞ� �6�"��e�8sv��Bm��3�~��?=���W���n�GH�c���a�'g���=�87=}[�Ӿ��%6��က��l�q�mq��L@�ԥW��a9Y�/ҟ��V���깭v������n��G�����s��������7���m^?��$^J�g
E!W(b��	G��d�a�����)��d
�)h ^�~�FDQw|b�˃C����}
v��7��� ���YS������'m�"�/w];�h5��;]�u P���,�C�SV)X8|�ur�n!�|���y�1�`1EFj�� d�l��:d�.Fн066�كǎ�"�S@�0��H�%K�,,���D?��FB�
�,���Ut={������O=��ȩ}3���ٵ�IABj�CPp���տ��ȡ��_1�������U�vg��*&$���BfH���8���^^�ǌuȬ!&!}��$� ȿ՗�=z;ٲ�����[������q�ſ��ѻ���<��|>�Q�CV5�K�P��y�y�{13����,�5���N�i��+�+�b�����[����Y-����g�r���G�>�X0�~knf����EҠ��
H���_5<"z�>.�M�E�"�Z��6��Da�����'=
pS6ן���ck��n���O�٩�{U�كI���Z��E�Z�>vR@$,v��� ��t
\$V�f�����T�gg/93y�G�}�C'����?]ݾ�J���}�w�^��o�Wy���/;}�������jo�OeUÐ�C#_ �����P��j� �]
I7�-��F(�Ad�7����ul7vܰ#��+�m�����G׍���[ ������~�k������O���M���5���p  �%�ÿ���ry<�a�� Z-˦h[�er��֭_��k�|���č����Rp��?�8@XY��W����,K����{��R\X��4�p`�,u䦡`����m�5�:t���]���a��A�A,L�%�&�	@�(C%�Xd�u5h�B@>J���ddd<)�J���)H����@�b���S��RP Нz�Ob��$d`˾�uU��������®'N�;|��s۶�L�����I-�_`?����<��Ƴg����=V��#�JD:K�h$�b�|�~��88 �{�M0�q2��#�ޫn�
�=���ն��a>��o��ꫮyr�.���!�/>���k��[��������P�tP*-KL}��.OA8�9gZ%�n`�.�kF^�'� �w� bK�׫C�o���w<r�'o]���IjobK�Aj�,�i����ɧ��/c��Ʃ�j7�{ȶ{�HX`d�@�D�s(8����"�-Γ��
iԗp1�鎰�$���@�$'�)�����ڭj�����pc��v��ȱ����m�����`y%��`�d8���vh��x�_����Ь/]u���WN��������Z���Zb��~��U��޻0��N��.w{Dd�l]�P�P�ߥ�V� W���	�ޔ#B��ʟ� o�ؐ#���&���G������������޴m�O����Պ9	`_�����o�c?z�j�������I�̄af��7��,,,�Vž$r�e��T���Y.kY����2Ʒ���=H��\�Y{�[
R��؍�A�����{�]7"a�."���M���=�� �S�d�k�h�t��y�s�n�
����!� �
K�+��P��L��8f�ġ��U>�T�FH�ԬG�#�.�"�H}���V�A�8�%����,�D_iUđǑ&D�`�	ʎm�ﴛ��?�ܫ/���ͯ|s�5믙_{c
ުv��w�����\977��v׺���Ua�A�A���3|�(prT]�.� 
�� �q�;�~��r�1��J�R��oJn@>C9��o,mۼ��}���>T9�����.v�wf����~��S�����|y`$�A6��#����ǉ�хs�8�F�A@`��X�}
t���o]{ݕ|h:��\����~i�{������_�_�я�����Um����'�+a�.�*	��aL�F%�qa�hx
��1��g����"!Ձ
�apн h'�Mϐ��ŅH�8��	P$	Jt�cb1�4)!A1�pN��1݁ 4�.	�����B�UYj�7�:�wOO�;��ȋ?���ҫ;/�|zמ=M��0��.^B�SO=%�ffr�NLn|�{w/��������T]?4)@F/	���'�}�ez_R� �q���
��;��AA���	Y�҈�}4b��ޜ�׵�S���|�����F�������g?{�q~��_/|�K_}�+���G�lq�/
%�0e��g���t '�@��!C�"<��Y��h�vL��[(珔���sã���?9������ �_��ŁK�ْ��ֽݻ���>�J���v#z��c�\�c7DF0sa�e����	�ꫯ���$9�`YF.��&aP��2,\�V��e �����B0�"�X�!s�a��jo}��_��0 tT��"��c6�R�ࡼ�P˷��U�zc��3g����kO���+��t��}3�#�F�2$�]����Ӿ���T�=���̹+��nh4���0��ڄL
r��q�� dr�c�ĸ޶+�K\��!>O�*��	�����H��ݘn�͚�#���ڲe�3����|f���X��n�?��~�޻�;3��J��ݏI^�r���4��������/%$e8N
F�x`�	 � �L��b�on�����'oM��Ef)8H�nK������K���E���N���>T&='d�Ht����Ap ��Ry �ݮ�Q�"��K��aX��R�(&�
Eb긠��Xi�B��y$7*�~���q�.ơ��c=E��D�r�� t�R�1v^�����%��"�F){~X#'׳��z�ҩ��ǎeh�����_���\��$I�Mi�}�k�N�����GO��v�����z}w�q�z�_���8��@"xIe,)��s�!�{I�X�*�|"+	( ʈ���ri4�i��dÖ�����L.\�a��K.�z����{3��Y`�~�>��-�N���\��΋��� ŁA�Eqa���&�bW �}}��2�д��إ�`b|��j߾����w{
.JK�Aj��u���Ϟ�ǿ�=t�@��h�kq~iU��Ӏdm�Vhc��ԩS�Ci`zz��!smy�"��5vZMTa��T���^ZZ�Z(�I�����G�b�@�%>� ������Y��,.�k��� �H�(��U�m��>$`%�AS�~a+�q�c�Y\��ڝ��3�;|���U�F�lܸ�'����u��[�Zi]��a'|P;�����Ï_2y�������f�2��׸���%A�UBW�$�؁ 7�E��� �;g�Q#���Z~�+��H掀�8�&�΄��(ٰaS���G�ձ�
z��g>�?~�������~���˕�����j��M� :&�H>}3b��tT~<��d, c�S Q�7b�0�r���a�߾�|���?r6��� �_�]s͸=�/������g����Gfg.���@��	�6 +"%ҁ��Xu��,�n�ԗj$kf0��r!O��"xd�e�<K:�G�^Y Z,9��49��B.����	#�[��&8`d-X���>T�x)�B3�=�:�J�yn���L�ر���������v`����?��Ys�Pkc:.�g��wKO)������7߻uzz�ʹ��ݶe��L�&���F���$^w��c���?�/a_����}p�2Q1}�G�C PFP�r`Ji�ץ�t�\�m3)�]��Ӛbܷn�v�3��������pg���寮ط���e27�iT1�*4(�
z�2�z6�3:f�B�� Uem�2/k@)D�����6�M�-^�ƍ�~�����dv�Z
R���ZAp�s`b�\��O΋���S�3��"[p|}j�^''(@ز�RRo6H��Bg��4����>�rx>r��&
"A43Z��X����t7�t�T� �	���ɀ�1�>��B���O�& [�Ǡ��N�S���LFI0� F�A/�lO�4U� �T���Z�gN�����3��X52���������e�]�N�߬��������h���ܮ���+�jK�)�Dy؃ԉ�a	u+��� ��"�0f:�Wp����W'�@���A�H��-c��pu��\�}�4#�i5;�GGG�߼��W>�]��q����������<��bqwǃ��M��F�3��ND��)(�q�H���d�d�"�A���o]ˊ)`�������/ݴ罏���n�O3��� �_�хR�gyd�7�{�=��������K�5���k��F6mނ�V���^�	��ei���,Ҭ7H&W �A�d�&�7�,��L����"SS�c���8���a;DsR$�k0ڣ�(	y"��������f�(b�(�������n�k�|y9�D7�J�Jc��t�����o?�9���+//��y�W��s6l��U��U�V��J;~E�B����3��]����<5��{~�ma�~u���b;��=k>�%Y���|&GY-y)PF >
��6%�L9�M��M�ǐM��v�%Y7�N m�>/"�q��z,�bmɫ��O���g�������!��?�g�����ο���;��n�4���*�D�Cث��z\�C��u��jȎA��I23�DR�pl
zwGQw�ڵ�KŁ���={����4o���v�[
R��h�?{��3��y�④�l^�o^��]�����u��^�G������H��v��0$	��A� �24*"}H3WJEҩVQRd�c.U��uK<
r��[��B�0xD�k~,D�k03
.���Đe�GU��ѡ��W�R�b���z`w�h��F�
k�cQq���:�N�;����{ff~���&�������#�6l�_�nj���Z��4�)O�n�D��D�����C�����cS3g�k���/o�Z��cq��x���SzM�`Ab�%�� "��qZ#��ZB�/#����g�`��q
)�!t��0�A�S���Y'��0��#G�����kן)d����MR��m}��_V��O�l����y���_������4�Ē�/M7�t8/�@�N�}�j�ޯ�j�(��>�:@[��s Df6�za�Z��M��'����oK�Aj�v�f|�>t(>��k?�o�<��(��z��xi)w��q󥗓u�/!펍R�(�Q��<�E�i�нPo,��z�A�}�R��
�ϟ'��t�`"������lp��b�������ś:�B�}�}(�[���c�5Q�l�A�B�` FS�K��pn��X��_��6�v=�7�ѵ��u�"]}��L��'�9�Hux������'�M�~��V�S��{�n�'���ف3gΨ����cwݗ=�8�j��������Z�~i����E�X�E
��0�e�f  ���grjoiEQ���� �)�sbN6d@ �$@�!d��d��?\�pފ�{�[`��z�����}��#�L6�M���G׎��h���������uw��W�����?��e[��2�����T�%��Z�E��~ATT:T�7�K���g8���m�'��Mlz<0�<7P��
��l�d˝�|�?��;R`�V����m��.�g*��o?�Ѓ����1�U�ѭ�:yZڶm*v�-�9άDPXp��b��f6O����F��,i�sH2�(-C��HH�0>��Œ�-ig,`�'b{"j+��+��Qeee�����X;�c��LuL.�'@v��2+a�n��De^� "cdzNhڶ[�5Z�,^}��T��}�T,�8328x�4���'��|���714�n�S��C���NGo����TΝ9���l�m.5V5[�ݎ��F������C1R�(��9p���9� ���V��^{��b}� �� �L �Xd�0x�OI&��`p��C`Q����Q��K<�j��J%�e2�cC�'G��&֗��7z��^��7��=�'ϼ���IY�U
UU3��I?�� �
J���e�/�� ��hbI�����\a)_(�xǥ�������=��l���R����~c�7�U��{�ɗ_}�c�f�3�ӫ׮[� ����%�	<�����Lc�Z���Y[�K�c�iu��ET
$2f��Q�G�q	�Y{d�Y��X�5�C����U��BqE�~��.��pbY̝CRr�0��<QG��&0��<�ˣRQJ���B2�O���.5Z�5�ӳ����ƒn���ba�R��V��J�c���ݳ��`7W��t��ݻ/��B"HD���xfQot�|�{�sK�۵��F�5�:����Á��7� R��iA�y.+1� ^.Ba%F�XF����.�
��ܙ@�
b!�<0 �KN!a�"�#~?�}�ܛ�D��@�Tʃ���Β���Jb�"Z�Ã��s���ǆ��˗�G�~o��������ݬc��12�aj%Ȍ��@Aq�R�*�L���� ������ �(��4zK�������Û�m��o��K{v�i�ܗ���� �ߨ�E�I������Gy��(J0==�n�Ν���!���
�ı%QQ��p�~,�K�C��� 9� ڰ r66�E�:x?}8�L�����"�>[�è�!��)`�U� %,�|2$��w.$�v"O9\'q*��*"�Sp��|	�0@�����>��vMWuE�!��ڮ��|kT���b��ɞ��mC�k�|n���Δ+'���|�|�`tF������Z�l�ڵ+x3.�T��X���ڔ��͟����VmC��Zӱ{c��9�S�����A��OA �����A�
����],��M �'p�LE��{�#^ъ��!�� �,�Τ� ����}�vll�`Е���
\ʊ���|��K^�f��=����/>��m�"�O��	QQuM6D#�GEC�$b! j X�e؏�������cE��b�8W��ʷ��ۛ��Gv����Gߢ��������g�y���|�G�<��s��\7<:2��t�V�!�VO�&��kF,���ת�F�D�Be��+8�t�A@t�W�)T�0�d�,J4b��mX�čx9@d�Qد%G2�:�*�16U�;wQq�^Ҧ�D.���.a�u�;��B[��ۆ�K�h���t�0��T��s�� j���4!�$��4]�躶���b&���e��*�g{�������@.gg��r>�V����i�eY�V8p{kLv����A���	��R/?^� 9L�^
��ǒ�`~^my^�����^Ǩ/4������m���v�[�u����[eu����~P�]'KO�!ʂNO�R 'd-/��"k��Ӏ}���)a��+��R(�!�V!�^C:�Ā[r�XL��y�מe��!p�Ж���W*L��>�]�!��~|<y�4�W�����ҽjF=3�p~䡇^�bf���=��U�d7.k9T��]F�Q
2C�S��s�k���{���s|�-��bEQ�j�z*���u�{��W���SB�-xK[
R{C�u�m����dx⛳�_?z4����������̌b9]� �aJ1̔ouiҡDq�L��+lH��`� �r��e���Y�32]PQ`4<��#���>�1d-�8�G��� �e����i�~X��D1�F�X����?Y��{����P&�I�Z�eȔ�t����2=��K9�9��Nwu\�,�C��(}�G[Ӵz6�Y�uc:kf��w�l��7�uu�)�|U�t5ck�l�3eK$k�#?�ԢL}O� A
$��p��}�;��^�v[uEz��zJ�]W�p<��,K�Hm�Z�纪ձt۲�^��YV���uG-���9�n~��3�����A�/K�����X
,q���p�-��hcs�zV
_����K�e�c.�ɮF�dY���	Oϣ�����V���'Z�'��d���-���P��͚���O?v����ۄ(�*)�/�\%��'���3��za���'��EEZ���-d�����bI��1u��'R0r��n~�}��ĭ����}��[�Rp����t�c�=�j󅗟? 
��^���Vk���Ca���`,�縠�NTc�.��4��dp�#��Z��<t�6s��ֆ(�Y��2.��#
�~jRБ'�|m �~�2�� ���/3  ��,HWG�E0�K�&�NL ��6D�+GJCI$��%x#a�D!�#��`�g��$K��X���	����Nz���>ݶ/K�/+�K�����M���J����(JQ�;�g���H�ň�'EsKR�D��Ht߰C)�@ÂH^�ka�g�9͂(T�^AG���tz�5��T���CP膕���gSD�0�Yo��<��,�#�t>?��L�%v����A͐qC�r�`�a���� ��\ ��F�s�S�ɽÈ���H���D^j�����d��[�$�1A�3�u5h6k�V�~S�c�˪8DϙI�%kd  8��p�p�t���2 `@)@4Pj�y
<�`EE�2�|m�Z}i���=��G{��WN���Z
R{���8�qc���K��4�l�:��_�ХB�X`�0X�!E��g�{![(�b�@��P4ɳ\H=�&.�ܙ���.�2�w/O��L���f(���	��7�:38]����EQ�w��l\MQ��eu��+.G��
I����!9�BT��<pP�N�,����fE洒������'B@9��2�:
:�(�}D,�͢��GQ�O�C�lEM@���_�Z���7/�1~.��'0WG��-D �  ���B�+&��Š-��~z��8��,��!���2��Ho S�P#F�xM�u�$�|~�R�x#0������`p�1SȄ��&^��������dz(�Ӆ���)��)M�N���'��Y6KD�@:�#R(�a/B�^ϻ����5����r�P�����2Upb����(�j��'����� �C
F��!������c�l���>���ܺf!��H-����5���:c��=�KK;[�λ,�ɸ��Zv�b �r��Z�f
��+�ɒ*Ly����$)�"��ɞ�є�ɸ��B*F�@^�{��$ �d�$@	�.�����̌���=��8��9�Hf�
�m��1	Q=��J@����p�u�.3
<|���	�i�F���Z�y q���1F�	�Q�J�Xaǈ^�����Q(�HC=�X�g�?�G�
܅@�_E>s "X�Nt b6s k�t� ������I�*0 �$�gd�@G%6R[b��EC�h	�$|'l �,8w��a�!�0چlB�!e������q["�7 ����Z���^�|����AZЩ��e! %"p��)��L��	�q�F�e���3YSȘ� ��T��R3]8��(��=`AF�� (!sb[.�wh��@��)���ɗ�F���\{�u���;�{��K�)� ��������i�C�=|���� Zk[�f�� �"��<�O�6�r��LX$MC'�]tm�@i�zF2b��}%��"eq����9䈳Σ>/=������X	-e\`u�.�`q#]cK��Ɍ��/ϸ�0Xno��s�<����1َ���~��AP��}#Hd�c���?�X{�&OƼd�$��\{Ϛ�b��c��X��3,�B�N1�*�sI��["qM�2�`e&K%p� &��Z�b�5H8	�H�MKx(n$���1���b�:Wpra���E3T@��rVCR�uphr ؁�0!�$Xz�`�7��/W���C#Ě8}Ѧ�������&��~��2��J!��ԟ&���|�R
܃��4���K$p�8��w��FT������߿���i� �_d)8H�Ma۶m������7������s�uls�~�!@\X�a�>8>��H�96��ebJ�����VG���x}����E�g������CZ�����(�:���� �^a��\�Jǧ���Ls2���f.�9�'�_3��
��c�3&�܈� و`Fr$�vΜ�@�>�M��ӆ�,�s��JE��Fb�Ȁ��	{�	:���^�<��$X� cP�9�����:���������C�0 ��A�I@�y�I�Q"S��\6*�����9�����H]�͢ �2�$ʗp�����"�z�1�28X�������
�0b�Rx��X,����?�� �2�p���|?rc(�HNF�6X�2S�TE��b|���+	�������Z��g�Ž�V���>v�7]�c!���������={��8z���>���u�H+x�GI�ԨӇr@�Fo:��L�F�(T�E�}��a�[���#�MB��-�>�1���j��� @���S�%=�HU�:(�$�QK����P�ODx-��a(�8�  �	�"a܃����"*^_��8���Z
}5F�Bd)t 8�"f��pi�N$�����d��O���UP��Wpt���dc�~$,��Yv���D`;L��E���G
��PJ`��Aq��,��{��Cy��p��r�@b�Q�X�`�e��˝:l�'��~�#$*B�A���U؞H�d�H��|�^���^�����D�Ō��gY����.)����f]0�9�6X�b�t�28�ؕW\��[���C;v�Hj�������4$�W'Ǘ��lg���m�u*8w��F�auZ���� AUh�h���x�xR�1����]v����d. P: �b+�و�8��jb���k
cQ�]US�������xNP�Ql�>�{A��HR��0t$�a�"�h9=ΦP�Oء���J�q�A�Z��<!N~�X�N��xfb	�2}�@�c֮�ҩ&��	������[��|����O~Ϙ��a�_�LV��\p���B�?�0�`���"q��0�N��@X�z��@���K �`� �V��,�v�=�ԙ�K9-CѦ�Ԙ�B �|�!�� �(���eC$�ː5k�  @�l�����ld�L	� ,1$b��.2݌��%�^W�N���B�H��mv�__5���ޱ�ɫ�x�$H���R�{,���l�b����^j�6ږU�w�u]��h����nu;�A�n�� D�
]x�>�zġ���U�D#"u��L�K�q���,�� ���E���8��@��@�Iv]O24Pm�͗��O�(���H�ꮦ�WDI*P��`��(	
oq�Ҽ�s2cb+�e��&�Y�I,��L��b� 6�:�,LF7!	
���\��)�$���äe3^v�%?��ĕ�`�ujp0��ȸ�)�m��� #���e��;Ov��ǜX22���h���|�DBF�AL�AЍ��F����uNɂ��e�<�������d����v)���k����c�a3e�B���޺�bbnn��qG����٩�ke���>�?�8%T^��@0rm��Q�B�l$?�/�M�O<Y��c�������Hgp������2 O��s�,,���v.	��&�r�kхҧ74ur�3�K$�s�nB�Y(�b=D���#j���u����p�C�����)j�
��#$��PۆR� ���
 ��񘝞��A�\<86��qI���5��u�fskkDQ24%���"QoCK]�!�����W�Ӹ�Aҭ u�X�N"$��L��t����2(�����s~�y+a�B֐A�+���_x���<��#P����DI����D���+��o"?ZƇxݝ)&Q�J�"��I�P�*X��{�S#�<[*W�O��8<2<t2��7�����;�^{�ݬo�:mzٜK�l�ȗl@N����+0M�4�M�0��f���%��,��@��4��p�B4�W��}�L��9��D K��X	�).�C�:ZbQ�l3�?�qæ/ݹ�߻����6I-���� �7��(��}���ް��g��ڝ]�(�A��VD����t:-�X+Ā1��e(8(��G�Dd��5.�(�q�����U�ԐDw��c����d(���*v]H�
�ah�Y��`������3�MNNΖJ�#��?޶���s��������K۝��V�]C�7�(r��W��� *w���Q_�R2���K�B�D���F�\g!����%+4P\�;�~����u�!�;䨟�_f���2����2��) �����1J�$c�T���$�
&"�,I�=��.��C	�J�[�"�B��myӢ������l=�~Ӗ���D]�n�k��g�v����jo�Y�5�e�c�c�����Z�1�#��844���������`Y6����j��q�\��A�3X��õ�, a\�9��� ��HpP�Tb�ԣB���/�_�v�w�q�;��䇮�����p��˷����ݻ׷�}�У=�/xQ\<{��z�`�n�؍����p��Y7jK ��|@��s:����J�X.��AӘMH� ��u,�&�������������;��*���tM��Fq���(�	^e%U���U-��p��]G�>T��2:����]{�B�{fgV���^٨7/�]w�F�C�'�)LЩ����E�����.�'� ���Q�=F�fKB�������I��"$Qʲ�Z*�gWh00,����8tfXf��cP*�<��O �L��'T
�\��{6+J���]���l�"n�Vd'�Sd�ADa��A���F?�L����es�l���Ƶ��T�b��_�#}��wK���>;{��۽KzvoO�۾������\h%44��E*�2<4�e��Μ=M��6k�UTb"_E�L�/�3A@� �D��6�3p�bg��ܮ��,Lc���FDz��tG�l�.�
�������z�}7�v��k����&���O�����k��V���g�_j��َ�[sSSc�N k�BzN�3:		�� )�DQMR&�\U���E���A��vz�`��
��2#껔�E�P��P	��B?"f㗱���<���!g�tE�5������u�3���������Ucc��n��,OP�XX\�_�4��q~aq�u�	�T�E�����L�l�q$�bAdY�a�m�碃g�&el���KUՙ���'�`�����U��.�(��I��g��wP�T�ǃ`+i)䭐	'�K	�Χ$��K��pm��"�\���{�1� �z6�
B���C�hGյ�|�p�X.MV�Z��h�:6[��=������(��ϐ;�C}��{����cq썷������uV������U!4B'�|��1 uN�񁥩ZU����f�n1K�g:$8��Aa
/�s�hX�lz}e�I�rb�Pv��130Pٷq�����g>��w.�ق���������v��.,6�8=k��uo�+l��iH01хvEY#>�2�]�:�"k 8c�\�B
���T�����#}#�0�f/� �RA@5E¦�	�K~^&��cP)�����(<�.�2t/��,}� kgg�n���>��f&���#�Jyzlt��͛�����j�gg��,..�4��
�d+��5Lz�:�u�:ݖ&�#��E�v(�
:� LH�x���$p�B�@&N���Lql���Y��%NL�H�5�|~�G�,�F�ق����y
��F"��h�H���a� ��:Г�J��� u�!��<ۢ$6%I]�r�r�<_)4FFF�JC�ɱ�����BA6ڥ��~������$ 
�S����/[����;�ںV�9���V�h�@M��6D� 
Ο=�:��3A�BU���8_�GL������%��de���dzB�m��F@ �!�M���j]�dU�G�����}�;w�z��6I-�_��� �7��z����f���U�0�.��LJ��4���E��Hmq	ӻ`&���N¡!l��Z��a�R�{�s��O
%L+Ȃ`�v?�K�Qc�БaD�P\ɇ��L?G���u Qo9{~�S�'kԃs������������'w�<��Hjt�zc�QnZ�J��l��Z�^mw�U�N��ԙdY1��%�T�Ƥ���B=s�	]�i$������`�c��S���̕�
A�e��yI���%�������\�15g)���6��+�G��EA�E?O���G��ӕ�������������B�4�TU�)u����|~Ϟ�I�s��N��)7��K��oow:W�a��u�J�X2��#��g�aBZ�9{�,D������R�DT����Jbd2�:)À�dT$q����H��<��E�dd�L��c��X��ѳ��=�m���o���>��i� �_��� �7�m�Xi�pd�v�U�,�(�⮥�Ec6���E&8_ g��p�Y
�<)���U��3�x�i���@4���L��}ޅ����,jG'��� �Wt�Ё���@���L�}���tc��+X��k�O�̨��I]7����cc����.lܸ��!uNB������Z����B��*/.,UZ�ސ�8UzD���Kv�[�axIU�Q�*ı�"��D(Q����9���BL+y
I��yH��Cb����b8&@��0J��LQ �D��= l�����MQ�����MÜ*J������j��/u����g�F�hU�A7�Y�?��G���s�$�����=z�h����e�*]���K�͊,�T]���$��aaa�t{6�P@Iȭ�]Q)��k��+���/؄{�J�I��qYbbp"+�ixa@EF��Y7Yi��TUT���Ѧ��?�~���m��gv����FF�t.Bj�lK�Aj�]�eU�'?y�G]�6_y��[�®��i�8ޗ:3�:��KT�n'�1C��{�����*td3������	�#���H
{^L4�} ��҉��5	�S��Z����5 0@F#��A�At�e���b��d��c�Fkjj�>55=+I/�3�W˕ҙ5��.����;��n���QdOl��2���k7��V�^�7����F1��S� �5��Q$�H�5�:=m:=H�y��D@;�����}�!�ѧ�(���BQ b��Q �H�`i�ٓť����1!�\1�,�ˍr��,�J��+d�V�T����Ҡuv	�..Ƈ�����������#��/��/d��Q��]ܠኡ�ʮ �8�7�xnvqqA����q�^a⡦(t��Jd^N�(���@ل)&��{�=�~� 9\1k!���	�RA���g�1�/�CCգ�b��M[.y����UWm褠 �_��� �����˗�l�{�V[='��C��n�=[�( �����!��I�Q�\��Y�\!�
x�HS&7L�H�1�C���3#ԏՀ�T�:��!0%6�Q�D��ߏ�����A��y+!ԫU5�߻�+��)@���$	�\.3N�s)u>�
!u��S�gN/O��Y3wn`hhzlxt�4PYX32Q7�V�P�r��7�3���M�'7�@��)���uD۲�VӖ;��R�b�e�n(��=����LC~�F�b�c%�{@�Q
���( �cA�4͈�"9RC�4LA[���h����ǃ�Bhd
��e�bY�$���[����w�w���x��w�+���ɤN���.�q������ڝ�.z��u:֘e�ʵf#ױz
����D7aR��'?&"D*����2�(��9^X�U!^�qa�1q*�����:p��"K
��ުU�N�J��׭_��u7\w��^�����~Ֆ���.0�����}�>jJ�|���s�#�W<���A�3x�V'g�I2A�Ry�:j�i��!
T�x5"U��9��<P��d���~�ȣjq�cX��&�|;`��=�v�z��h��
H#�Y����#��;~�a������N��%Y��~���ɞ�\8\Z,�L)���K6)�^>���Jx%�?+�z�;��'�'x�[�n�X$���7��ޱW^�/*�BG�[����?g:�N�^_�#�Ns����f�R��W�z~�) ����dr�>���|6�J� ��������4�क� �!�(@|E�&d���IIVD٦a�.��[5>���_�����J��S�uY
R����8�w�|��Gʶ[�O�]iܳ:���D���8�0DR_Q<�8�OF�V�,u����0��ז����`b:��0EO
YkD�غ�1�$���ԇ��\�/�����Ȉ��A��s`?@�)k�Xy�NBTHiˑdA�F"8%�0	���:={w���R��<q�hS��y]7jf6�T5�],��K���l1����������Ɉ�$U��!ѧ�(��k������ ����9��?yJZܺ(�)"-j�te��/��ܘok?����p~a��Tq\{���T�k�gYc�k���Jy�-S�4E�AR�x��ca p�`�D.U-0.��WB�de0l7�מQ�6�*�#��YL�sI��=�Ȝ/�˯U�O��u�s��jj����fR�uZ
R��)(��N�.��̥�����`8�]��#��'��8״��M$�s!�\{�Y�y�W>Ē��H��3۲H����0�gP �:qNV��_r�֖�r�ؖ�~Vpeԙ�|@���b��JH4,�&�H�H�[��E�_��w@��_Cp�v�%�pg�M:��vEIjJ���M�chzK� �Ѝf�P��^/��?�c�����݌�qL�tEA2f&�?�����H�홽 �5�EY�$q�A��h4�3� n)�'��עTP�Q���X���{��ZN7�:^��h�v/���2~f��Vŷ�!��(B�AW9zNz�zg�^%�Q��
�s����'"��Y/O|��j�.-�$\�p��u��غ(r�f�]0��)��I ��d���:u���g^,�ϼ�mW�t�����jÆ��#/SK��k)8H�ݻrr�x��}�'��h�x�����ƒ�s�3L"����	0<+]�#���42P,&],�� ���܁
B�R��L��:ֺ����*>�mi�˅�d�?	1�����;��p"�g�+!Ip81V�4	`�/��8�y|��P8I��ƔQ~7�B?�c���������C�жa��]��Rm���Q0 �4��[���TU��w2z�kf����Őۚ��%E�eI�TA	"1BP����T�~�v�T�O�G���P�&V��"�wܢ��%?2��d�/x�����B�p�P����Ǫa`xa�Œ�� �tM5��'� !�TUY`/I6� �hA�|I·�?��w]���Df���Hp&��&L�:Pb���c���+x�$��!�/�㬙�*��a�?)�O]���n����v��C�R�MZ
R�hm�ڵγ�Ͽ��W�}�yR���O���kK]�'� S���F��:������*J�u;@�8�N�
^���"�\�`i ���C���e��A�ѩ�>�x�8d��p���������J0�X���G�l�[�<�~{���(����
�8��:_��"��s��8pr!������v#�)A�!����&�cz~�s�=y�42���$R` �Mw���FB�]����"��e�x�ѽ��odzb�8�x`�����g�`c�'�	BL�%��P'�膠"�b�{-.�G�D8/B�J�!'��N2�����)��LfG,�TX�`y�4�Ha쏻��m � $z��B���fL�|i�R�{ɖM�]�+g߻}{Z>H�a)8H�6З�;9�J D�O�z��L��p�ݔ� � A`JtԁC)�Yo02!]�@ȐR������ԁ���	$2B�e�"��'�Zc6YQ�Yt�>��sj$P� K��-�AZ�h�s�/H������kP3�.�:F}~�2=b�H��J�/�A�,������0��������D���H����PJ/4��~��c�$2�E��@�ϔy6$0̩&I��ȅ���4J��xD�07Bd-� -�j�5��A)��Q>))�$n����I �1�d)$�(��_�(x%�qQ�0(����`���%94��TmF3���|�b������]{��殹f<�����Rp��Eo7B���hP��g�~&Z�n����v���H,��!��ue�{C���J�:�@{���lA�ÐI"'�,��B��!��u�D���0	|8��~�B��ك����ȉs�8�>�� $�^+J}��tU�'=r�cr,�%p�gt$$�6� ��$4�Kb���,2vY:I�
;��UI\1�9q������TB�y/\��{��t��&
���up�0�5dEf@��i,�(�{#yƬ� DB���r�
��}%L�.N6�"(�j�1����|.�w��կ�m��N^q�xm۶mi�AjoHK�Ajo	��lrr��(���\���|�:�	������e��d�:~Ǳ�3�X��Y���A�N��81� �m��0d�2�B�j��{э�(�ms�$_⠁u8�c[I��;�d6A22�A�]���#��5��,��x -v+�m�V'�H?��M/9�lFc���E�@�SU�Q���F'>RѰR�||	�"N���ؿs������Nv�AH����.@��c(E8�:cj,e2�����S,��$p�[G�ㄝ��C3 PT���xR�6	zy|5;̤����e
6NZ�D�ERTG��v&���u}y`�ŵ�6صu㩉�w��CRK�l)8H�-c�A8q����_~яB�fm~�%�$!�,��O� ��h	dj�q<�@
E
�Y�M�܌a�V���'�٥NJ  ��]	t{�b����}�|�� =�;��R�FՆ3�#���À��(&&-�,��I���!IWE�B�8��C?J����c� ��#��}1-���Iw�ò�8QQ��r0����M��_��>�0G�rNc�U`�1�(��	֞	�''&� !��n)<�2 ��N<�x�|�E�B��}.�-`�M��(�@;a����H@�`���(hV2X&#<���^�PVTK3����ۯ�ځ���[�l=r��k��6X72���R{�[
R{K�ƍ]
���ҷ��1W�W}��T���4E��d�n�Ol�M�8�E\�&m242Nt���ɪ*i�,��l��8d����(�z��:�`�h�Y5�u��ӳS�L���%mX֍��Q�A�I�	u���]�F!�g*|b�S١�2�ٞ��� ���1�:���,�I�o�#���yZ^�����z�s � ����M�Йz^��-�)�@Τ�%�;h�G�1��������/�B ^q$1��� �{H� ��V�8)�DD���� ��d��Ь�4�;q���  "�\����,p��d�#��N�$H � ����J�}_5�N�2pNW�WI~q���/_z����.��ذa���#��f����3 ���;bdK_����K��;BM�Ա:F�,��s�4K�e�4���QZ�즙!9S��*�Q̺A�B�G�N����<p�m�Qr�����V�I&���ꪫ�|w���C'Ol>vz��^���z�J��.�[���PԦ�+c�DWT��:�υ �	���ʍ~�18meJj�A�\�cR�e{�"�r�?\��'�"p�B_&���'�� �dp��Ɍ����m%N���;������0�>�+Q�'oB�l�\ւH��ˤ͘w��,�D��k �[Ʊ�$WȽ`] v s"Ũ�I�)��2r��R�����J��v^~b瞝s{֬qӮ���̖���ޒ�{�n����$M���>Ys���&_Y[ZȐHM�@�}�����f�x6h"Xdpp��J%��((0���$�5I'k���&�N�t0�H���Q�Ѷ��j��mo?r�������ju��;/{�+w?[�8�����]@l���U�n����(0��:|Z�C���0B�G��W��!���[N�*�
��
lDrґ��Tٜ�dAgJ@F �R����숳����d���%%N��l�d߃�\�e �z>�&#�]�3n;������jD�0��+�ā%��p�0P��	��϶��LE��������v4U�+�Kg��b�������u;v�?�g��j�v�X
R{�O�.��{����v�?�i����lw0}YV�L\������F������.�暤48L�L�h�N�b��fF'fS=  p4��5�T��{���g6�>~b��Pq��m;μ�ګ�k����k��ӓ�OM혝�]��y#A��i�1hFF�� E`僤� I�G�\�fB�s�W�;k�v�[�\���ڡ}O���1RL�(�9�g�-a/�C+��5��!�?(Q��E��DD�l�A����3"f>�m���?L� �r kL����B>S�����["3������Me��S�b������5��\5<}�Ƒ6d�Hj�]d������v�m76����z�~�����wۖ=x��� a�<D����.j��g����H._$�B��fK������LK#n�H,�z 
���M_�̜�;�	�wn�/.��G]x��g����ܸq���n����v]s�e7�z�Y:wnj����湅�M����:�AMQ��4�W (�lG�f�t�#�� X�Iy̧�6>���~�!��&�h@� p�1Snį��H��r�?��j���|F�� ����h�\�aXi}���t=��4"r�a� �P����XQ?	!zD����d*��f��Ɯ�)'��G&V�?1�v|j����5�<��.fK�Aj�Q����C����^y��s�oi7[���F AL���4i� G7�N�D=�>��AB&Gr�.�>�N#lӌ(P��W{g��u����:=�}%	B�\DKVHmVb�q�T��%]^󚪔���#Y4c�")	� � 	` fzz�rϽ݃K�[�����V��������r�v�J/e����� z��(�����k/��;U��pza��ɹՉ���Wοt5�����vm�pfc�ɩ����ϛ���0���X��j�U��F9pa��U�Y��o�ͷ�˵Q���`9�Rb}�9O�W���j�����%�s���y�BiX��7��0T�EQ]�S�:
2�V��;,��G(6�H�ui�2��
�b��T*�dE�U
��ch����Ƚ���ۍ���Ϟ[�il����������
(�dii���Gŭ��T��{�?��������K���C"�i�,��}M�ҘP���.K���uۤ�9�a��6:�6Rs&H�G��:dŋ��Æ>�L��,��Q�}���N�6=4:E���W��wWV�,�l�l���X���||lf���7�'�4<��ܛ__�x~w{w�:s��� :4�ي*��)�y�Ōr�۠%]���?�̳��]q03�_�\���� �|�zc#�W�� ��E�T��  gBe��2� "��y4�{.ݒ���m�<�����"�n�X�TҌ}�V_�699qk���G�ss���Ў:ީS$EA�|Aq� }��4��݃�����c��:8�Z����I�Fu���}�y3#$�J�i��:�]��Z�Ft�$
p�*��a��ͯ,��N�}���	T(ص��]��v����1I(H�I��|���ѣ����-�4vk��6s�ģ���'/�}�zI��������t���*>N�ۇ�i�N�E1.'��$� ��"@�d%�W����t]����w@��b́:�����E�}�b@$�Y ^7p�Y8�/QG����YB��4-�<�2��"@���#�-8��Q�sfY֎����������w���t�j��IY�c�� �n�� A>�w.���`����ۺ��z����OeM�~Et1�f�(diH4I#isKah]��T$У��2�V�>Z��:	,*L�b��P����
� f�IJ]LӀ�IV�4�iqjE���J>L�8��8�k������,;�saK��.}_d�F��Իã�w��F��w��q/R�1D�����մ����e�Fo+�oEeuն�X�Ų�A�H�%�'&J�����T3*g:���[du�l��|�}+\� ��<��:��P���Ǩ։��(���گFG����wW�\� � (�P�m���[?�k��k���󶠨�Y�;�_(Q�6:)�~�#�u�6�#u;��.��VV�&&=�FlK'��i
C��0ӕ:�}_"4�s�!��̀ )fYb&ad��@L��ɜe��s��^����v��w��� �^�J�o���V�)8"���ҤV�`�N0����Yf�[�7�;!�硎�
G]��w2����h�<�V�Rok�~e�<^�[�:2�v��?pTA �� `���V��T��<˖�����|p�o���W0C� ��������J�������W�޸w��ݎ����'I��{(��,*�a/�f�U���C�!;�S� ��m��N�`�2���Og�-c�z���bB!�" & &y�
�D%!���,�U8�h�i��$rq�C`����
r���������fLp�"��a{�VAR�x���M�dèT��(q'C�uK(G����N�������-fi��'��?�	U#���9n�6�s�C�el��pN���q��
�Cz�����߾t���7.�q�^?�����Aq� _��%!���ɉ'�W������;�?�x�N��ߓeq2�B=
}�e��
K�w|* ���#!�B"S��v�,�jt�kY�L��,�İ�x�-96��>�,@d'�' ���| �(&**�`8X��`���J9�*�܈��޴ǜO�����A�X,'�	 ����1{l�
�:��*�rV�,�,�P���>APmT� pyUe*�Ǫ~�Q�N�YJ�(fߓ����న�0�{�"�=u]OfǦۖi��u��/.�� D����S$�l��iP ���f�H���˯>�y�7+�>�v������a�|�����'{�K$�J�n�Q��N����!�!���p��˶��A7,^4g�Ā�*,,*��/�B@�1�c��F)G�f����@0�R� �PN�b8CЇ��`���,���s%"���]��D(x]���l%OX&���SpU��������2�#���VN���Q=W�0aXΐ�� +R
�������14:��C�E6:�hS��ЮY�����w~��͡��I�� A�8(��H��օ��k�.�^����~t��ۇ��U_ee<
B	��sBlJ��o· ��g�#A�#�e�����D34Y��U�M���*q��l0��}�(������	��@�20W���$c� �36Ȩ� ���3u֖N��%�Cbu�w�4����&F�q�U� ��o� #`h:�~�%1�I`NEe�b�E�(3!�Y����!�����P��9�l�i��#*��_ZZz��Ko����M��}� (�Ϥ�$�ip�~y���G\��͛�����[����x�u*
�"K�$�y���4~+u���O��� `+m��[��Z�>oJ*I`h���H�>�i9Nl��4<l���<����V��X�j`s5հ���~U`Ȃ�(p#�2� 6��3 l� 
�r�Si���D��,З��0U2�0��"Q2�nlt�M�`��$*���f�~����u�N��|�pf���o���3mG##�_��)3	-8���|�|�����|i���9�k���d�����4�{��F���d�it
9�>��`���U�ي�@0�=��0�X���R!�*4@K�HT&
zu�DBR�CKC�n -x�#�N���;�;����}�Zv�y9'��-��>�,�����q)���oC�["�{��p�f�ES�������j����q���3�7Ϝ�v��W�g�n ȗ����g�ipl/�}����[7�x~�����{u�<I�_��<=�"Q��ދ|����`,4��5�tUs���ìL��?&L�Ⱥ�R�UA_�G �[�Խ�M�$���X� B�aJ�h
+��C��f`�u��R� T�vme�K1 �sl,4��`��JQ�3!����w^!��$��=H,KAʺ"Ʌ�(9D!D>=�X��`ll���_X>}��{gΌ�{�b� _.(�K�Li�h������>�y������=h�bX�~Lzݮm��z�^z_Tu&�8#�����	K�glN@�Z#��2��jEل��(�Z��Yʿ�8��ΒB�|���#��EQ�tx_^T�N�Y�c�ꏳ����^�}/Q�uI\�"�|�UP��9k}��
 
E�m��ؖ�RA����]Ǳ?>vl���������5U���� A�:P �WD������un��f���[�y�֭�6����Zs�j�� jgI����$KX����|D1���> � ��7�X�V����X�^�_����A4�$��C��{>��9!V��?���M2/k
*#�M����!�w�
$�kU�gB���,����k���n뚦,�>v�����Ϟޒgj�Sg �����)W��Sx@�e��ym�ƍ�߬���=�8���qoo��9�}"I"��%
}1�A��e�~�m@�GÉ2PT+v��:���_;PM<(�	��d����.���p�����0�P"�Dx�a�j2&h$fz�I�*F
��9)�a�i��a�͚S�4-�]�oLM��������\{a�֦�0C� _/(�k�r�^ׄ��?\����hd���;O��v;�y����t��I���4S�`�#�l՞�$�#�����h�"��d u��P���	e" �f����+�e�{4ܴf)�4ǜ���Q�p�
I�⢮�9�(��ȚѶt�P���F��v�,K�r�ݩ��OF���������	� ��uAq� E��>��q��qe��cs�`��������v�D���h*��1��Z��J�J�%"��]�&B��4����J ���@�� �T$|�_��b�O�`[b5K����"s1�d�iY�sA�rU�SYSc]3UU;�,�jVmۮ՟�굍�Fc��؟ԇ&�ǜ�;3#Ƣ8�<)�A�o(��iA��	(f�~����Z����[;pg�v[�;��I����n�7�U�H�`$�Z��zc��TγL�8�E�� �m��)���A�p���
P �E�/��R.IBNϠcQ��TQ�D���*���J-]Ӷ5�xb;��e��ѱ�F}�وS�n4��Ԕ�LLL�hN� �lP �7�ʪ���F�Px�I��ޞǾ�
�p�5���3�{^�u='�F�cQOdi�"o$YV���L�L˲La������<
�{B*v#D����$��51}i(�����+�R���C]�[�*�����ul�c5jm�vZV���O��R'����X� ���� A����)�,�0m�)!��PX_'b�)ݜ�^�i�~`$I�t<5H"�
5#5ˉ��LE�6�9��B�B&JR�(R&b,(Z��R�HJ�(j��Jd���v��1��($�����d��y���k����R߬<*`�ޭ~(�B ��{��Ow������?�s�9yA>� ��� AA�P � 2 �AA@q� � � (A �� � �8@Ad � ��� AA�P � 2 �AA@q� � � (A �� � �8@Ad � ��� AA�P � 2 �AA@q� � � (A�����}x    IEND�B`�PK
     �8�Z��[?:  ?:  /   images/b75f5fea-d559-4623-b1ce-f8cd504066c2.png�PNG

   IHDR   c   \   z�   	pHYs  �  ��+  9�IDATx��}xT���;��L&�B�P����&
F��"*�(MT@��T� H)ҤI��e�L�����������{AA�{��s�d&�Sֻ�Z���;l���/�������Cd��!����o�����B@�����b)0~:xrU��|�(5�����r$���������D�ر#|.�b�u���6}lZ="�����_
:LU��
�ӝ�P/�����:v����h��N�P�h)0�vN�/��vOK��oc�ׯn�߶��e�0��)�
6�R�5�K�ѯ_���+����ß���o�?�Z�N��z�&c9n��>�|>p�\���/�"2�O���x�S��4�y)B����]���`s&��T�A��P(��������-�C;d�4�Ñ�fee0ig3l&���3?��|�)<?��J���6�ߏ@0�-DQcB�_7�|'9�9�{-�|.a�Z!���W��$$G����n���p8���C��I�(���^��
L�:��ixa�Xl�q C�z(��C�KKuHO�7�a�nTUi����2�o��d;Z҂����Ph���\ZQs~��i��[z;v�u�7��O'��^�~�zr{�����s�.<��8�|�<9n,&lV�z
o]$ �y�}���ȉ-:vh�5j�$�8����Vt�\��QR�yΫ�4=�����s�E��+��Yѱ� �;p$�K/���g<����?��
0h��^�����+����B�j7�¹����;1~�?�8��X$�HHNN8��,.��Er��� ��1p�#}��A��	�\����(^~u��d�6�qV��ڵ�S|�d�:.qw^���fMs�@,^�^�5�Oa:+�؂��YN�A�9�E���b�蘘~=z�y��ɦ��7�
�u�����!�B(|��D�hߡ5$�wg�粚��������#�A���x^_������G�Ց�_G�ĭ�ܥ�����'�b���<���?��G/c������	Dx��W8�N{q@��#��}������S�9�x�X�0[Ⲉ�)��
M��K��y�,_.LL\���S��6f���£�����^g2 ��@bBBv��i|����'��1���+�=9vj����k��	�O�p0��ъ/ѵ{�3�_���?��3c
^��l��.'�����|.�"%��~-Ij%"�zE}K��#}$��)���=~⬠��2?R�Z�b1$a�� �$�<=�8>>q
�:._�"&.i)�`�C�Fm��}Fh�4{j�G�ݦC����ɹ3����?�ÉY��F~~����L��������]v3(�DH���C"�@&���(��[#IV&�EYZV��y�x\��'�'@��i�$%'V{=~_��<���DNz�����ı������V�EYyLf7jJzJ<�����+���'&O����S�<�O_����:z�����R��_yJ�T�^��2��TW�Y�V�fL�C] ��(eb��V�����0����sX�R*���%X��d�ec��?��ӗ!��^�`0u
Cc�d��'�BL|���A�vm�Z�y�t\Vx�
l�4m����)/ݚ����K��|z�d,[��Z�C����b�·Ah%�\�>�=2p��a[j77��6i�q�|���$���a?��?���WI�����0|У�w>X�O�pz,��� 3����I!F��qN�0�B���6m�1���6��d0.��~��BR\^�Ӆ�9�Y,���6�e�ƕӦ�  ~���������gL��P�C;�g�!<n�\��v��N��ӒѲe��6������w�&�y*xd�|��*xJ��OOf��/�ӭ[7��֓$φ��ۈ�{���S��n�����O�KĐh�ȡ���~ϑ��&.�(ùKWЮu�;Y�j�>nҤ�aÆ�ێފo7�è��>0_=P0h̝�>$2)�ݽ	zv\�v���Ԕ�b!"��@�G�]^+�g5�N���������?�5BSI�9wsޞ>��������"<N�-ě�|�N�a�E_ ��@z
���|吁=�>�jsrtT_����k�Ж� `�ի�2�F����~�h6�G>���
�W�C�V-�i�z�l��'���f��#aGB� �Sҡ��^���F��JV� ;8�?Z
yT�=]S-#��!�e�.��μ/ӯ�"��Е��E�������5[<z�?�!���J\�)F���,+V��j>9fTϋgι�|����z�/����xD����y<�VW�B�h @(Hoiݲ9�S���h�g%'�����6��=zv��w���	�"�D�T�f5� �LޚF@��L�/�8��CL"y�o�O�xj�䒊ʥ
�$�����(B}Sq�����]{_�TU,�}l�����&�����X�v��l.��t:?�h*��f���5��DBz#h�4'��G���7��j�e�7Y0�H���S��fQ� �������1�� ,�����m����6��?�p6b��v�-��t�:B���Rn~�w3�}�H�`�/�Za9Jo^CTl�6�%����~�D?�&'!�qKTTV_K�U<VVg$RC�^|�����hg�9��׷��'�N�"�3���B�9D��Yp�|ϟ>�<:�s���o�^w���r4�ʀ���d0�<y��	�ť��j��i�����Oǡ����6�Yo����!�w�����n�>SA��b��1j4k����j��K=QU�����c��S��>� <$M$#�$�.t� �'�g�=�����p ����Ek�.�R=����Q��~�V�
9�^�AÆ.;q��-�͎�m��S(9	�n�Q�k6t?�C�ˇ�_1�2T�2Η^z����W�������F��-�7�^��i��]x��A|�v#��3�PBZ��� �����gv�n�|<N��n�nrL�8A��*���p7	r'��NȢ{�-ry�kEvW�⊢'�S�B啕Od��C���8����ڔg�=r0a��_���0~��^�8r��\�C�h�ݭpXA���_�?�ʗ��6m]�E� I�zEI椁�y�Ӕϻv������B��C1�;t�8~��o�#�a]���� �#E�q�:{� �bb�V�g*����M̗�����!&	O!lt2ǝy&a\,.��Ψ�bΌ%��*o���I�B��z������<��_�{���k�w��vo��a����9p����YP���xm���gj*F��s�EQŤ�i�2� �� ���7��$O[�Tbwy���xg������l�
��' �p0��=H���@2[E?���=Ϥ��[��_�7@drLZ�`��ֲ��V$gL����Gz����c����l���y�f��ٹ˛kWm�����E"I&�'�����A��WbR�n���ȟ���{Og�աr���9
u�&]��tz���k�ӄ��N��;��1����˻n���uP�kў%D��wI�JR�5�E�z+��2��J�g	uN�+*����}��Y�-��Qs������ѫ��[�g��h-N�*�'ʫ _F��8�������nL�y/��t�B����W!�8Hv�׮}���iߍ¢���m�����jv~�a�gC_xi.���p?����":���_��_�|s��Xz��U]�
<;�1d��º5[�;�f���6���H�8���{�?�<i�e���/��h��a�`�^<q�ۊ�oU�z��*��jX/�3�.}7�ÖwO�v�h���X�VP��A�P�(�g�bQ�����zGX h����%�;��>�X<���$)�@`��'���`0,Y��¸�1a�H��k0h|��<�-o��W�����>yE��'1��q�Y�+?��`������� ��@v�&(�q뚏ϙ�c���v�틝I�_���oe�B�!�cԛ�\ۻ���dy�UEX��_��X|](�.Yd����e��Ayo���t�P^S�H���8���w��,�C,\����M,R~���3.>v��v�:�����,�sv3�<Ѽ���co�����iGii�ӓ�[���ټxq�&4�KD#�{�]��g��ѕZ�윋Y�?BN���s.��\���B	>�E(a&��#._pZ&�O�X�+ʞz�Ѥy�F��p�!`���[v�C�~R\f(����1�a��Z��I��5��{�]�{~P�H��J⻗0�J�����\�=�L��A���q���PD&�թO_W��+\6�q(��t:���[v�}�һa�6��k0�d�m�X0D���~��Ǣ����}�[�ǿ{��ea0����C{q~>�s�H,��eEt\*Jjo��.m~��X�ه��׋�D2ѳ�/���s8�� ް��Z=Xp� �����-խ�*L!O$��&��e�i�����9N3F�p!8�3��:��%Z�.�����9��٬S|�qz�EAtG�b(��/\,����}��]L7	���tw�CwY/�k/=�8F��CM<�n�������Ջ�r�������sH�c���tUDӖ��^x�'=ӊ��="	5@��|��u�/U�im ��C����Q��`S���Z	���m|��l���<��;��9���i����!��Hh���Ʋ� 5����L*�L'o���t���`�J�"�V����2{���N}���B�&�r�J1 !S�H�jZZ涱�W(���z������ɍ��8$�AzDZN1ذX��ϸI�	R.�����^�	�4��:�^�-&6�p�����Y����\�g�j��
��H�����V�fp��@��B���Ù������U�5iS�b���@g%ξ��?�����`��a1�iVTEZ����no���6	�[�qK���3_�nP� Wv������l���$r��]���OUE�U|gFyi���g<��=�2�}��ؔX&&-BjAe3Zh>��Qt�<����G���B���=�%(/���I��uQ'6����,�U$�*�q�ڵ�?<J����f^����H��Us �"/r�L8���jy�Lª� l����/<�㭡M1b喻~�L}���>,V�^*D6�Le����ܤ��I}����`&,L,�b�Y���¨�3�I����)����V�^$I
��j�������=�A��Tb��L:?�\��ߴ
/_���O�0�.��1t�����3mN\Nj���GKd*a�v�B���q�%�^�#H��aܩ�"����%���9� �y>���݁�9J�tĤ�Y����|c���V�ʅ賝�z��!�1*�zpH��^�\��[�|��v��*6�g�;KXə��O�bc�(�)�fjpP�p����.���m����rȜNɤ��ʗ'N���a���ta��z�����&�S��NԠ�~:L,y�c��a)!���i��u%�B$���n��u<��}�4#�cH|�8�{W���B�iS�V.�<Q��P�~�"�R\�Z�T&G#�ɂ ��x��:�:�$H}q�l["�%�?�|W��?EW�[�fx�A:��I�m�N��k���N�;G٭6��\�bb!��$&A��7ۭ�L(Zaq�F�^���~�m�K6~��P[c��ڽix�d\���a�������F	S�V�۸q�p-���Q6�S�$��h��K�!�ӑ�vI�Gn6��}�쿎e<!r��`x�$AK��	56�����c�x�Y:�M�`!���f�|uI^>��Ń]}��2��J�띞 %w���Ą�;�f��~,�g�#i�~Z �px��㓒od6ju��U��/7p&My�!�H2h�DE����e�Ux�Ib����>�'^_��C���{��^���[���!!3���T���W�%�h��m|bRo|�b-�N2���HX����Z?���{���>A!��R6J�1���2�b��c����d�$��իp�D�b��\��z�ǂC�"!��	j	I(2��*&��. ����	1�Z�t�ɚ����>��~�	�=��];B��/�����T��\�/z���ZÐaCw�LK���G�',�.���`0�oւPz�f��H��ۼi��O>_�_}�`���OhGϾ����lSC�i�ఄ[�`�wm;)I؄e��L*���3��\}�m	WxتT�R�~rU���*��B$e��R&W`�EZ��dXw�}��w]���j.܆J���Y-p���������B�a!�g�OP}sVke�{�m�g�X^�����^�YSU����'�#���uGu��u��П���e�>Cµ�>_������*��������	����alEyE]IE%2R��Qj���"��iq���ҝL�I
)�Fs,��IK�L*����[�;��H[w����^�(�}e��PO�4�
�x1f��@%bPmA]l��#��Bo�0U@SUb2m	X�)8�`���j�7�3H	�����M{n�F>��x匁`~s ��}�Ϙ���	�ш��˺��m�S�֭�8;d?"
£��p��.�� �m�Ʋ��z��0���B��`lIBUݕK����{c�G�!�q3Z�]��D�!	Z8x��T")�7tF	]rI	M%���b��]j���W�����Yj~�����i� �z�@���.9
�b���R=T���$I]�CuM�l&����h K_�̨u�+$a���)��Z����fU�tD����&b��ױ���'��k�.��E�,�A����!%)��`�;�{џ	)��Pg#�-��U�?1B�G��^*��={�۶zp`�P��?_�'an�8\"%��H���-��r��S���{�<�����fw��e7��1)�l��֑�e�^"���A+��]�pX�DX�4c{��V	��j	H�#I��U�^S��2���F&��vȢ�h���-��C4pPL�w����hHwiL[bd��i_l��e۾A��d��z#���g�S��p����v7�RZZ�z��&�,r?�������<���¨���/�IoR[���cG}�t�ŋ��*/�r�,g�T$Ngg�%����$z��p��$V�͌H�L�f�:Z-����a����'�ʆ�<,���4��2��'rW���n^~�R��LC�u5�z�jL���u\I�jx�lpzp�I�K�Í2+���L-��n�U��~J �8�@��(s��E��5�/�w�� 5-	b���a�L�q�]1��Uh	x�;H+b�L&KLzn�᣻��y�`�}sk�،��F��L�y���%E(�b�P��ls�j�����`�t�=��$�s^�Q�y͇�aH�����1c��O -}�s������._�XB��6�����CX1E�!�I���p"":2�4ي(l�v�!�B��Y���٢:$Hp
�IF�{c�$)����/��Q�X�X�5f�X:p��)4u�(:gPɠ�yv��Dȇ�Acb2�V�%����?Z��}�m�'����牸�P�$z҃|=����:���:���J|zx:HB��>��b��P?)�f}� ;ߺ�#H�� �b�bUR(�R�j�Йh�z�����ȄTIE4�R��+(�䐰(�U1c(����u�!�(ᗩ��"�!���.��x��h�����{z��o .J�����a�D�,.�������+a�p�l&�E�g�x�y1Ez�c�������Gyl~��v��Ji��wI�'ظB���op��;���� EE�hu������#���^��'b��<'	3V�J�]%�	)�F5�\�h!�qIⰻҊ��r!]eb-ը���Sh������8�ʊB)%���&�HhIQ
�e����x{`�����Z?�_�1J˫�-s�YI��b ������`%9Ҭ�#퉴b6�AQ���=E�{�{�N�YV��F\�]\Xh1�+c҄)Y�k���c+�C�_���@�Kh��t���pf�c��q��hk��F
!��wϕ���`��M�P�������Pcw�Q!�sB8\�MR���!$8�()+'N���������kG9ņ;Ć����Z�I\��d��a��=���:����RZ�<.�&����$����Oz�1Q�I�V�a>=�%�˙6=s��p�l3Ȥ�ͽ��Z-ƹ�ZL-xғ���Ϩu5�%�_�P7���Ev_1�py=N�R��Y�D�����	O'�:�sul|����"��DoAb�L)f�����v�� %�"�nGF��p~��|�r��p��+F�h��DX�[U(��0uV%��ѾqΛ����!�~R3���b���Gp��,�p�b�P����>�^j�l�rDGGB �x�n����j��E|<+�u�$���q��2.�|���qhra���f�^�7՗?t�MH�n�j*_�ی���њ#�#��	�)"w��jɊ��E�^���8�4�"��=�&�W}�����vo���]�Kk�:%B�"�M�V�v��b�,�"��0aN#�
uxQM�8!��:�j4�Y9�v�
�	
<>Qq�{���	љc�u�$��bG�7{��Gr%�[}�z�iL۸˟��/�u�scp� I�,f�Vo
���FD"�"��O���K�8BLn@LS����L��N���K~����j����^��w�)}��sbz�hi\�a<��.V䅠7�����K�GŢ����*��#g��l�|���ʼ���^��oﻈ-�N ]���m�A�\�vc����J0.;�a�Fl-g!M�ߪ!ɽ><U�E�  .*6?[��M���q�ԍY��C�9+NbK����R�ښ! ���"�����w�+sg���?kc0���;�$�ED�2�Q�6��Ee�m�B!M�J("�̓#'��I@�c?��*պ����l��":a�k�G+]�M=�g���PLf��:VmE��ÆǞ=�.��?�l��7�>�Z¤.iu+�G0�;'���˲��*�6 C��!�"�1�Z(ak|.l�W#c�p��Ʃ:�I���ѾQ���YV,���c%Xs�67��=Ukd�m,�������a�8r��͍��V6!.&ɕ!"��$iw��R\|�|fz0`��,�a���m����Alr�������k�R�b#[�z�g������ڠ���p��62R�tm��d�wr�=��|��:��:cю��lZDGj�l�r+c���ؖ� �nbI�j(]vp�n�#�a2����:��[0$#<��kнY#p�A��KH�n�!�r\�YPcwF���8����e��͛���yV�=�民|a%Ąh�-|~��j��M�0>�����)c��s��������|���5�Gx� �YsJZ�׺������<k��]�ǫ��c��Px�<Z���o ��za��w-�����鼯�y�Oc��Ukga���]���<�.c�Ydd4�Kc�Ir	Mq8��p����v�g�;+3�@�	���l*n�E�Fy��Ew�d��J�ޖ���Ȱ���hۋ8�� B��z>�YeӧLǶ/?�|bb� �,���)���bb�m���U �βUhٺ�QqkL���ZMmLbRb�/55ÅA�j��7�G�k�# �v�s5��=y����s�M-�������Ò�G�Ѯ��TW)�T���)-[�n���h�(A��$�"��zX�(ԣER�ݺ�a��лKgD�x�V����C &���&GR�f鞓V6s���o��Q�͛��|�7�_v�٧�N�#�;ag4|��l&��}�>��@(�+�ק{
����6$<v�wO��]`���)2�:Ԧ�g|VW[�fNl4"��\���P�A����jhh�:*�ź�s7�r\^祉�}}ܫC�❝�0{�&�5N�j"���ڶ�!�i�9Aɓ-El،NDŨ�L�}$�n.2�ӑ#A��
.����8"��������J�����=�A4��A�zx}��chܸY^��oD/����.x$G�X<o}����[����l�P �õ7N�>>�ۃ��ߖ+Ü7?A�.]����������J�RS�2��?3���}bqؿ��JMu%��-Pr�:�������O�x}6^|��_=���m���g����@��Vr��6W��&%#^�vXI\~�ȤP(���2��L>j+o�d�W����������{,3-�,Y-��S��~��=z���3g�����I�;�<2�<\K���n�<��Z���J�(u8]�a��Z�~'�������ٟ���}lAҒ%����1*.�MM�*�����f�t����/.+Fn~G�b��GΝ�����gK��������{`[���N"��)�$*g�yLo�2�R4$������B����ό�0�I� �1�w�bqI�O�I�8Z�)�ONI��o��`̰_���W�����p���}�UTԀ^��w%=C�VASW��ѾC)���D�D�XJ���Pώ�o^+�F�N�Fki��`�@,^�1��x�i�:v:�������LV��aalTt�VWy��ud�e-�z깦�����{��5F��3��b��^[H��VZ)�@�2	�.�Kf�$)�p�q٪H�� �q�����k56z�=Q��ڎ;	6�	m�r�3�&����0�R�PC/#�_�q{S��Oh����B���[��ЉX�F�k��}y_X�:�q��<�|���^�v֒���VEE��z���H@�s�����Q��W��O}��곯N�s�f����K[�sb�ݢ�����d��~��`���[T˳2�c���JtKSAt�����T�B�cK&�߾i�YP�cI���3}�|s
7/�_K�~��bB��6<�#�(����ʪ�=٩I��z�k<&��B� ,�u�RqŁv-���^8x��{��}�NT;�Ő^�h���v||�lMyɪ�7��,���.㬨�D��t���8�w����.���+���}�#~��m��~�C�C�[�X��qʡ��tO��*dX��2�HF�FrDHEfO���,�Kʆ�`��@�v���>�E��͛d��r�<B,�R�[r�n�V��d��Yb��<�9"ݒ������kX��ǿɏ�m�1Ĝ��)>,�����k�3Ԍ������bUuuȱ��P�aԵ\���v�@���k����=��_=���M@=���G� N�l��'���YCbUqߏH'�oWp�H�~bv�py��Ħ����	�б�^Fp�����bR��PH%O���6���* �����녫|��`�����(U�=�ñ=M��k�I�����&��u��>�����f �c��߮�<�l�v�UG���
<>�e%�NH��fa����C�6�/_�����|ه����J	c���_l�O�j�^/.�Z]c�s9wX��T�ǫ�e��l���h�+�q�wm{���'�AM�V�ע��J��J2ӓȽ��,)���`McJ��J(�bw8�������/������`$%���B���,���9m
n^<{��dDDF���
55��IH iU�S�?v������G�w�N��ק���󤅶����⛓�ݱڼ��5��ݿ��^�.a|�sPg>�z����~W��w�^�~�5��t@zR�c�Ed�у��++#��d�QTQ�d��ي��/J�"���x��t�<t`;��؋�?l�����;$t�k�/7����
ж}�ʸ��ᚢ��L{�R�@IE9R�Hr��̱�h�x��ė�����8� �����`�)��Z�;6��C�0q�*��e�j����𯘇���}�`l���y��{�����ܶ��QҪ��闯��du�ws L�**7<	��ǔ했��V���];��Ը0m�����-�| �U��K>�
������_��j<DSrc�,�s�l(+-AzF&# >Q�u�h�ǵ�_�����YPZQ����G`��I�>d��^kb�,>q	�:��c�6B%�mW�у�����s�W;p��Y�(��{��g��ӫ��۝N���@�Fo���6�3�DbQ�"�^@����dx���s�?�`�F���%x�h���������۔����
]���"**��tuLO�?s�]�Ur���/>0�[o�t�8���c�;K����&M�y7�6O���
*N����0d��<�-�"Z)�h��x~IEŔ ��
�f���*���l��O(�6�T*����l�h����;�̌HII��>{��M�@Lyi>>yo>���Ԭf�+�ontY��N(���������
Z�o��ux��{t�]&���å�����;����R��r�zt��+\=~���ź�����a�p��mrZ#/+��7�F��Q����M�8ಘК����p�ܣ7z���"�<��_0�1�~�������8y
���/�z����@�x�]|�h>a&�Ҷݻ�9��O+-���%�j둙�edj*K��3�4�����9]��=:t;(�J�&F�M���)�yS�Z�;w����E~~>�t�|�b��B�/W�����ؑ�z��,z�:�u��K����\
���GN���-�!&=�Jo�ŪU�6ꩻq0�#V�Ȕ*}� �e�Y��6��ӧb�s�譙��WȆ�,z����vlEy�mӥGkߡ�5O4�i��]D{4i���:��z܈P*@
���9=�t���y��E�}r���{gk"S��c!	����es�C��=����vPX\��_��~�����/خ{���˫���Aޕ�����#���cK�Oz��։�l�z�D*eӳz�@��/�Z�/�=������-��~�öR]4�l�q_��cƽ2[Lo�hs���()-k�GZx��l�T��X�&Q!�Ŗ8�d�ߟdw{�s���s���Z5oR�f���v����d�Xl]���()��U�D℈U���~�8�QA���œ^K��+y��z���W���+���O󤪮4� o���1c4���ƳS�`�'K��M���E�i=>��=�?������Ii�n4�NT�K[5�&4�!����^������N���fs�|���iL�3�<"��}��&^��.�/{�W��)T��=���A��O����t�8^����l�G��,�J�'����3�~ժ]��^8c�x�0f�� K������j��ۭ[Ǆ��Z����BZV�ki�Ysj*�>R)$hժN�	��ؘ(j���-Wy<n@���qY�(�S`19�%Bt��-'»�0~���
o�CQ�"�`�t���R H��dT�o��`�"%BxD��t�W�`pꅲ��O���::�|�շxvܨ�?mc�IG��v���wL[ޮ��&�n�Mj���۴�ɓ'��X!�K!+"�~_O�/`��e��{@=XW�BPLNIo��{@�D܇��g[�z&�]�b�ʢ"�u*��iu�F�]�,6'R��;�{$���yɆ�����^�zv�Bhj��Ѳ�ק��ɟ�/��ꎏW�����S3ߜ:o�Ј+W�k����;���'QW�I� �\!?��I�|�P �`ȯ�B�� ��C��,f(�f��&#����d68��4e��"�>3<�"n`�9.�@�G����ם@ѵ�ݷvo]>���`�o�{~�K?���y�7|��'��Y�x����ٙx�h��W�AWW��xLe|�PMB��K�2��P!V2���t�J8GЛz��X/J%����l�>xV8t1A����8��)��E;*���;�^��}f���%��n�^<��������G:`��}X��ۻ�}���';v\YXX�jl��٩u����פ���pz\,&3��f��O>�����;���]F���61��(br��
���J�<��P�;�Q��v����B<7}�i��5��9;6}����O��	��b���X��Z�=#x�Ծ�=��>Z�׼�7�lM�a���tgr|zC���`2km��f�Y~_4�w �����G~��yM��$�ELB��-�TǾ�w�Sߍ��Ѽu�kJ�`�����!�-�6�rpp��-���P�A��A}p��oU=����Ϝw|����77<�5U�<�R*E��i$C��/�����az˦7|w�֒0E1�,6�,O(Y����USY�8qx��p 7m�k�ǡI��a�ݺ��T<4`�֬ٝ�����P��?��X�Ƶ����f����l&}���(g�͈�9z���Vr� �i#ٸ���^�
����q'�|:�f�.�BV�۷~���|��6�jI�����=T`�b������װa�R�xqa��v���ן)�y
s������v�T>�����x^�Pd�GD6L�>M�<F�kߥ'�q������1������3�sfO��f%���C�߇<6�.�D�G�c��Q[[bt�lF_8<��ɚ�QtxrZ�X��
�Y�cF�Ɓ���4o�{��z�xh���ٶ�?����Z�_�П���C
�K���a�������`�_����?*�I�    IEND�B`�PK
     �8�Z��z� z� /   images/00f35920-432a-4227-a0de-f9ff33566dcd.png�PNG

   IHDR  �     G!��   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^�`Ve����9�Μs��sO�{��Ůc�^Q�		�4�!���;z�QDT{ņE|����{��͗˜��.vw�v�~�j���'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�x�'�xb%??�/DTUU�W�MMM=E9F��؞x�'�x�'�|e�ĉ#������exIaa��O����ǔ���1�L�o���'�x�'�x���E�1����O�(((M����d�\)�9۴�Nu�����95�?��䘯�c����?O<��O<��O�c�����@�N�h�!жQ@�!>���V9��*����-�Eg�N��ͽ�s ����'�x�'�x��w%~��5�ik+D_�4i�{z���2���Je���cя����|!//o�h�L_<a�)��ߙy�'�x�'�x��СC�T ������-��ˢ'���� ����ʱuS�	9�/.��p������S����x�'�x�'�|["@�������r�R�U���2ߔ�� ��>(��T�q��`b�\+ǟ���s��{��x�'�x�'ߦ �eeeW�s�w�\m�d���5e�t�8�=Sun`�S9�]�����d�����?���'�x�'�x�'ߴPW2''��hѢ��^8<���	�N�|ʸS� 0��ߌ:!S�K��w���6����-@f�~���rO<��O<�ēoCp���) X#���O��6�2�Z��>&@,��L�.��NT&�o"yɋ���O<��O<��E��� ))p�H����,�n-,���S�M�u�px�j۰�������A9��2?177�⊊
�ʽ�E�x�'�x�'߄,^��O�%�n ��&PF9��lB�����(��9`���+�rrrʼ�S� �O<��O<������ʺ@�1`Ԏ|S`�˾�e��n�@�����h�:NuBbo�O��� �rn_��!�������ʴ�U�'�x�'�x�MHI���s�@W� �N�π�3L��Km�C�ZHD{[��e2`~"p�377�^��)P�ommm^V�'�x�'�x�ɹ����R ,B�k��+2}�t�i�-�2��e��@�նy�Ԃ&�o����;��d<I�R�����x�'�x�'�|].��Y���������_t�x�'���f��ȭv=�VOm�9�9�7���vj�e�������'E+d��322��9<��O<��O<��B�K����
b���VN��y(++�$p����	�<X��]��0{����Nu�o��=���E������ܻRSS��x�'�x�'�|]��[�~E�rr�ge����(m�N�����\ǧ]�j�q��Ԯmz_="��+p��^�v�`���/ʹO������E6��c~�w�޿~���N�����g�i`�������r��ڧ�x�'�x�MKFF����O�����R swnn�g��@}y̞��u���븧��L�����
V���&����dL�@([�'�Vپ�6��i�m��W_���Ç�m�������=���7����7���K7~}��@������5�^��g�y��̘1�p=�t��?��7`�s�lԶh�ճ�O�m�|O<��O<�v���-�Q �:?�p���g��I�d���sm;����W�Ʌ�T�2;�ʶ�2ߡ2OU��\���B�[i[@�+�O��
����:����ί�������l�#n�Ѿ�������WUU�8Z�o���_q�y?��+�y���{tے��������_�_�?����z���R�}�J�{��^x�<�����@�}�Z�u�,�k��裏�>}��gΜ�o�^�O�~��D��U��[���;_~~�ٳgw�e˖�x�=?�#*���~�c��tۣ��ѝ���7��w�J�uH[���c�������s��O<�ēoG ����rs�+��
v	|�4��!�����}�"��Ӻ��0Q�G����| �������&Ȳ�999�SS�oOHH������?%%�lll�ѣG��5��������W������_q��/��2��~��8���A��

���A�ׯ�k׮�g�}v���v���{d�˪L�:�9��E�}��w�{Dw��⋏`�۲eK�ԩScsss��9r��;n������rK�V���.;�>|���(�ixxx�E�aaa��e�y�= ��*��`��a�������r�=tv��?##�QQi��ⲻ�ʪ��I>��okk��ŋ��1��?}O<��O<�椬yo��L`6���=�sj�m:�*����X���L�4���L29�y'3��?���z*#3{���[RRҚ��[��S5ާ��^.`��2��[n�ᆖ�Do�ׯ���/o���K{�K�C��w�U�����<lȐ��%%K7nذs�޽o���+�>��s��n?z�S�V����gO������g�K/�������7o���Ҳ<~|������v�mͷ�zkz筷�Чw�~{˭7��r�M7��*�0[�[x��-��U�����n֗�#ZBCC[���[F����]w��r������F�7n��;III��O}�$ٖ�.�e�����r�7��U����Ĵ�����>�3f,��E�j~�����O<�ēoF������`����&;'Ϥ�g��ԣ)�iS�ҞKIIݗ���l|B�>������Y��v^rJ��رa����}W]qE�^q�e� {���K.Q�������K�����KNL|}���������7��:d�x���F`=x�`��h�����U���X7P�NԾS��n�i�2���w���[�inj::���aߵW^���]��q��]�o_����w�UW���+�������]}������o�u�]����w��7����	�2dȾ���}�c��ޗ$�Hjr�̉����+���WU]����d_ZZھ�Q���x��.���}�^|��n�u����[����껲]��OK��\NN޳%%e�WWW/oll,mjjon�|Gkk��Z[��������x�'�xrn��4i�\�`���ҭbII�4���>�����O����s޹R۶Sݠ�S`ff昔�	F^ʢ�'��~<1ѧ	�����X}�(�v�jRr��ذ��w�~��+��������_v�*��������2n�?�.8.r���?���p��̧�~j���K��矛cǎ�cǻ����:��i�|w�g繖�ԦS��Ծ�hڽ̭,��/t����2�'�_y���/��"^y��$�_q��e�/��]v��
��\~ǫ���������[�8�8�DGGϘ8�xiI�qi����ӏ/Z����+��{���?��#�W�4�1����\s�����}�z���CCB����݇�{�/�/O:'Ä������yfVα�Iş
�����Z]]��������)��m���-�'�c�O<��OέX�$�|Ҥ�]j~�,��pi��ԗ�����w��;D��g�,0'f*\����0���ZU^�_KSR�M��q�L��o70F��\�MsCQ�u^/z�E鶷�t�IKI1�|Paɓ������ɭ�f�ȑz]�����e�\"���暫�67�p���������A�aC�� YwLH����0q11&Y~�	&��,S$�SeE�ijl4ӦN5sf�6�-2+�/7kV�6k׬1�֮U�9s��HO7��\u��/�}���1c��KN�{G4�}�ML�m�SMڄ�&'7_���LYy�����������ꝵ��'OnK�={�f̘�/�J7y�'�xrn��,Cs�$����I&��'�2��v�9�g�����U'L�B�|̉
����:LJ��p���
�w��	� =��N�9�֖�N�<�w���5W]m�+����b
�����2S&O6s��1˖.5���u�TW�Ze�.Yb�ɲ��v���l�e������5ro�(�������#̝��q�5ט��>�����?�����,�^���j�//�4��5r.զ���ʪ�5�u/�N�2���#d޼y�Z�h���'�x�ɹ�.��$�9� �O�@�q���?`�˥��\������H��a�R��P��2�q�^"�����o4����|�"_}���7n���sն��s�.B;��}Va��������k��2,t�"VH r�c���{μ������T,�;w�4
�X�̴O�j*JK�Ǆ�����䷺Z~s ������W�2����̯~�Z~S�m��[o5c�!`������L�ϋLee����7uu��������7|:��mˌ3�,Xp���뽾�=��O<9���"/�u�ȭ{�awh���U�Ι�-�M��R'`����K�Z�<��i�&������&L0򂏕v�s��^(;�i�:�պQ{L`gb�m��8�����i����r+�mH���t��N��Z���[Ltd����3+W�0m�l�ڳǐPu��!��믛��~�<��j��jY[]mrsrL|L��ѱV_߯�~P�&�_*y������¥��wg�a���h�1{o�E��K���	�&;;��w\SSc�LSS�ihl6M����i��wΙ3�tɒ%׭X��o��O<��O<97r��٥�y]뱝Uێ?�:�0���Թm ����(>>ޤ��j\]ZZ��Rڙ��ar< ����~�D$,D�`LG�5|��y���G}tF�s7�}y�9��g��?6J��GB�@�e~�zD�ٟ��mZ!���|��w4�嘙Gہ�q�ɓ'5��ȑ#�O>�Q��},�N����>܀i]�7\w�>t�I���X�*�*�M��03f���J�,�**��I�eA^����1ٙY&sb�ɔ�=K>,Љ������X7�I�X+��~�K0�q��Na���{f�q�ɱ���P6�ɓ'���V���*��bZZ&�蘱k޼+W��~���`z�'�xrn%`�@fwhs¢�u~꼮���;�ӹ�K- Zv6j�s+�ɋغ��:����#�ǚD���.Q�����%�X��t9�B�$�8`^z�%��+����zKA�u�2ֱzB ���9�N�B��H��Лo����V;,x/���*��KU��q��Q�>�eŶ�< �S9���~ۼ"m<��s�fF��y���0��l�w
��:��<9��^{�S_G���8�v��a� �m��.�睧�	��W]q��w�
�7�p�����Բ��q��w��Ç�@P~W
���֚�i�f��Ef�����G1��|��޽�l߶�l��^�h�"���n���<Gi���� �p�w(��{��އ����^��N��O��lk�&�����̙��\�pq��5�� �O<�ēs.0E�1��L�;ծ��.�]��҄:���i]�Ĭ�b����ڊ��}OHK3ÿA�ư*���Z�q߾}�����O<a^|�E�"@v���W} �a�C �N�i`��8���*�S��t�}�;v�P�
d����zU���d����)�\�1�Ne9��w�^����\�I�pl�'1�{���rCO?��y����g�1/H;���7����m�o��w�/~�3��?��������0�������;s�嗫W6�J}}��?o�@�F�./��^�O�V޷�qN[�l1+W�����R3N�'aK�C�;�4�QQ���׻���˗}����F�Y�f��g���g
lN73�̛7�%��<���O<���%%%���d�`Zh�M-̹���y}�oJ݀	b��ŬMP�6�����쯴�Dݤ�]�%* a� ��<��N�y���� N���d-_��,X�@�#����6��ѭf���j9�H��.+
������H�>��fKSz��C`H�J|���Yh��1�~@�y��u���v'nn��_h����4��B܀	\r��{��]f��O�@, �.|ه�q�sv'�8-��\y�Z/o��fs�@�G�wLt�IIJ�qg�L�b�ΝkV�Xa��^��C��{�l�T�@N���3Ե����7b�0��/��1�cr�m���w���W,�X��˙3g����y��9s�lΑ�#�/ٹb�*?`z1��x�'��c	��%1�������6;m!ιܧv�L;����u�`�.���Ѯ��N�z��=`b�LMIU�䥮�@�l�kWQ^�1y�( ��/���]:Ԃ�s���e�c)Tˣ��.-2��N��5޲E-h:ܶm�Z@����c@VJ�k��'v��@�8޿i�yr�j�.�T�~�4��)�Y�$̰_��8���s<��;:����F��.���X}����0����,`	|;]��J��7������Ir�R�?�Y�|�f���$)W4���4��+d�}�/�Q��L-M�����6�qqj��b:z�5|��g� �^^s�U��-�w�e���A��긟켾�$SZZajk�>�<�%K��ŋ���]��,>�l�ʝ��m(۰a�u�w{��'�x��9������j_f=M��¤]ϧ�y]�8����B�b��9�vK��Ҷ���%]��pa�M�O��s^`-�����dge��$`2N&��G�.X�w�ޫq�O>��Z� F��7��L�n�m���c����:�����J��a�=�����
I,"L,�$᮶��X�L���i���@��pܸ�m��ꪗ�p��rm8g,���st�ȹ����o�:g��r� �֭[�������m@��*I��ITD��V<X��@$�����@�}�b�&܁{@��8C�;I���D��y��2SVVn��jLSS��1c���ʕ��W	0���KWY�z���L>>0=�'�x�'�X �����Y�- :��R�aѭ]˻�/�zN�m�v�[�j�t���y��
�>�x���y1WV��I7�Xuo�^������7���<�S\�V.P�� �{r�;ݾX.��h�j׬Yc�]�^���)���� ��@1����D]Rb�L9M�y�U�^Z��6$�g[��	�X+��0���@�S��b�q����c a_��f[�� �^��	��'1�XDI ��Y�7�p��.p���c��j�� '��1b���������s�;��yTHH0���iB��^!���7�˾����iW|Zj��(/W�(�G�U;�tJax{���L��n�U�֘���x�`֮]��k֬;r�}�v>��Ce۶m� �O<�ēs/N�,((�%�o0�۞��S}�|s�������tu��Շsmm� b�Y(������47����B3j�HL���0�8����=,pE �$� n�KZ��Z�t��6�H�6��\�n�ZDW Q3���:�H��	��cqd;����iw9VJ�����.V�#G}%��V@(� �� H@�6��r�XS�K�q=�1��cr&��vI�:G4����mM�K��llh0mS�hL墅ͪ�+�:���2\�h��5s�.ǲYWSc*��L��gY���<!.Ό;��$��O�9d� u����aR�J���*ۑ���2Yz�Vnذ�<��fs�����_>B��td��v�u+�{�LO<��Oν�����\ �2//o��&�X���?�N�s��F�u1�ۜ�]m;�sn�6zSb�u���ֲ0Ԭ,����5
NV�bccs7{S����S̔��z�A#Gi̝���N�0��N֧�ͥ.�����דXX�(���c>�>�{ "�	<:-�n�Վu\�t�Y�v�!�v��@!�K` �-�'���J`�T ޺��8��$ƀ%�H{m �?��9 ʴ�����[�"Ӹ�7n�h��<��@��m;c0��6�k�\`.4��.�q����,�F�ҘJ����V�Z@� "L�y�Ѵ��W��s�3I?��F垰�L�I1���T�Ƚ�Gʙ�ָ��˹s�իט|H~����*��#:-zD�w��櫯���'�x�'�V,`fggW�����9J���fW?���sz8�j�n�T柾���&%]&��z�))-��skg�@ ��R�ک���י:u�i��kX�@�M&I-�l�XbUd�L�Ҁp�a�sB�S�O +�*�6(`��$+�&0`�z?`��!��@+�F���2j-�}��eNf�|�S@��Wb���	��.��E9G w>��`:%`b��ZS��[n�XJ���U���������lR��@ ���7��g��J��͠����]Mu�&�;����Fu&�����t����d�3ש
�d��ԃ�r��m�O�=�C@�q�͇~��֭��yerm=���O<���K��E.�U����+33�(/T���n��o�c����o���|? vN���T+�4�:��g�m�1�	>�Lfv�����L��>}�io�З�Oyٟ�ӦuW�rڡ�`yY�0a�� y::%�X c��\(1�(@��#q��{L��@@H�r�}��!}o�����'�M�cU�J;�i�	Х�&e� Hzr'���
(��Z�,�% ���!\�$�p�/��3������U$�I�V�8��0s�,��d��by]�~�<�S��S���E\�E�M�|��aA���%4"<\��q���ȱ����=�1}���Dg̘.�Q��:��wߑ)N��n��iv��#��nU�4�t��2�==���O<��܋̔���䴴]���Gs����x Ӫ�xNU�6�(�kNIM3�99������fΜ�Z�������Ky�;ս�̛7�T	���,��g
��� ���db1)�C� \Ƹ�q/�X>{L泼[) i�"� �?����}b%��M,�>����E��(��Q�h�@fO�d��\�v(���ʹs����)������_��3F pΜ9z�XUI�"i�2D�
�:��\WJ@�����׆
8��-@?�m�B%�_������Pd�|�M��4G�i��+���?��H�7o�Bkw��M�Ǭ��!�/[FmN�����xJ�ٳ��I�ګ�;w�:"й󩧞-ۿ���`:�O�299��n���9���<���ߜ'�x�'ߥ�"��ξ!!%�2!1qWrJ�Ѭl_Ws�~��zM���nX�cw(t��l�o�OXRG���u��sLJJ�IJN��7��Mf��fѢ�f�_Q���]:onw]�p�Y�x����3��C4��Bj���vک�ۋ0�.rj_b!���} pEo< �XF$��Sv�,��!@h�������;�8J��
�f�
Q@�*�G,�����k
� +`���k(�.��,�UV���r�XV�X��XS�!���|��_	 RR��o��c�I���M��X�DOooטQ���W�X!�D��S����������d�_��
����
����������`i����,^�� �K�.7K�,��T�.���Fq�3d{��7o&,a���~9��#�8VzL�p���ϗ����~�����*����y999�3�*�=�ls�__ZZ�3Y�����Ӟx�'�|�	�II��qq����gd���s��y�-`ҝ^bb�ILJ1�E�u2qrK�N�������V��K�t����U�BB�Q�Ұo�)��Y �~Ł;\�$��0<��>,�Eٖ�H��l�;�Y	A!B;Z�H�͖%�Q���·�p��j�t��q�l�Y�<�I>�b2T���"�[��0�+$}���:�1R��2����Α�J���RJ����nn��f���?��#�g�����~�[���o���-`�����F�j�j��5k�i�N���k���9o�*ߐ�7mz@~w���
�S�����_��yDt��Ͽ�� ̪������_��!)�,�*�)��d�ծ+ϥ�.,,�F��h���O<�ēo[p�O�8Q3&6v���أ)���(oS���R`��]@��.��N(Z�ۏ��.�� �~��gdd���D� �Y$�3�}��^�n��e��Wu�����ས�e�v3`Z��p�	>V{ N�)`
��"'��� (+@�Zʰ2��Y�CO��X I���'SxR�\b5� �ڳ
��'Ɉ����^�x�f�����n �s�J��D���e�zXd���R��� ��7�<0��N9��-�~� $�5���Z���jkMrb�B�T��pB̟��Kzl�7w��pnĝR_�(�/�Ų�we��0a�c�d�W6�}C)��7_9!�2H-.~�Q���b��+X�_�!
l
h��Η^z���W~��)ϙ���o��2H�Rt��2o����n��u�ɶ�D�d�vi�'�?���O<�ēoS��i3*&fWxT�Ѹ����kJJK��<�;��*�N����}�¡�.0tjw(dh�k���i�
��$�81���ƛ��$9�r3{�<�B����(�8�R0�߿ِ(46,���"{S"2�u0]�iA����Y�t
�p=�xt�VA
��[]�ԟ� �m[���|PA�3I?�������T�t�0����AM���g����
-Y�X�s$�=����XOqa�^�Z�-�8peیt�E��ѧL�U$�� ����o�~H�inj2�uuZz��K@@&+�eԾ�=k�Y,��>m��_�f����_x�>�����{����`ƅ�5�:��)'��C;�i����6(�H����˯��_?hx�s��k���W�|�7�|�;L����MAAA��}����v��=(ϗ�d�}�/�çS�Ce�wd�ei�^�Ε����3�.=��O<��$##��RSS0#Ǐ�v42:Z��0K�>�;\�U�]�>u��5߷n��m�tBawX����]��ަKq��M�`��c0�+���EK��[Ѿ��D��*/xڡ���L��qZ�&��AԂdgy"�t�Z��� ��h�=@Ĳ	�a	$6k�SV��|'Q Ģ�n�m���t
m���_x�E4���l��_tT���	`�X�\!�����m9�ƽN�# �REXV9n�+�~i�*ny��sf���Gr�qs�o8����hoW��x���*۴ʐ�v�H���5UU��EO<d��Qq�wh��+������;���q��d���s��Q�
��R��'�t����7�|�Szۼ��!`�����v�t�[o�w݇~��)?ş�r~#�!�͢��~$������Ϗө|,3<)���|ѱ��g̘�?����O<��ے���� 3%�22*jW���G��&LL7��')d����W� x��H�:]p�0���Lk!%���i۴�wmϐyd�'	�EDF)`VUך�+V�˝r.�����'���2�7w�����02@ïn��VN�nwK��7T�$Xq��I	 �@`I�K�k�{�+p�&�`���6љ䃰O���Ｃ� �%K�_s,�X)���&VB��Էl�X��[k+p
dr�����!�%����y��$�s�0��ړ��2�z�Mf�!&2"�L L$7ה�}C�%%�J���w��}T�=&,LS�79VY�O��*P�h���Zc��{���^t�0)�p�"�k���3t�����3f�SO�tOߔm�\k����1��y��wUg�@��˝2���>���Lq�����A�����<c>��\@�q��ө]��2�^�3�H��p��11��]{�'�x�m	����tC|BBexDĮ#G	Q�/�7�%��a��vAߙ �[{L���K) O�|\|��1�5u�A�ھ}ϩ���(p@;�<��,^�X{|��~���,��uD)�~&��W�H��<@�֭[��	T��C��+X0��s&b�ֺ�m"�m��'���Ll���)@��n���5��82�q�c]�]�q�����y���.w���r�-`bm�����ѣMbBBg�<&2�+��U��
2'3S���[,��ω_&>�~Ʃ�IL&�)��L]�竅3f�x�|�r���Q�sH��o��%np@����(`��\��:��;�{D`s��+���. �	`^.����~y��o��	��T-�J{��n͓�W477��מx�'�|[��<..����1cv6���QAf|L����4E�������i��9�w�2��/�i��Z��FW[=��;ւ��2:&ք��,��f����I����\x9�'_V}�e�yQ�!:2�\y���ik��f���@�K�lG�^O.�Ӊ�>� m@ �a�(�3`����w���-�8���E�{�-�)@%��}���;�d,�d����\�ā�!�¾(���a	%�]�K(Jb�X�E9^�ɹY7�7`�{��{����]#5(��Ι5�4�ՙJ,dr��^z:U敋�3�˗-SK/�yc	ƅ^[]��ϸ�X���;4\���.������S����3kV�1/��ZU_;��9g�l�;���OT?��c���8�Ç�?"�S�S ��o0�y��w�<�D��~Z�<[��LyV�6wʰR�f��w�]{�'�x�m	�~CXXX��]C�=:L^�a�ƙ��d����o�=<7�X{��.��t�kaէ]��*�dH�˴	�&"*ڄ��3�ɩ��u�&I�]{H^���ȩ���]_s��#@p��7T�|�-�n���&&:�\)�}L���6ƱT�n�M]����i:�mڤ��$�P�t�@����E��nH�ٸa��ω�$�3PSHR��I<(0���s�b�: Wƭ8�c�	�\W-�~��79{�lU v�
��Tb�>s�`�2�#�Y�uw:0	|�\CBH����Tkh��=��� ��t �)��!��շ�#��ہ�Pϊ�+��*`~L@�3��'Gt��OI���RJG>�����	`������]�"τzy�<#x0��x��p��6_�����YFmL/��O<���\�c���R92h��a�ͨ��&*f����T@0A�k�흠�]�h1�Y��=��9&9%͌��2!c�
@��)mS�c[����Tw��Ss�}�w��]��� �{����@�m֯�`bǏW��d?`�
��x�i��&��{�$��.I����n"��d�+�-��`�$�Ȗ8ڵ{���I���Ib0��a_C�	m}���z<w��24P&:�L��~��_+�џxKK�B/���J3f���1l�	=Z!jBd��=(8��-"���KX6G����}�������^k�$�G~W~S�|�7���7o��y���>��}��8�m����i�e[ �ώ�u;!��6������uv
p�}�����|���G-�E�z�g��_u�*��_J��n��e�K������O<��ېB�6(4躠ѣ+F�zrȰaGf��aBǆ�Ĕd��G��<���<}V��hw�tZ7�&d
`M�s�7�3MBR�	�0�C�6�M�0O�ة`����?���G.���{V�z|�+�cy�S��}-a�k�0�9��I\�
ﾫ0I�K�`�߷s?X/I��֥�aʶ��q��d|�qN��� �\�)�)���EN9��f�ԩ�Г��b��TS��g��wZ.3&NԾ˱P��������j�"�2釜v�R���P`V+8~c�����.?��H�����ʸ�GV��o;m��lP~��	��_�'N���!�������O?�L�ر3L�tlkk�s�E_522�ϱ".^��/jkk�E`�N��F��E���DL�}��ez��K�����q�r,��xѽ{�v���s��?_������x�'�x���� '`�j��bf�E���&����cZ <}ph�{~�r'T�> [�����ƙhAa����1�i�&.!ٌn�CƘ��	�c:}H���4,>G����Q��^�=�o=yi����
 ��������K���`��|N�}ɞ+!@I� I�O?�D�5g��Lb(�Go6�	nl�aͣ&`JB]-�CO8��q�f��e�}w&���%�w5�р���k<��U�t(� /Z��,%6�.�� j�ҥ�.�2��v@�P�K��Թ�} �}�
��i����Ï���^:v��N��Q�U��mU>�T��DY�g��B��W���I_��4������S��}w�t�(66�_����k	?���4!!�����?����ϊ������\&��)����9q�[H%����>"�)��ʺK��w���Bsrr~���������>o޼�/]�Tu����5k�/f�^��9s��D`�K"�ē�n"�s���9��\�n�_�;bD�ͣ��kF�v��Q#ՊI�u^~���L���� ��H�:�w.?0�C��&���b13�(�LlBR'`�`Θ9G���O�e���_�+�l����_�������*���0mO>$��H#�4���={>I���򾸵���,D'1����]�y�H')�"�X2�O��s!n��ba�:�o8�H� ������-�����5q���qb}�̛���~�z�����h�bb̝�߮�p��������|����0��{K��:��=(�|�K���zir���:G�^�)�l�S��~����W��LOO�}�ĉ!���Q2�xO*ۨ
`�	�����&�����m.((x���䄅C'0���6,����1��˲�����E���
p��N9Vy6�WWW�755�O�2%\`3|��ّ��.[�p��e˖]�~���$_?�����zz�����_�W�?�^��G�Y_K�n�������<$�����������1����Ϙ1�o����f�瞟6rD����#���XS�1�d��Ǜ��LST���>=OQ@�j��m��M7DR����99f���(���hB���Es��y�A~�ڀL^�g�X�؞����?7oy�$��+P��T���L
h�aé@PM��0���@#� `Ԏ���%
(��	"3�}���w���ƛojV:Y��6�I,��'�T8��r�2���t׮�����e����,`��UWi��Mԡ����
UX9R�?��Ƃ��%I<��o�u@�<��R�^�n��:s�����g�!:o�w�����ܾ�q����'��ә��T��)���_w����z��E��[`��
d�%�X P9[��d�J��?���K
����cq?����g�.-`J�F����������d+r��uYO*�u�@�29�e��e���w^6mڴ�g�]>o�����-hЌ�?�m˖�9ٲ�?��'���'��1
�����O�'w�/�WM�>��M��z�s��z��>��H����φ��˛���PW7��-���q7a?�!�GOA����Mm����񪚦��O����=����Y�H{{���/��jj�r��i�.���)��wya���Q��AGC�?�ED�>|x�#�>r�;Æ?���F�1acM��YvV�@[�)-�x)�@P_	����$�.��O��ٓ���<313ӤLH7	)�f||�	;N3M �n"��N�?V�K��^<�emչ�7�7 r��xF��r�?X���Pz��i��7��n��#���T�}X=�هRH��7�P�ߞ��R�&��m۷k�vO}�#��]��:˜������� H68����ڒ�����#���?���K��'ܼu萺�G��Ȳ_Jl@.���:����z�nOI��&�]>R�©���������m�}���ѝ�}L��i�8/��8%%e��!�~�ao*�[}S�9$Ϲ����>����@7,��L�C�O3���2��x���!��@s�
���>$m***:$�š��Ʒ�Mk?4k���OO�>c�ԩ���	˗��q����;�o���O<�#�?��熆�~U5�1�U5�U��э��� ��%(�������8O��͏�a��0��7��J����5���i� �/�q¿�
VCi���&='�����wi�^"���eʔ�+jjb�K�3+kj���:��7o�?�W�y��Oi�?�w�<�%m��De�G�������QR^�^Z^�VUW7H��!��¿�
@)��z��9�OLLx� �|�_�>t��C���jȰ�����#0G��ѣMxd���)�wUU����2���Zqz�����h�h����r��r��ҲRSP�+����n�R�L|r����7!�A�C0�̝k�a�sK���S����a�S�LH���?j��q
l����}.��Xyo��q�! &�))CDQv�/�|���_�~�\R�+���:��/�m�9ݺ,s��-�.'�-���:d��t�ZJ�?����7��:�K��$q��Z�緢}��/�JY��*L\� &����~���e�,`��{R+�i��y��)�}L���<W.�g�܆ɛ�=)Ϭ��U�:����=���� �z|��{�� ٓ:�Ҫu����%�WM��X��<����I9֓999'�xOVUU����IyG|�����ԩ�ސ���;:f���`Q��'��/_~ي+���'�|�"�������!����!%��hizF֖��IK�S��ڮnmm�,��r���Y��pqqq�������������7��7�D�jɌlk����_���QZ^՜�����̬M�B�3f��`����XW��AsU�O����2.""<>>)63'g�<�ίho����� �6m�e5����y�Kʶ/n�֑�`��+g̨�|�_����^7>nxTLL\rjj� �����w������<y�i�95}��&N�TRVQ���>����?��וc�Ӳ���ML�5":"<66>V^�sr��wv�V������b��'�	[%���#�>�6̸79u1���J���h�L]}�_�k��C;���;��?C��E�ê�j3���d��y�$����$?`�	3���9W +�� fo�L@&ɋ�ʴU��) r�Wh<�m'��r��hHn�y)II=�`~Sr�k�^n�q��Rǵ(^�u8��n�@��&�[n���.r-�~���EdmM�ٶm����.3��C{a>��:����
_�h�"����H����߫v�ȶ�a!�Z}6�)G~�r�
t�d�|B�DƯ�Y����\+**�P�'07�~�uP>��J�XS�e{����0}��L'���}���O@eڪ��i�� ay.���<=^�������9k��h��J �i�:M�2�)�y�ӧ�̟?��ݻ7{��'�w��������kl>��tZRJ�K�c�L��z���aq�ԩ)������wrSӔ�&���ff�LNO�\9qb�����²��;k����"k[;����iDeM]}fv���c�?�OH��������ӫ;:fino��c�=��e���D\�##���C��Ư���k))/��il<�j���7�?��u-mL*�KL~9z|쑬��W�ZZ͘1+iڴi���e��Y�ddeō�&к2)%e^vn~Aii���dRZ����ʲ��	�["��>�������d��i�-S��ni�?���e�~RX\xϸ��������11+22���X"jjj�L��G��	II�c�,=��Q��'�g��f��!� sd�(2�DFG���\��mSL��V���PY�^n���ݹP�~�@00�+P�"/�����l�b��h��*/�o0��K/��\%�Bv11W_y���/̿�k�\���#��o��q��cJP��-̳��r�c���9�C�uγ㈝FYO�9�=��tlv[+vu��2籹��N����ƒ��0&$T���{7ܫ	;���G׹V@��C$��⧤���D"�}7jL,������$�bP��� �܊\���O�)`uANN���Lx@��_gm��"�@��t���;ݥN��=&.r �}�9V���Q^�2����^XX 험��jL�J3s�l���o�̙g�;f|����Y]}���M����c.\x)�z�e��O��BLaUU���
&Ŧ�MX�Q��y dY]S�RS��ō��	�7�5M����.*5m�ܨ��O��'8{���tSYMCQuSk��涫&w+������y,6.����h���BI�[Z�/�j��mW�Ϝyw~aaiظq�

: ����}J sVecݘ�����ZY�xU^Aф�ԍ�""?���!�������mSN�6=��}��s�,���u���	��G�<;f��C�II���l*��*��������g���,//6ab�9�BƌѾ���߯oj���:��i��{��|[ffg���	}H������C�Y{F�WTT�����V��M��iIɩ+��W�G�����G�!C���C,`��H6��'&���b���lڦMU�l�2Y����)�3O���(���|]�.��_�7�؀��IE&m� fr��IH2�1�&8t� �����@��6	��
�X%�dB>(�=Z��9|��R��辮_?���i��}8����L1755+)�3���u(�����lK���c9�n�	��s�h��m�b��Ͷ����q��[X��H�a�@����5���0�<C�z�������Vk^gy�M7����7񱱦��QAr�E:�;g�f�7��+���7��
�X.e,;�y����-�gr�v��S+��6�uڮ�����?��� Y�k�����EN�,l��0KOL��ww-+�=��J����w�*��(h�e}}�im�l::���?�,^��,]��,\�X˞	d����'�9��eJ��9/�ϒ�'�W��XYY^bJzJxD�}�CB? .0'7�TV�|����\��ŭmm�����Y9�sǅG==|�ȣ�&-}��F��pcucK]m��I�MS���>:>.�p���CǄ	H%�M2���Nn�2}ƌֶi�&�WU5&���4:�M\ƚ���w���⩊ں��������e�u�SR'L	;v����G�#"MFV�)-�<��<yߴ��䫷l���Ҳ���11q�1�XhX�IL�}�Q^Q�AP�����qe���EDF��s94rԨ� f~�$S]���斶�榖ɓJJʚ�9j�[$���ƙ���O'��直��YQS[,�V�����syQ��� �QA��#OL��36<ܤ˃���J��S��)�a-dx:m���n�f>��c��:v�U�:=)��1�%e�&=3C���(	0��y�|x��ӻ��k���$$K^x�'�85)S�2Na�������[n��>@�x@�i��!�$� _n8�XF������� VIb�:�������@�[��c�d=f�w�}Q���{96`h�i���0�� Ӈ�=������L�l����L���tܺ�{����H�b�X�|�Y���H�cRa�*������
Dx�Z��`J�
����\�%����}1N~�_����2��N�zAUUU� ����r����@V@���nݡ�w�D�ʨu�Z��	�Z�%��iI�O��X-�q�uu����U��s��5�-1˗�4+W�2+D	l��u���=[RR>[>�c2/]�x���忤�x���E8�Ú����&���I ��q�&+'�T����Z���2y���*��KL|A���AL��&ff��Ҋ��uoU׷<Q]��peu�әY9���A f�<��ON�2�3��i�:mKN^ޓcƎ}g��!'�F	�$�<y`�VT~ZQS����~UmCS{qE��������:l؉q������)G�Ϙ���9s���7m��>���!c��5#��$�M*9!�y������چ9r���3ׄ��>?pР�F����7��0�lln}oʴ�ݍ--[���w�;�{��v�����'�]�qYU�seU��TV�n�T\�zBR����f8V�QA
���3\/�":7�H����= N�ϯ-SZU;�]@h]�v�o���\ֹܶa�i[�y����j�����6�>q�g��h9����ͨ�P32H 3�۱`�^���<bƏ�J��ax	��KP^>Z')!A-���v��0�� ��G�u��g� 8��7�X����t����b��tl�O!w��t`žX�d}k�t
�p\X^{j�u���u%���z!�	@�Z���X1�X���lCf8�豇�iӴ���5k�C>�1�e�M��;1����e��\ ��t�s��7����W�5�!״N�}�O<�_�R�ܞ"�?�7o�Myp[�>�H�s�]oj��֦E'M*R��@��):�j(�j��}pL�G�X.��>2�IYH�MMM����'p9mZ��=���k֮7��mP]�j�Z2[Z�ȹ�����_ZZ1��eJtKK˥555￤�x���Epє�T�����1($��X̉�%\	`�N6�-'����-(x/,|���1���I��2��UF ��Ə�*k�-(�t�`�ѣG�A���8.1�������6����iMm����ɟ`ѻ{��fĨ&6!����pyuz����`qYž���ã��<lȗC�5�fBF�0���Sۿ�<e�a��Q��?:t��g�3:$̤���M6t�W�U��W0�ل���F�u�s�4ѱ�&����4�l#/��ɟVTV�+����Qr��V���Y//�)��>^R^�����/����0H,�#F��0����R��5���w�)�����A�ȉ�'��m&.rb��5ccb46�7��%�TW� &��qaa���R0����,r����f�Se(c�14�˂F r��)�і�=�Y�8ܠ��ql���F��wΓv�F�tl������1���=���,�m2�	0��0��Ɔuy��uu��� '��6��fϜ���X�ɖ�:S��ދ�H�w�5����N���'�D����Ç?,�5O?���Gy�?	E�ׯ�(~�n޼��֯_��۷o��U��ko��VWW���ґZ��\�Ve~�j�WT��%Ѻ��0���X/��߳A~7���@�r�=�(���,�o9�K�[�\��^sߦ̦��!��|�
] ����Yvv�3E�%��|�4e�E���+�w��'����0!!����1��	`�(`fd�`��y���/̢�ү��R�=&��g�0�	`f���ZY��TTכ�����'���(3B^6 ��`'/�"���&7����Z��'#� ���%@��yHV�C���(�23'�XBr���А���VPÂ���e�*�[LM]��Z�W���3f�$p9����/�:S&0��W�yJ�c��Æ�s!.2:N��h����o4eU&3;�dDT�2bh'`� �y��ڔ	�N*�*#3�$`!����s��.&�>�+m�]dRR������?�a�t]���.���\תo��m���Z���=o�}�VٷB��̤��2A~kQF>N:]�s��1����'��/��)��u��LC�C�8>�b"I2ĒI_���c�kb���y�&0�L�y�9���K������5��%���+��e|���u�;�fO���:�MQq�{��CJ�ܺ�g�p��S��6��r��ǐ�X�С7�m��������9�{iKq|/�8u5<h>��C�-��U$.k~#��<�		Q����<P��(��ʇB� )��C�Q��8"p��Ν�]N� ��)�P׸.��<5��y-�[����jł�\�r��ݻ��ݻwW�{ｃ�Ηg�˽�oh�*0��ٳg�n�ڵ��gϞ�Pk���Z[[O��^����������\�E
�n�T`��ɞ�v���D�@N�<�L�Ҧ��S�X��ʺ]J���1NBϼ�o�f�:s�}���=l~d��C2μ5��j�O�<�� %���0q�%e�[�L%��gr\^1vO<��Ȑ!C~2n�ya��%����3��	�5���f�t&[(����
��`5+ ��#�Wk�jM� \^^�ILL2��:t���0�L��[�@YA�$�t�7N�x1r�!�P��˫�M)����r|L�@Y�/{� ��Db0+��v�sL\l�	1�\���I��T,��jy�V��)_�i�}>dذN�/�`����9����j���z�O�q���&V���,.�4��E��'&�0)K�`:v�� /К�Zr��=w]�gA�L߾N�8���J�m�+��1���`Ǘ���zX-������ɺX7#��d�u���{L�����yR������ 7o�"}?�u��!�`�<f w:�裏jMG����q ȴ�	�h���}�"�plX�v�:엌���G��K;zl�?z��*��5�ylLG�Ԟ=�;t{�KM�z؞n(m?�vg��]�6��	�aE���X4����:�?�wSE��by)b8���?�TD=ͼ��N����L~k�0�ZQ�s�ʕ�
 ?"؜���������2433sH^^^��[�,��6�����g���1�$�5c�#�f����351�U\�t���_`���	��0�؆�F��Y3�p֬�tv@e�����rŊ�fÆ����{�ީv�����q>��q�L�/\�D���I�w���inn�#�����q�k�%�x���E �~�6ncph��q��yj��mlV+]��A���{8�0Yٹj���i0��%&Y�,��*�
�LLN��j2�~aQ� V�Ǣ7��d�4!K'��
K�vI��0
��XY�`� ��� ����[,�@0��i&�)�J�
�_P��es������|�f��"��Ҋj8�O�� (ǈ?.!��� ���$i��D@+:ڌ�s�k�	��:S`��$3a���ֺ�
��rp��-ȩ���cܵ�U�]�|p���e��NXu�w��W���7yFv��0�ZR�hdP�|8���} L�ڊs�{9��-��(���H�.T��X/L�v��������q\�7:�Y��(�M�@�~±�a����$�0d1��t�4,�NW3F�@o�  JB���o϶	PZ�D��[�)��[`kÆ�E2���ѡ_�4ҋΊ�+��۷���۱�ې��q�?8��& I����D{'�J�(��i+�,�r]L[��>)}�k�R?D�떲��~RG�b�0�j�#�+'�;�;c0;]�?����=��~tO�r�-	S@95;�N��澟���;55uMrr�\̙2>#--m��_)��DII�;�����?�Y�d��.X�H�����EK�Μ5G�m�!7/O{ܢw0�ye��wN�,Q�I�hb��x���Űo��S�-[!�Z��X(�ly�l߾��ڵG�!�W>~�f�.����l��6mS��8���>6.�����rs����kF,X����_m�x��w-]�?`����̚�&uUc!L�?h�.�K�#ۼ��F��T\n��"�#�,`&%����V ���V��N�g,���@�$p:I��,ț$�܂B��1c��,`b�$���Δ��c�UT�;H�1T@7}b��~�K{��3�L��9�Q� 3_�U���YE���1�1b}���u 0��xu��,�
�#O�!r�Կ�J�467���?����^~�\CrԷ	��&nnj]�����.��^"qX9K��9¹99�v�*��m�rv�)L�1���>0�G@��G�!���{�l@Ú�r7`b%
�7�{�-۞-=���8�v�Jh�#Ǵe�m@��؞�UڤKI ���P+�G����Ժ*��Fg�?.q,�XP����-O� �v�C �yVzL'��nt�W+�c>���A�a��R���#pi��T�v�`2��|$�M'������Xb����U̗QƓ��ސ�'�3�j&k��C�īW��]�A���b���:�j�-�������L�1�Bj��}tMz��bO�K��i���3�6=`6o�"K���򩧞�{�9��_0ϋ�{/�3��!Е��PS×x�ȳ�������%ޟ���-�y%Y��5<�ē�H L���	`�	`�`�GF���|��\�{�Zk����q�]�"�	db�T��V��ܱ�aq
	1I)i��[)��h*d]�$����X&V�O8a_X/'�W*`��M9���A�d<K�S!�[��zE�%&#S�1*���U>��p�R��R�L�s���R�F�i76�+�6�*����r��7p� �����'Л_$[Y�P���p���>|�B����&�`ʩ��zUt�'��P��~u�w��ʞ�}z��T=l��E�d��6��y�%����2#�C���7�`Zq���{>�L �*C`���$�fY���'�r	lPO��]�e�"�N��I>�Cc�4�P��`�Lw�?�4�B �3@PH<#��nW�m��ys�����Th
���^}U]���	x/
���?�˱���\[��J
|r�
�@���'�R�h��y9��<�mc�u��L����Np�[�D����-�-�iն��(����ma�����}���U���;�e6J(�@��wͽ7��/^�'�e�Î@嗢'�����	�/���}���7�l�h�	�͚=ה���yXJ���p�w����@�L�ɗD��E�.\�ǻu�c桇�Evh���~T�ݮ�{�S��O��!~U����+2|ᅗ�~�o�|r��c���>s��Y���h�ED}1n\���ccg����������U�+�O<��$ `FE����SYW/�X%0T�Ev ���� �b���*y�U�¢I�)j��Y�B:&�ŭ�Y._�|U��6v���`�����= �H���by��F+i3'_ ��Nן$_����x��)��������J��Qb@��1���	pb�0�.�ڙ�:A�#둰$���	`��W�!^s� L�?�	�>b� &1���}�9T�S�=/W�^ĺ��
��a�KX��/�9�[�S
��u��:V�p��ơaaZ�� \�Z�5�8�0�,�B�0�'�pX���M����M~����ބk�;�m�C�&I��-�ܜ�A�`��1��&�[�|Q@�3S�� ��	犕�ZO9zӡf'Ǌ������zO��ke�'��讓i�*Q =﷿�T��2�:VI���m~�_��ɐimï��q������o
0O�l��_���	�����l��h{�Aݽ�dd���S�R>4,Xh}t����=�����4;w��q��z� %���CX)��s�X/�a ����+W龱:2�I��@ʹ�- 	X��!D�T|S��^�e{�<m�>���)���!>)��wȸ��c��gOvqq���:��y�'ߕt���sX�`�ih2� ��XY]k�����Hމ���+,�
d�a(�#������PYwth�� �*���f�^��$��j<"Ј�8]�����eg�i��d,c)ÂH�"��T- �P;��v��D��^d��)n#`�Y3��8���O,&��j�h�2����t�e���<I�`f�
dOR�)qO�q��8LY���p�KJ&"�)�#�П7�X��>���AcO�y6j]�X_I��(בD�A�f�(����{ �&��E���)V��d��x
���8�	���.u�c�(I@ �@���D,X��@ZUk�@��/\� �bzڦ =*ۢ��|����v�=6��c �P�<�<���: 2�����u�q�?�k�ٴi�ٸq�vӈk�9�V@�f�4�s#m�f�D�VH��V�]��C���t��u&����&���9�1�Q��4���	�E���+����Z[�h��"Q����k�i`�\���k��������������l���Y���d2�YZV.�X��.��>�K�`�;�!e�p�sܔڰ�^�7G�=)�إL��a�|�W"��C�ޖ���W}��4_�u�y�Y���'̽7�9s盚���w))Es\D�ф���ӳ�Jگx?m7��x��7,� 3r|�[}� Y�� ��/F@/99Mc&(���ZE���q�U2�_P��ln &���&S�@�|A`VK۔$/�E\%�Q���HeU�L�$����6�&jF����I�N��čΐ�HJԄ���S�"��W<p��_�;fi/OP��-`&&��
۪Z�-���`�Rw:Eщ���e �@�73���J�XY��1)��0���q��n5Q��=��.�$6�aA�	 5��cyJ��[���&�{[Ƿ&��>I�ɑq�
�#{L��tӁ�	����h�ذ0�yIQu�,I
a7:�NP��S����oW8q�u���9�����\�(b�ú�no1@-�:�9a1$��=B�7��@�S(�����¶�q\�@"�N�p���={	A$� �$�l�i�K���uϹr�n�6���u�����徏�������FU>��@8�!d��@�?��F�e�M��7�jMoA|p�O�� �Lα/��o���	��/N|e>��?�K�ӯ�{�h�m{�L�>Ӕ�3(�rA򁌋�j�<_���,�i��r�))��|<�!����_?xZ=pP֗!ж���������Y�<�0}]=���i�N*��c 3u,q�cq|��wuس�٩��@%%���$v���O�#��2_�� @?�s��oӃf���t�ar	ϑg���h<(G�R�vfd�O�����'�|$`���˙"�<��P�@_��W��L<:Da�z��V��"n�"u744+�������cv�in�b��'���o8����q�gX/K`��Ģ|8-mTנ�:Fc@�byh6��*X�@cUU���2vl�>b��m��ب7	`���U�V��K�;�y��ɩi����+(R����`;��� &��r���
盜|X9�|L���<�J����)�4�A��H�_N��.`V��?��0�5�i��Ouڂc��v��֧֭�n#��6�m\�ve�zyѐ�J,�0G�0�j%�2�)��u�[+�������(�� F���(�=��E{��������Z!����!V:\�mެ.a`
e>�F�0 F�$�q�8��@��5!K��qi�pAio�R&�,s���˗_y�<&@HV;Y�Q�	H$��L����@3��>�.�:� �|��(VL���2����緹��;M��"��iI=���=E��t��l�2�x�b�<�z�:g���z�*��|�I\-nt~[�"�	0ݿKob�e��'�˓�P��O�c_�5�D�|r�f�SƧZ��<�(T+�V���<֙={��Ǳ�}������ޡX�N����e��Y(�BJ��ɡK��r����쏜i��y�N���Z�|ؓ���d�qwW{�]��s�a9�>��|�
(䏗�s���D��ӄ�|�VL������f>׶����&�3�^�0�$$�<���U6f���x�3Ӗ)�?ޔ�Wk��)>�Ы�kljQk}��DC�#P���NmH_�𩦾�Q�0�$��@��h�<��d�� =�a٣�{v^�c�jIF7���i
z<8�q���Ni�c��#�n�
Ldd�n0'˲jݞ�0��[M�<�#���~c��g-_��
��5=��>'�s��Βmk�$y`ge��yWʋ�^�#�>T �8p������d��> �����w ��\0h!�������}`���mh�������蚶�;U��&��y��@�=! �s���b�z�w�[�L�zn��f�(��e�O4'��4y�`�2��I��ʰ1c�����j��y�M&ڳ{��$�$�Pnh���1`W5�@�E �yԁ�80�0�5r��V+� J[*��"v�.�B��{S���gY �'�;�9�' �&K�5��I�)�L�p�l[� ���CW��C^&�ŵ'S\����@
�_"P	��\O��d}��t+�����D��\�9�gk.�p�1X�tZ[����o��[V����/�gǾ0GE?;~�|��	��/���O=�W����ak��=��j��S[d>�ɧN�f�,Yjv�|R!���c2����U����|j>=�������c�}��8>f�)(,����⻔i�P���LO*�g]�IM��)�;k��;�0<*��	~��[9.�k�'V(?��0_oSǏ.�|,�T�g�y������;�1��yr�-UDI&�E���Mr�1>�D�$)%m��e��g��ē�^܀I�u����\K�'	�d "�Gz�!S�,I\� 1�Y9yjE�1s�����72h�		V7j����I�:��)<��
��D`���(/u��W}�<�gΙ� I,$u8ǆ�k�m�Oڨ��ShU�i\��kZ�Ċ�y���G��K�k\�i�L�<8�hs L�Fy9�[\!8T 87���թ4++W��@A�6�W
��K��ry׀���ib����Xd�{�S@�? Z0�a����hU�9������O�ׇsd�l �Jo˝��1���tZb0�*�'
�0�yJ����X8���a�����X�w�}W��X�4��;�(�hY�ȑ ��Z-{�J�B����)\�_����l˾S��cC��n߾]A����iƹ?y�	�=	�b�����.1�6��0�����b�$W���)��X�I�B	q�(+S��}J&�e�ˇ,��`&����C�D.�5.bJQH��	̋/>'��u����W���/̑�����g�>7`CI]G���f�ўj�c۩�G��[��{ȠO`��|z�We]�[~Jgm�����<}��K��5�՚�S+�T��5�ZK�c�:���vu�[����G|�&8���k�nٷ��@�q�m��K��n*�m�]�3������3��Q���ʫf�&�J�E��d�?�(�9!3�LO<���鬃9*8�0�+�*56��J2�'O���|q{I�6�	hd &�ωa���$����b��Hn~�l�O@(��Y���B�1B3�s0I��[E0��;���+�y��Bb7Nc=�Y��$�Pj�aI����%�`偄��<��3�|&ff�!C�i���ֶ6� ���,��2�M���=F ���A�M� f�� �+/�!"2Z�җ�3`�=殻�ȼ[3ГSS�9G��� ����s�.��`�i��m캝j�隶��	��m;���a�Ǐ�?=c�		�/�Qz�}���I�/��2rZ����jH�(�A� ��#@
���Db�|b�tZ�%m��\Ȧ�j��K0I'� �W�M�M��NP$�Z8����zlX��H����*�~8F�$@"��*�:�Z7��r�̳�LgO>\c�ր�u��iY(U�ke�4E�)����V� ']z�h��1/�X����M��]��I�L�`: ��	$�zZ��nu�	P~���:��G�'�ҟ�g7H��c���+V
�3��uӎSǒ�=l0�;�}Q���+�~'5Yl�|d�!<l����,�.4˗S؜B�KE}��q�����e�U�Y�j�Y�x�<�k��1E!���c��Ór]P��N��-�s�w���5d�����w~MK�����n��<��_$���:�#!%�4u��k���=��ē�Zz̪�j3���0C����̨� }������F�����5k�*ԥ`�P3{�<is��.\�D{f��oԢ�X1�7`�����6n2�g�21����>���ZKVhy�~�����5C<dL�0KK�y aq�(�X���L����䜛��I�"�M�O�a�2}�YoJ�%H�L9���mf��0��FEǘ����B�X-`b�� 2�q���
˵�FI(��$`:�`�K̕W\a�� `�H&X-�Lܳ�Z��сS����Vؿ�o_�n	4�),w��l�*�'�!׍m�m��8���¶@�-�d3řFwN�XG��R ނ����R���ʸ�"�2F@?nn�J	5�;w��N��|P�~�@Sp�$�t���Y���߻\��0O�#G�	L~�Cb�ĥM� �7��!F��H��ۚ����%pIY��ߐ߼+7�qR�����M���Y>�I�Y�x�ٱc�^S��g���Y�wo ��M�]�{�9���'ͬ9��y'?r�'��?a$���c�i�{�U��\SJ�����D�ę1�"���G�� �O�/��__�c�6�
R����>}��ҵ"�A 
@��E}pCw &�l
�WWי�6ꃠ��ބ��QK"qA��/�vf���Ij	]�l�~��Z�r 33'�4�W7���&'�Ys癇~��_�H�K6w�� �Y����ju}�6Y <k�\�_X ��fY��f�����D$z�X�v���RBC�(�M�sn��f���0g�Γ������I`��ť�&5-]!�s ��*<` py��� L\�v[��\l�~���;��gc2�:����9��iW�_�������`����d wAQ��#�������\�nuK���I6�W]�K�,ZO�Ri{�,�44H�!��ڃ�^I>�8;ֳ� �
u\΅uz+�sB���� �E�C�g�qcӃ
�Yȴb�s�E�f�tO�ܞsa����v��t,� 1�$���ۚ� �Baw��M����l	!`��;n�����.�V��.Ԥ"��֯�8L�������L�1��KNv<��o�����I]�޲��u�j��i�|��!|���\�.eudb�桷5f�n�O���O�Ъ�s�p��ݚ!��;��b�N=U�?�L��I����Ԣ����V(��V��9�rOq�����f��U�f|B�<Z{�ގ�.s_S�u�R��/�*L)# s����hni�%J�E�� 3tܸ���`z���E� 3L s� ��$�� sF'`vL�)@�^k�Q��ln�y$�� L�c'n�8��$��c�����:�{@���@R[�3�W�����s�/4��!�|�*C�v��Ʈ��V�{� #�簾V�t�r�x�R9�23V�͹PC�fFf�&`KF"�
Q��E>U �I 337Os���u�S�H�!$��C�'ׇ��ȣ��e�n�@lHh�9*X��@L7�c�Ǚ��|��`RϳD ��/CB��L\��ωx����|}����JzLINN�%���D���4_y�\��M$�M�!�3���)쓗-���K���HY:�?Jad\����:����t����E۞SXαq\�t���<��c�� �-�7�%K�tB�h�Z6�K����֭S� VL+=&=� }���g�~�Q\���ot�z�-腫U>0��>(��|�23s�L3���L��R�j�*�7D׭]�I,�Ce�Q~���%��j�|���̡��1o������l��.���2�DckZ2�JmH;|�����ԁ �}V��`*`�����l��;������&+'������@ ��g�KO���w���`v��N�ǂ�#<&�415�LO<�>�0G�	�8b���dhO$����4��%K��"y��͍E�8Dj�iw�3��і����3��C��G)`��`�>s���5k�	�n�6�kB���њ B�Om]�f^a���h�yr�S�(���N2ر�����1�M����jy���ךq�X�|I9��yߦqϏ
k�ϔ�v-ϔ!`��5\��qs��C�ty�M�ڮ�X/�ٻ_�$�x���0!�;H��ݢ�I
i���|��B7,������}�Z���R;߽^�m���.��R�v�&ע��J]� x��̞�#����LLt�杷ݦu��Hy*j`�. K\��U�jIb�&w�q�Z/!g�OO��|`�#��s�Wo� ����)#Cm�����8J�7qm�&��ɺ�{j(�m�H��'��)�m���6I5$/��a��\��xK���U��Pjdb�d��n�)஀)׷`
D���J,�k)��P��~/>r�7ͧ �|���s�B�7Ԏ�tVi{�
@�N�u��u�>8p�c�<H�3�oP2h~�Y��yW��x��#�v�N����dS�<��[[q��v�G���?�]���Z���ه}� &�b'`ʇ$.r��ގͩVz�v�G�$l ��EN9�m\�|��n�`@ޱ��"]�%�x���A܀)��@�0��X@Ԫի�*4��3%jp�S0=M�
W�[���f���w;�If��ՂI	 ��֮[ov<�Ӭ^��P��*Eȁ�ZBL��������+_���t��!~�Ă9Gp$�g����ª!p���v��	�XY�?�C��q������SMCs�Ɠ�E>O��ލ�����װ�R3��|P�*���{^�!~����c۶k�y�;�U ft�x��Y˟��X�c d pظ�_ۂ��|�	��\y����5#�9@����\b�LN�X���u�S�>�m�u,^}L��@,��A�SN
�b *�\� q�,���=��Y�$��:�j-�=] �(�>tI���pnh�C���q�ۂ�ւ��1�w��ՁX,�N�u[05�\@���wݥ��� �Ç��	9��GrY�t�ɼĸ8�X($᮰P��|,kIr��%^�VK\���j=�}��y\�W������9���7���F��;�?��#G>3�x�P���CN�UM�b����q�i�|�0�}L`p����@�������æ��>r�r_��/Y���"OJ4��o��̗0���Q���fXdd����k###=��ē�Z0CB�	K�QL�q�VVW+Te$�Li�&��Q�p�&׌��EDT�)���`����2I����=g�ϟo���ďH���>S�9��p,�;��e�oؠN 3>1A����� 37���_��<#������y�>�q�s��`��z�r�j��`dT��ǃ�u9�c} �qyYҋ}�:�P�qJ�T��$��l��r���ŋN3��89ƹ�����Q�TL
O=����I��� ��� o�6UP󹝭v��.H�_'�Y�󯯐�Zǽmg��eNp��u�ծmfi�s����V����F�)�y�@�&����s}L����{���	 �
ns@�X>,��iL�|��dg�� �=h�0���O���1���>����H����{~�|G��n�pus� 7`��k`�.��Ⱦf�@1��k�s9�O�K�����s�N'C�k�$�p\'��?'`zZS �Z��x�"C���y�zU����J���׫Քh
���58-��q���
�2��"� l�����5��b��cu,_y�u�W_;`^�i��K���Wˑ��7�<ϩ
D�i���18�q�����q��%���3o�<��g�V��~�>�����o�f���i��b�<	�I�a��3�]�Vb�ZfŹJ\)��/�����ē�I{�0�` `�$Y�c#�v\z��'��̐�Q��7ʃI s����ָK���olim�Wa��[p�����[]G��"4b2)F�5eᢅ&V@ ����QX�M2���+4��x�}�B� &u"q�[������?X07X��C㸪�E>k�~ɒxDf:�H��
�EEGi{FV���㲀�W��%�.Y��w�M��%�&fd
�j64h�u��!/��1��@��{�A�:m�f����:[QU��0�N1�-���g"䚧��}c�	��2E�ELJa�L��% ���n��#Aݫ�E�?9�(�@W	`��`�$���:�e|l o nv��������e�.-�b1�#Ŷ�S������˞������?J�������!�
d��w��{L�<j`R��^��qg�9f�f���fzG��ho�T�I��C�jj�b�|�OJQ�q@)"��<Ӿ���Ya��ώ���~G�j��K/���/�jo<|$��	]�W��V �jݕyvߧ;��ֳ�I�%�>h�����p�*�g��̗��E��.>�D0�~;�����^|�<�c�z�<��ē?0G��8/8$8yd�Z��ƅ���j�1,)+W7ЅK[���"!c��7V�֘���T��G}Ts�����f�Bٌ��Lv^���)Q���'��WK(���~��Н�2L�
��g�C�D��f�F�ɧC^Vťe5���l�
MD��n�c�e�`���.�[)�k�4��%���
��u)�`R�I^�|	�Μ=Ks�ʕj�0q�ϑ.@Л��ƛ
����#�O�'��"���8�vB����;����ƻo�[�.g;���n����:�`6On1y�t��*���}��ȭ8_(�en0m�u�xOI�n�d�]���Qۓ�苜 �m(m`��"?�q X&�>�n��ڴ}}n�l_z�E��4I*��ޢKG J�ht���m���=�J�9.x�/P�t>@,�b@$�&�`8Q����Y�B�m���EN_��	d�@(�I��/�L��x��QQ��E�8�>�ȵ�W�X�Y��%��<W�H���z�Z*_|���/�������~��jq�"v{g�y��V-�i]��=�f����j<{k�d�����Nm���m0S�96���<#�锞�1�|;ϭNa����ͻ�6�=��ٶ}����	�L�q ����h0=���"]�9*y䨑|���ʚ�Nx#YW��5k�}�6�U�x±��h��X0I�!S{��� ̥˖����N�\�p�f}���h�L\�@%�I���Ղ)�3IbЮ=O�-�<� J��uR&hZ�t&��ɲr�d�2�Ж�d?3����39a���0�tMRk,�i�
� &���Q`��2�5�R s͚5�/�!�Bf�k���~��y˵-/N�cbf�>��;&��#�ǵ�6 �8<z�0���k!uQ�����E:%y�%�^}�U#x��ן��q��@���E��>|X�%F��]�R�vOs�X����K�����6����>����b� �'d}Ɲ�H�[�8�'�G6i��8��}]i�&�`��T��M
��r��@(I���m۴�",�V��Iv>�gc")z~���+��׿���u-Q,�(�o���.����u z��8Vh\䴁[��L
�s]|C��E���pQƟ�E��枱�i�l����=H,`�L惖�{�7ͭ��H2�3U�֩|`�"'���E�1�|;ϭNa��c�5qj����c��0ã���GG�� �O�/��9b�y��G%�9b����2�u�ء�>j=[�kV��q1Z���e�r
��͞)λ|�r�"_����.X$�)����or�
���5ɇR$a���NW���C�9G r��
��e���8�J�!̒R���"�[l-^��;g��륦����
��r.����R��d��� d
�746�E+&����hWt��܎g:�w�U�70�R�O��-�>K���NU���N�������@�@3��N�t�m7��,/�0��Df�����y&`�2EԾ��%�!��(����� 0(�)�m�dR��!I�ٓ�=V`���4�V}�e��������M/4����)`��X'%�q��'�(�}��-K��>@J� g����x\ �ޅۺU��$@�c�� #0���A��m�R�(��2ڳ��s�� �� �D)���s���8P�~�b�e�%J�,�L~# �$�ٳg�M��׉��1��Ͼ����r��н�q\�$��������3ϊ2N��˯�j>3��+�e�	��C�+�J<sI��ol��S��9����e�K��߹̹\Ʊb��~#�����|�{Yo�Z�ZL8�S{�ݯ��(/7W �I ��Čl��̨�Q�cK��⮉���=�� ����1jD��0�Ц�� #�A�K�-��l����ǚ1����U��t����M��w���1�xqSgdfʗ�|�Ff�䙬�|3w�|} L^YU��9.2\����&�0���.�YQQnF�:0����� �y��	`�i�MrZ�)���yp$+~��uf�9s�f�+`&'`�i�@�3.s�c0�>M*���9v�X����G�l�D#�x�S�\S�������F�u_G��T�����=��k~�ud�n��mv-��ڗ�s�o;�<��OH�������&�� (X3Mk���u%	��LQ���Ml�$�L,�6��%J�$I\ 5�@ �8E,����G�� H�ď� C╙��J@k&VN\����n�"=����:�JmJ@�cz��X5�6b�2ݠ�Z�$0K"��~֡t��r
`�����\^}��sno�o�:�L�{���lC�%V\BH�!6�.#^�d�)�w��+4%�.���ɯ�g*\b)C��)�<�w�yF�q@�_1� ������wN[	4���c�<%.�.�4b��"���o�޻��}�|�S?^����-���A!+7��.�m]+���@	���yV��mf��O�֤
�� �,�1c�>Y���ru~C����<�ē�J���8"$�Q��
���G 3ԟ�<�N*V���-`N�q��_Bǎ�ghW����KH���O��AN�'N4������Y9��cf͚cv�xB_����a=_1�-+`bq�F`𡇷�*�W�|���>��ɱ��C��I�<���k�Y�|ɗ��7��,�I�?$=&/��3gh<)��8~�`
`&%��E��|���c�f��OSwbo���)`b��|/�*�./L'��� ���;�:���o!Чv�vW���zZ�.�/�pJ�0��ę�:w�<�}H�0ڼ������LH0y99Z�ډ$�����Ӏh�܇��>nu��A�7�.r�Xb@��E��xq/s@���]GΓ�Iޡ�1�
�V��
xn�{�Z��cM�Mͱ8X.�r��nn��,|�L�Ǿ���}���vN�m���M�Ͻ?+��kJ� ���XvJ�߅R{�xJ ��yRT-��g�Y3g����5/��5$�����7��fiK'���K���0��ݓ����|&��;�g^x�e�@Ϟ��
h��WA�XLb���@���:H�����<��	-�F��X�B������3��<�@���h�Y���3>e*�ڪ��|$�m� `�@�f��6߽�{��O>�p�=O=#�����}P�cRI���Gl|�3vܑ�ѣw��[:1;��9��{��'ߵ,Z���%%�EDE����{(`R*f�I&>!��Y�3م�V���j\!�t �֭� ۽Zߒ�1�|MϞ3G s�I����Zgs��O�m����Sp$��3,��E�T�V�-[�{Hz�0q�[�{F��;o��K�#`&&� �� ,�e�ǝ�۶),?l�p��I�%Y�546�M�m�O�� f�\��y��&X� LΉ�U\LX|�����}8�0�����#۩����׹�~'��t]�:�9ձ��|�X�?%��y��z����Z��˗_�0�|��
0.��Q�;L���{�Q���^��q�^�&ªI�e]m�Z�pՒ���c0��a��
����%D�7@I5�^ &��s���v�36 8���Bi-� E) `������!��u��w5���=���cj.~��L�'VG��'xd>�Η��ϐ>��zN� ˜�	X��׿�L���V'��&���K�Z��oH��B���:�̘1�def�IEE�9NXVbJQ�ߵ�j��K�1��	`�W|o=�p6'��SC�4.Y���r�p����ơ�4�r����w�(�I,&ֿ��뾷�Ѫ�4��:=�w�Q��!vKc�<o薖�U�@�߭�9!����3�k�U�߼��b�x���SPX �H����@��:\oj���u�<O�$nll�,��O��`���=:*x��cƆ�f��޺v�ڿ��<�ē�J���3��?/.)!y�a��}�a�m,`R*x��E�5Cx�*��Ӊ�0)i�f�ZL��uf�t̌LuU�P���>��ɾ��گe�#jhP��z�C� �	�b=����i2Ҝ�s���K55G��偀���
L�葈�8&��ˋ��x�R�=!)��j�|�&6m��l_���1�/��(immU�,嗸��2)`��ޝr}����L'��_��v����𩳍���lk5@�}юLΏ>�� ̽
�].^��ĭ�o˹t����ׄ�tpG[�,��S�l��$ƏU �qb1�f��z� ��L��\�����BI|%�g �}�ٌ5�{�������jm�K�1,~��L�r�|�`�]����� �z�'�0 �tb����E��r<(��S�=��]N'��t����/~���a,��/���1:��5�������^~�R�@ $ &��Ӗ ��x��,�r\%��v뭚��i��0�mۮnm��{�ė�'�<s����ǵ�_��g�'v���(D,��o��-4�^G�V��HO�� s�|�����:� _�F}.n�߯U��|������ďS%�Jxp�I�d��S
�S�k�ЖG0�546�Q�xo̱��yq\x䂬��py���������9O<���C���%�	qɃ��xG�;oX�(�NO:��c�\��l��������jF`��C���R3��R5&��q�P�=;�~�}�9Gӧ��Z��ɩ��u�پ}�Ƒ�c�d�c��`&$'jaw�к�z�*`
X�N�"_Ծc��;Y���{��eje>r��&�G
�����2�Nb5��S̈�#u} �}��K�z��.u:�ì��6�����M4�\���h`����a.�N`t,�MǺ�ܧݦ���ynu�XY�ߧ�kYg��c�<U�Y^b�f|`Y�=o�y꙽ڣ	B=@^��	���S+�UYW�E�C�k�bp��%�HRH�@.rz�p�]�]Nb� o���Ì��5�rS�488X-a(�$�z�C��%b&�>"�E�R W.e� &��XY�K�#����� � &�&�Xe{`6��:=Y�`�� ��)?�x`�M�V�ϲ�=�s-�@O�I�Q ��$��$a	���/�O��_4(?7W�� 3����h��^$�Iw�\[�@������	�
�0�.r�����k��G�j>=��K�??a���|&�PozT@2�~���o���X+�x�I��h�ܻw�9���
Gn	Q����N �C�Iu{�0���ߨ̮�����M�N-`�.�ђ��A?`���w��<� f2ȟ�e���zجZ�V��tO<I�'�P�3.����!GEG?���[_[U5����g��y�'߶8p��3g�</3'3y\D���Æ&��?���I'*:F�	�~�1���Mڄ�N�,���9�I������ny�[�����)`��zX-`�v'�f���u]�p4Ja#X�#75]3��"�0�9��T3c�L�+W��$j=�ظXy(v&Ǹ`��ƒ@�*/",�@ .l�=d��L�r�޷Q�R� �H9Fb)����Ùvx�cY ��{���o�w�9{�f���'�$�ȋ��^��UU��c/x��� /y�`�$��X3�'+#C�Ǆ���AA��/"��I���kƌ��I�"�d&;��\��@ .m��Lc��,��R$�9VE��"�E�ո��V�'�,履zJak)��zOG@�8K���O?Uk�����>��1�oZVH�@z�˽'�i�9�o~�+��\�K|�L�1���2�
X0����4�8w��x͠Q�4N���Qa�岥K�w��t�)���+`��ڢVG�E>����?}�i��=H���pB�%.��?��s�2M�oz�;�]�w�3�g(U�=W�I�"������&��"���N8��<�y���O�1K�'.r f��q&8$����.�4�Ѻ��z��aӧO�9�8������3y���oRe�/WO<�]jjj~8mڴ�'ON..+��1��^��BI���Xy`�~��.��V
�MPW1���"�p��MH7��,�/i�Ԉס=�-�9k�<��+����+��(M :`K�6����'������n�I�A�%� Â5�$&�h\'1�d�'%'�!Æh�cqq��2�k��t�	��G4���F���'�������{���Z�t����{5,�$� ��lu��Z������/�� ����Ӎ�9�D���hz��5�q�2mK�$���XMHf�H���w����������Ï����1�<p���5�,v|����H�UN<���#W��:nROO����a[`Xqg��f&���zf�e�6@��ĝ��L��0��"@J[(PJ6:�K ����#��|`�d{�����
L�d���5BmMM���4��	l�g�W�Ͻ+�-s
�8��A���r})?4��U$�����Fo< &�W$�{ʵX�b��̽%��I����Z�����J��ҋ.ꬳ�	�2�E�`�A-�t��;�
d~h���B��߫rϺ�mQ`�8np\�@%��V��������wrK_��]ǽ�{^�u��ؽg�>��$���ߥM�9����;�q��օ7������H�r�n��|��G�>���g�+�ӽ/=��(J�d�O��J 3$l�	c��,*.~����19֚���r�\�_^x�O��_���ÿ�K=�������������o���_��C��S�+�O����[Z��7ђ�ӦmLIM=����?bzg)���Z�F��Lzv 0�E&��PP��f�/")���.�˗/�ظS[W��Ƀ�z�@#BJc_��PII�Y�v��B���"ȺtMH�6��p��yY�^�Z�I��"�۩�	\��������\����xX����^Z��I�W��8F�o��}��c`D�U"�h�դ�o���Ym}���$}���h�#��ߔ�����~��w�Zq���㭷����=�P�f"�c��&.N��$V���J]��&Y��ˌ���n%I 2��Y�0�����p/��8'��S�Ku�H��e	��!�%��B
��~_+W(��X59�t
��1<'`I�+��E�����5��9�	(3���6 �#��8J(ĺL�!k3���i*���2�0�w�zwI(PZ)�%�1���{����� �^�P�,�Co����D����7�Y���z�d.�G}L3����v�1e�%`�,œPZQv�����G�K��t�w��G},��h�%��;������i�,��̠ѡ��6II�&��hxd䔑AA)7�xc�E]4�.u�%���
D�Z�
�K�!/���!��k��⊟���������������7H=�俵� ��E~�L0�`��ꆠG,�3f�Ծnq}�N?�dhca���6I�ij!�?��H�],@6�$�$k�L�|H���M0�5u�r�����nF4b!d_>f��OH6EE�f��U�:,� fv^�iഀ��(@׮��f�m��D.���z��r�3gΖ��H^`�ZW3.!N�@�"OJ�~ ��n���#�lD2�X]S�ЛЇ2�J���+�����=��!.~�v�w.�iZ��tsw~�;e��ud�=_�c>����-�i�,W�u\������%�y�5�	\��՗���p�y��W��~��!�ځ7z��{��@����{��D��a���3h�@��H��d ��u��^y��&:2Rc0�J��M��'�VJ�\�H�P���#D܎���@���$�ºl�� ���w���
O�eH��r�ƍZo�!��lc��/j��6���d���_��s��}��$		� ����l�ۦU����)�#N�Ԟv)S���˗-3�f�ҘY�.�����w��XL�s L�ӊ��5��q�J��vK�2�ڛ &��U���=���!���k�+�ʇ�(��}U@������&&��U�P���;�N_�t�7�چJ���#w�hWVY����N�m�U�ݡT���3=n�����p������~�������)`�~�-^*�i���]K�{i� fXx�b�nʳ��[o=y���p��>uŕW����K
��Ce|��P�KU���d|��Ds.�첡2�L����?��aU���y��Y�39���O�?��cO<��%��5
��g�Mnjn���txt���łYT�Lb�Ϝ.�'�2��KHN�Lz�IMMxK��O<�ßy]�������C-��Y�f�<$j�AM!���r0B�U]��B-��X�y����a٦�-�CBL����Z� �;�� &	F
�C�K���uf�D_{����b߬]�эe��	���F �^K�ׄ KScS�&X�������x��K��|Ȧ�50��f��%J������o�K���^���|ʋ
�^�l��f�� �&�r�@cXh��HOW�k��	 �2z�a���
u�������}O/Z��vɂ�
��b")��t�R�Xby@)�D�:ˁ6�֊��ᖧ�;�I�+��p�c����|B8P��nk(�<~�)�-s�0q]����CםW���>��Ε��i�w���S�����t�P�6M{�Y�p��"��Zh���Z�`b�^�|�yv����^���s����^�t*�q��$�`��e���;��Ҙr�Nw�n���]߾
��穧��/q��U��z��PzW:�v_��&��$@>��p��~��!�{߷�9�S������wt�A]d��96"Ҍm��J��/��"s�|����G���; `�� �����{>��Dߐ}�.�_����ȼ��u#2#d:ʯѲN��#�w���e�G�&�����2�����X:��kO<��b0̎����5����&X��� *,����(���:'7��mȶ���Tw7n���Ty��1��x\c&q���//񶶩f�  	CQ1�
��n}L��k�.�{�AX}nwz�)�"���Q�(N(��Cs4Q�ރH����r���ʚ�IڣkG@�V�0I���>�l��Y�d�bb��0�0伒L��qZ
�XR�=��	`2D!��g�[���y�
�R��4pi���
|v�t]��W�|��@��l��N��s�v�s�V}�|�雇��! $EQ��u֬[�֞�_xI>"���V���;>^��
�.�{��ۀ0C�
` ��_�d�I1vyX������<��ڝ����������Z����g���1�X�I>^p1cu$^�,u���Thk%��������^���I66Y�X���4w�#{lnu�{^�u��"'�����o��X�o��F��X�n��JKK5�j����+QMu��1DGD��K&0õ�:͇����%����)``����ȥr]�鼗 ĳU\�XӶmߡ�{7n��p�<�D��~�������H/	UN�jR��rS��\N��ު]WF}���7	���%����Z���C��|8��!Jx�x�fϝ#��Y=��}�qF*۞8!`����ͧr�~�=h�c^?@8��Z��pb�){Gop-���9Si�03�xy����|�\s�5���.Q�h3�'E���T����t �ii��
L��ؾ/ ���&�^%ۮ�\!Õ��*�5�=�dy�h� ����ߡ���2��+���w��Ϯ��j�zz�C��q�̶����ꍑ����y��@i5�Ԃ� ���J���噠��
{�#Ni�	���
WW�����7(֘�qc����:E!�Z�&ƒRA�=���%�ѡ��A�wXq��9����)`�,032�M}C�|�� �z��0������	`ҵ#��@0pK/=S�����mҒK$Q�3&6NΣQ�>�6N��\'�ɋ�^1(�>x�`ͤܳ�Κ�����ʁ������ŝ��0�|eL L,�+V���O^���aR���=/���F���Ux�݊��!�ցG��@
�i��fM,a�'�� Ӿȭ�����N�b�q�c]I1t`�5����xL�~���U$��"i3ۭ �ZSR�S�E�nTIB¢yP����a~,@K� �k�y�Nu�{^�u�L�ob|�&ǌe�M�~;2�}��x^}�5u�764h�,��7���$Eq���656j��������� 3*2�̗{e瓻���>�{���{NQ�&�S>��Sj1r?���/��u>]�����6���w_��	l}! ǎ.�ǿ0�>ﮟ~"�
��8!0������g ��A2��[=��� �5��f֜�f�ܧ��-X9� �,Av���I=o�����	K���;��_7[��0ӻ�]�Ay��י˯����KU�NQ�7U��٪�����B�@!���d�-�H�9$��bZ��J����	Q\�%�^�h*�)�M�h�L	|^%�?��s�y��z��7��L�ȟ��'�?��9yr[rYY�ƈ��ã�N���Ek���;.��<����ZG����XSZZ�Y}i�X:ѭ�3��<$ Xo�E�x�5MM-f��)�H�Nqi�y��G�s/</�9
���%�0��&3s���u��Hg̜eRRR0'�OTW:}���������tϐAjA�Ս��$�7J����B"��O��ZSU]�� `r����)m&H�y�=�������a�M��Ͽ�\��,N�B|�U3s�,=߼�]��>�-4v{�w��.���]�ۺ�������m�w��6�X�q�\s���Q�&����̒e���{�3�V��|����&�2��ǎ37�x��L�F����(/W���Er	�?,vH�!>�6l(�\
���5�q ���.靆� �,|$�K�5
�t�X#��b��Z���f��j'�k M���L����l�}���),s�u�cU�)MDS�K崶6K�zHx��(-)1���	�X���k�m�~��oK]����n�>Vq�_t��ENBE�۾�����.φ�;v�I��9Ֆ%"�LR�q�*Q�X#�5��U��|P}�����$b��[���8��1��@I%[5���RJNU@�u�Q�9`�w����Հ��~�2����Ӣ<��o�d>�;���y����C_�s%��& r��ɾ�2p��~P>��n�呭�g����_��H,��:a����7c�#�����]� ��K/9Q�6U�s���mϩ�_����N���J��(�#�/��VY~�,���M2�O歕�g�x�5�H�ɟ�%��" ��������'�	�Ĳ`��#��^r�Nn��/z�CĿ�l���k/> 愉0I�xd�
�|�,=^�����.,.���Ɉ�F&VĻ�}y�б��P��۰�̚=�PS3x�h�F�B^^��8��:����f�0��'��@`�V�amniU7��e�C�0��,�߄D̱�_�n��`v��=88D^����	�����ca���(C���ݳ_΋x(���{2�}��x�;t�C=�C����m:��O[�Ϸ�ng[N�ܯ�^֑v,`6�4���	`��p�b��@����:[e{^��f�GƸ�c��7ܠ.p�\b��5�M�j-\h��FT�L���&����d
x��Ud_8� �����5���$���C�%pI8	E܁N�� i_��@������P<��t!�~�b��و����eN�Ċ�.�/�ä;Ob+I�Y C����V�Xa(ED���=���7��6p��� ��}N69�;�. �LY��������Mǌ��G5�n�n}x�cg����!�����Ol��]�|�Y�b�Y���j��O-��~_?>��"��q�Q,�V) \\���E��������{>�+���)?,,@q��ʢ��������vZ�lj�%Av̘n}�1��[o����@�×�&ʹb�$��8m��N��y��]��֏��7?dV	�/X�ȴ��٦.�L;0�w�@�) �v�;Wڛu��S �4~!ÏD;�}�F�Q���p�h�l�#�-㙢����2}��?���+���COϵ��w#� ��|cdT�a��r>Xqn@����G�_P��!�XX�� &�<Ѐ�6?�	���SI$�t2����b���Y�f+`��{��'�vW���2'/����k0ٞB�싄\� &VLb2I�W-���e�� ñz�5$]S���ҥ˴;��|I=ŦX��#�2235��}�ѡf� &��|H���N�V)���f�ꛙ��T\ʝݶ9 ��:�=Z!�r����/��U��v~O��4ߩ��e��% �	q��L`u�^y1�e{�����d� �t��[@�D�Z2��B�"`�X>��+�p"#"Lnv�)+-U�$1��7g�}�L\�$0`u�:I���n�����$�K&�I1qb+��$V����M8���
G�'1���L��IO�̼� +杷߮��X�����(�rBN�J��:2D�g�$��a@�U ������P)�n���\�c��M���{p�y��G�[6�?����Q���~&�y���f�e>]��SO>��'z�g ��t3���$z�(��O�@U�@#��lu@�f���f�w��$:��g����tv�Iȱ���v��o>�3�gM�|D��:�5.��W^H|C��c8�I�*�XZ��-N8��ݓ,�t�
3G>L0^ZZ^�a\)i�&*6��|0ﲀy����sܭvYO˿)u�׭��j�J �O@�iY���aX�=$���t���˼�D�I�נ2������e�n3=���� ���^���bcT�0��rr}�������<��V�]Ă��|��'
��"��$�Rz�Ay��c�P4�D!��jLf��h|�]�����!�
���ye��ll|�Z,)ľ|�
yx�TH�KI��)O7�@)�a%������D�G��2�8��K�C�/Q��ZIRq=�f�Y0�L�@3���r�uJ���i�%b�x���ڇ���F&>��N�Uï���u�����\ ����_�s]���ַ^$v[ǭݶqL[��`b���Cf���:�r ��g�l�/��7�)��L��+X�ps��.��Q����d%kI-D,�ڳOp��Sd����B��`��.��z�����IV![��v�Kz��P:�;�� Q�(<�>N'lk�q˙��Ӻ�s�ȉ����Z�N�YZO�߅�D6��J���H �RI���Y��ܹs5�|&Yх�ڶȗ�L`R�R��ʤʋ����ozlj���urn|�As�̆M�w�}~u����nDYW�r�<+��EK̂������YBO3|P�x��:]��GZ=,�V��j��"^��(�lG�q�ӧ��a���2�pL��<�z&8�>��}D�M��ɞ��N!�&❉r� �M�,�y��=�>(���z�:�����wJIY��� �	&2&֌�g��Q��,���~�
`���g��cB����?v��d�?-�B�eX&��x�h�h�l�)����d���O�9��IO>�G�1���Rߒ�>��Q�ǫ�b�$_ȸ�m&P����.����j���ի̪5��a`���<��b�9\��"#4r�@#G���G���&<<��516.�$���F�[���.�U�D�����أL�T�x	��d�Q��o�1��#�J�g����+�o:f�Z&���ɴ��\�H���E`5D �i']{��+��^ ���f��gb��['k9Y���COy�0_�p��8�����Ow�<О��qڡ0y����:f�З	�&ĭ������e����˽����w*X�%! �<Xݲ$�`9��r��a�J�q2��0�No�vXI��=\�E$�$�)�?�<z䈂(H,�N��i=�$=�w&m�$l�L�+%��A\ܔ��Ir��/�$��`�$+fkk�B7���:ǚKԞ�{4!��Y�7K�& �	�V�I\5���\'��Z� \�n�)�z}�Ft-ʺk֙�+W�EK�)\�l��Ч���3�*��_}�y����n`��Z��G��c�s&��^����]�f�Z�i��Mb�w��D��c@;�����P�mC8�O2���$k�Q��ܨk̳:95M��"-`^w]`
Xu�s�n tB♪�ݾ(�&@��qJ&=%p��_w���~�a�����e?��^#�~'���(���ճpzrn�fmc}raQ���Ȉ��G�R�4q��w���� �\�|�B�(���(;��E��$�6���M�+���L���4�I))�ƚ8O�xPA���رᚸ��MF7�7�f�5��LpLךg��Y9��� �8S`q�� p��7��A�d� ����1��h�傢"��1�Я-�L������QHh�&͘9[_.u�~�����	�*I�xPZ�����*���r���>�u��a����>w��k���c9���@۸�%����*��$ܓĩ�3I_Gig��S_ߠ�y�-����,��=�2v���{kfvv��KAv @�M0ϕ _��qw#	h��MV5���>YޛX�� ؛|����	��e���N���7,��/\/�p�>�I���7нz�*m nv|t����f��Ӂ��T�@���H���b��iA��.4W��23zt���{e銕�D�UkWw*nn�U}T��!y���U���r(�\,���Ss����V����?��������s\>��f}6c]�C����N�ӧ<���2��ٲB~�Ƕm(|R��j�c�IYK�U���AI�����͜���2˳��0~df�DyG��1!cǚ����_ ��|��(e�}#
�Y8t�����^h]׉�u��>!���U�ʏEߔk�Mt��k���Bَ�H�_p�??�����w�����'=���O��X����M����(�wx؈��9��rbF�fDd��Q/Y�L��Y�f�� �0�,C�����^r�ٲ�-a���2�8m��@ �z�ԟ������j���^IY�Z/��[ժ���M,�0��	��m�~l���VS����|��l�<ŴMmW�&��C�F&	N$1/.>��s��\�$͜=G �s����%�|��^�!�E�(��W ������y1���+�꛿d���ݔvV���֙��`C�q��H�ܧ����ul� 䀻�V%�k&V2`'[>� J��H����E�}g�}���>۹�׿������==Qd�,w��������,�Ȟ0�,^��f��7�=}��ԳB����R��ޙp��π�y�0�jWWר{�w_-t�N����T�E_��͗gL �dX�y�>:}ʇh�:>B���l-v�� }ׇȶ(\R�|����`ұ���t���>�Y�מ�Y�Ē�h��?q�����X�ۡ�9`�ׂJ��y�̞3O���7Ż51+��'L������_[κ�@�u�כZ`t�{Yo�Z�i�q<���r���>+���>*� gх^8V���;��2�:�_���K��/DW��eӓ��@�9t�M��ǝ��M��m�͝���'9���M�:����Tx��m�͜5�3�qT�h�7,���C�&C���?冰 ��k�Bk�|����k�QCc��3B�6l�@CZ�'�I�l�������l8�NLֵ54�[&�6�{��zL 3�S��X2�Zz����K�G��X_7o�p��%�0D���]ݶ)�g`���a��E_������d"���:���OX�6���jB�@�{�/��x�n�<����_ /p�E�TAs�rSUU-��ʂ��' DR��9�~��
� 9L��:��+�
F\��=ty�b����k�9����Ab.� ���t�
t��q�;��C��%�p����/u�����rF��V��ޙ��:Lُ�%*/T� .���yE�z3��oXa�S��_�տ��ۂE����`�uђ�ju��F�Į?��>}ħ�տ�G4f��M*��M��]���X7�{72\o��\��)m�Jo������ԭ�����󹔎�c�@������ꥐ����o�k�3��}�V�����I&]��qI)&<z�	�w��;��7���>�\	@Y���*��#p�H-�E��h����j��v=�\_���gr.��U�-��f�\�f/�e�2}%�M���2�_�lz�6=9+q済��C��Є�i����#Lvn��>s��&_�,1j��7�b����y�gU�����j�����Z[{C�N $����ބ�W�ao�)�ܢ�p�*u���[�NHX��?�y�7'�7��m˹��u�s�sƻ��9�z�F��x"�2 �ĞN��)2�#G�d��o:i�,`q�U���Ţ	2����mک[��9&�P�p�̬���m���(��1q��`D�)��I*�n'��%��!�g� 3C���Hghot���^�k:��򴭀)�E���Ĝ.X�H��6n�]a�|m�)ж�>7�f̘i��w�;|ҤIfܸq�I� ���0��H�a�dI*2?����9��N�0/d������Å�%�����ѸJ�����/hY&�IQ��X���MN�),��7�|���u*�n�խ[!`�k�VD����d!�߸�<�A�a�F�MfCY*L: Z��@'ceF;ک��?�j��ϝ�<��aG� ,'�����n����
u��랻���p�o�Ā����ur���;0X�{ʑ���Lr"9ތ;���s0�#��7i�6j��?x��ѻ��Z�������	��Yd��*�v+�
�y˓�*��F��w[Y
���!�J�c��e�ސ����7H��2�.��D�=Zt}�5~qq�ʋ�yMssr.�6mZ���g+`��ݦ�&�`�$f�,rb&�h._�R:��>W�ۘ��ۙ��i�ACrL����(A 77�b���X�@��8��١CgM��UM; ��G:@@�n�V�˱�:�X4X�ˈ<���320����;p�����S`��ĆR"�'`����k��3q�Ϙ5[-���L��{T��]%.`�6��z��r����=K�қ�H�,����T��K��~Y ��+}L���*u<�1���+��5OmT�Z�� t`�2�m ��D��3L���4��,qb+����k<1!�$�l��\�JL�^Rx}���
� �*��"H,o{E�~ߓ=����s&�`6�- �au$�b^�Y�b�f�oݺUǴ&��F����d���,�� ����Z ����6�GΥ���#ɧ�<(O�6M����LrjD^����(���۝��-w( Y�e���$�{��XP� !���M `�,���c5-_��
�n�]����� ��W�:�/��U���9�|s��U�\�z�\�V�vj��%�*�-�Ϭ$t�~�%�-��&}1�&L�lrG8�w���S��r�i���y�l(�ಮ���"���U��V4˓�Y��*+/��J�@����%��;��jݔ����ߕ��Dw���n���	�̃E7Ԯ]�j��_t�_�*�,`ʓ~θ��Ղ�ݺ�f}3&8	9�,3I�I+X���������M��h���&��|J�,�Y���P��X� g��Y++DK ��J,�@&��� ! ����@$�i�} ?��X?-`���p��	 �p�՟-�L���n��Z�hʴ�Z �k���U>�ݱ�9��]�հ��X��L/7U2��w s�&�[B�޺Acmy��6�A`��ж�f��$�P�8L^S�:�Z�H�� 
�`)�T��h"ʷL����^Ѿ��d��m�����I�$ ��S�f��%�����̞�_&K��E�9s��>m�T�,�$S�"�l-�CĮ^�F<@��-[kȷ��[4��4d�%I��a!
�`Q`m��6����F�j���D;���  q��'`R!�2o,c��U~��7�6�+[�ñ�|����2���}�w 3g�S�k��V�L���<��܂f ��*�v+7�ze!�,Y $��JA�� �V�����ۼ�}�9-���c��r}o�p�����D�e���c\I�#�d�l��ũ���=n�@����֚���@&`�Q�X�Y@ ʟ�_�~:�8�#�7,�dfyX�2 ��B��u�v.Q%N�ĝN;@�䘼�-P�r<@p�x��� ���lr�y��l}|��?H��R㓢��G���Ly?�0p�ƒ�v\��I�F�  J�"�s����ܲV:>ke����i�NҁS�Ȫ^&�y� ���0���O�6>���(�R���Ƴ>���׳�]$�r���S̬�s��+�3ZgV�^+�yK�D�C a�X'�s>�
��+2��U��$���L,��Ժ�X<َ��&�K����"g�6��C�*�~/`�L
�s��"y�w��{N�-o��uw�M��IWh��'VK�Y�L��գ��<%��,5����`�<[~�r�J��5f�-�ͪ5�.L�/����*�c�n� ѦM���pї�B���VU��R	�+���ֺǽ���[�����˾���'в���sL���8�>��u_���m� �!3� ��w@ƪUk�p`�50�a�'�G	�{W�.k12�2�ۭm�
�V^��*tZYдX��`�|U`Z��l2����}!�ޔm;e�V��Bϒ�a򺶼�����ث|Xqq�89�̉�'����s��G3�:��D�z�Y	��Q�����mT����$~xc־��3͈Qc�:�VY�~�y��N���n���(�-�J[Tffb=m���x`v�vX:�Q����t;�J[��p2��x�\���y�0�eHJ��`���]:���_-7LG����i���VI'�X!���?����͇�/FN��f�|.ר��rZP�<�9u�4u��
lt��Y�cm��ݪ��ұ���Z�z� l������۔-�}tDĿ%��0�u0���<�'�~j�o�n��w�z2�qy�@i)��t�lC�22t���R�K$�T� }����%�y��ú�(�S�V�#�����x*�r�np��B �\�~�Z�W��[c��X���/J�,�.-{��D{��.����/�R��2tm^9��j�|�����4��ܲu��&`ic2�o�K��L	��ٓ�.�l)���WSrjԨ���m�вTY�tZд�+6�˓L/hz�ݒs��s�+׸K�+��&���r��Zڅ���\#��//�j^�t��)��34wg��]����2��i	�Y�t��!g�z���$Z� �� �@�2�w�F�2��XrL��� ǥt�B,��8⦦xzrj�!^�߀��&097�-� &VI���# ��X>��D9~Zz����}����\�#F���Eä�j/��}����8�19C�a�0S��d�Q�/^���Mj�
�����&Kg�'����t�~�tޥ����Yv�sw���
���y�u��w}Y��Ͻ���C�QFN"hĒɨF�F�V�QȜ$��H��)�&��� �r@����\&��WS���@
@�P����Ӻ�$��5ye�ж��ݷ��;~e��mS�r���6�g�"� ����#���ΝZ�s�޽f�<�QF
P�X|2��ݲ� V��$� 7T��Wn�
�������?X��X<Hz &�Z� 'ә�{����Z���nS�UT����r�|ۜk�o�r�WJ������[�P�`6�������Wu�y�m�/�e.�����3d9?��<�gZZ��{���R�d��0P�]��3ޱd�RI�$�!�ôDEֹ_e��J|˖&T~#@pY�zu��� �@���]�^�*6�r�&ræ�6�M����VY��]o%�+��9#:*���Iy����[�Z�G�<=X&�� h�0����:�yy��7!g���;�w�t4�U+�{�H:`���C8NW�y���LR#3W �&7f�X�b���]ǎ&]�ɘ�� �λvx��S��fg�2ғSS5�cؘ�.]�+�b�2�.���"�2d�k�(O� .�O���0�!et�>�����g��S�7q� �0}��o����<�S�W:��X�?��e�:b��^f��(�3[:���'� s���ն��/��%�{��_�����/��#{���gβg��/Cz�E��6��<�oz����� �����i]�f������:�,g�O�8=��{׮Z�r�ȑ
�+䜸b��K~'���E����Bl�f
���|���jW�cT4}��{�T�h���0�`Rj d�$�Q\���>�lp\�X�~,��GTpK��,�X0�Z��~�Y��m`�ϒ>b���E�oͦ�� ���F'�x��Ub����-�È@�ĨA[�m7k�o���j�z^������2����?�}u�J�_T��r6���!`���N�/�I�e�8m�b=��M�,��:����I��F�*�2����;(_$���6�.�m�ɛ�L�;wu 3S�-0CBB�j�jժ���;dhVV��3���W偧6�*8��M��@�$�p�{�����2�\���3�ηe�#�n��3B�V�	d�Y^_y�����`��Wg���9���ٮ}�������ѫ��]�O���B$�8q�����̔v$�S+#�H
���;|��c{ߘ��z�1]��=��ѣ4^o؈��.95E���i�6Y츩�ÌL�eg)�� ��Ի�H<�缨K����ާ__��r�=5��ט�ʹF�`r^ ���ɓ����䓮���b D-�\$7X��t��bp��'ɧ"��w���̵�vT�,��ʷ��q�ڑ�8�����Բ��O����9K�k���ú��J� N[nL�l}��a�(�Ƃ��������G�ª	`"��d����6��Z� p�P�29�mSV���VV[�>ж�N��2Ǯ�ۼ1�I�R��5��b�G�1o���y��53|���k9������$��S�/�$���KY1���MPn�
��2������[U�@Zz��}��cA#˚�p�D��xH^�|����C掻�6�nܤ�ɾ���/HK忣
|]�k[�d��7_ s����߹�������k9�z�\���d$��s��	���*�Õ�k4	��I�3�j��A�9=f~t�yH��<��(p�P����0�tӄO��x�8��@_S�Js�M7�ЬH����2P�P�^�r�g  ��&ræ[4�6�r��W.Q���_�W,�F��aY��l�)������:]�S����.����������9�6�Nn�Ȝ>�����X qU��3@@��!fB�du?S�?4�׽gw�5  #y�b�IoX�ڶo+�&�0){�C�?b�H����P�����4�S�PL���;���-��z�q2�;wq��Lj35#M�u6�{Q���̡�B���0�s|b0�v���TW:�٩�&�P҈N3g��Z�@&`	P-X��A1��'R��C]!��2��2�u��1� �#-;�+�����n��C�#�YO;m���[�oK�q<���d��̓����� �g�d�n/˕�k	�/�~5�n�5���$�`!������$F��@�@�r� �P\LL�$U^������rO�����kh[E�Nm/o�Z0m�s�Č�s˚5���W�}�]��C	�9�f�Y3f�Y�_	$�̱B�]buƲi��Ɉ>V030�
`.Z�T��(�UF0I��U���;g_�>��yP~C;d~�����nHXs������%�Ҳ��:
p^!�y��?��3w��=�/������k�����6n��N5 y����p�Eu)ˢ�c�H-��u;��q���ƶ�q��vbT���<je��'�6�<����#�;��E�-`Rd��ڵwb蛷ha�)��x��n�9�Y����M�Ԃ�@�@��N7tVd��i��V^�ræ�A+/x�������u ��BtX�����!�R�(Y�:88���/�|UVV#]���'0�����ӻO��m۵-�����(��; `Ҷ[�n
iK �c�LIKպ��nj��=E�]��`RDW��q�;��+(���FRZH-��0i�]Υ�)pK;�W0� ��\��%VV��o��
�~���k�͟"�Í�x�d�L�
�brD��mӿ];~Y��rڕn��,ߍ���e]gۗlw�� �\v�V�nˍ��LgX9&.vʧ\��nr�䁤� >1|()1ѩs)�+ Q�h�|��W��=�W+%������~��i'�2�]W��Symm�Hީ���M� ���8�,� �M�&
��2D�E�c �3}��t�ĉ���6�֒�l��07�IL%5]��a�dXCF�z��}��||�yH��ܿ�ܶ��[�?O���_���儑��K�Ŷ@Z������(���Y�\��)�ͼ���ܼ�Uz~��S�1����$Cޢ�K>WB�l��~��Q�<w=��y����cO>c��,p���v.�쨀�Q 3K ��i�H������u^��ЊT�z��Ve��[^�,8Y5�N �$�^X�0�J�rY�x[�}F�}P^�"�GD�e�0Q+YNֹ̯���E-���SN�\���t��}gv��G-,tX���A~�̛8E��$6��ꇻ;W`��I�PkN�@�P6�0��o������urԷ0�<�Ӵ�2�U��<�9���}{+آN�uJ'���+�f��=M� EjZ��,7��}4�t�.���K	��ĉ�5��6�X�r`�ط�G����&Y�3fkй�"w���I,"pI2�S��+���'q
���ݶ)��"Y ��[,}�-��Ḥ�}�+��dV	�������]�K�S�dxH��LNLP��ݻ�־dr���SSՕ�xm�#0q�2�5�|*1e����Ӆ��e��)
6	��o	 �V���)�I���_���`��Y�ZD0�u0�L����������}�9�D���^���	�P*�R9�_����y��'�.�xڏ>��y���2�O�s����[7�$��������V��v$ː�H�Ġs�$v�4nr�o��߀A�����ʂN�6o_����_0g�/���M�S������6"޻�o����ZC��{�ӑ���#C�>�0������|��]f����y�y�k�fӶ}�o�5�S����������o:�H�hE*J��i�P�n������^�fe����UY��*���#�C��焈�����C�/���Y���\�u�^�(˿��_)Hl^��[& �o�Au�v�ӮC���2[���P��u��9y��&I>n�fqF�q��c�p�+`�͞�� (Ǵ#��dr����~�Ԃ�N�$�$����S;׈(�ۗġ>�MwiǱmf�޽\��U��8Q�p$�pn+k[���\+`k�1c4��`Μ#;.��RNr����}>n�����Ă�0�0I<�T�%b����`��7A�ېE��tƌ���V�
��A��kH�a����N2�ID��#���Of�^�4�������@���˖i;\�֯7wh��m�ֵku�" �r3�0y��a����� �+�r�/�^>����ɧ����'e��ci���cf�]��uo7��+��`6 �b�-gT
<�T �5����O?`���{Lyx^(	����N9&G�^}�<����læ���[�0��������Ï��v=a�|�Y��s�0O?��y��0�(̩e�p�B�_��Ws���ܫ뮻�� Q��B'��<(-B��@�Y�t[6��YhZ�!S���,R �,K�}9����,�&ˏ�u0BP��n+ו*�[����]+��b����)33��N�:��j�.'#3sgJz����t���ܴq{���j&M����z��L�c����Z��<u�Z�����d-i�U�XM��@我��$�t��IS�C��U`�� �c�M0&MR;p���5�9����
vXA�^Q�,q���::д�F�p8���/��y�Ӝ�z���Ys,�ƕ�A�B�&�z�t��	>���,I���w���T��[����Gֻo�.g��9ˬ��/%g{�u��n�z����&01^>�)r���z�9�ny�x*�I>��+`b#�7*I?$xԥ����
Q:_Y:Z4o�	>�i���}[V�";Yˢ�������T����+�T�v������|��30���� @��t�=;Y��na�D��R�Œ$ b5I"1�"��g�.]����%����`2L ��3��a���[��+,s� I(d� =�����ϛ����yB�;�������fͭ*�>_�n��V��>ݺ��]��f ���ʶ�}ֲ,�F�YFY0�.���]����z�|�]�m+"��C|�b��)�D�$�ס⽊�Hke�u7�M�ڳ}�������=d~�q��SO��.����͓���`N��Q�0;t�l�޴��Fl\��W����_��s�5���+��,R��PZ|z!�,�t�gE�N7t�nz-�6ݲ�門]@�t��V� �ʽ��r�"9O��h���:�r�>O4\�'E�o���%Sff��Z�����*'%5}gRJJ)�Ċ��=�������-���6m�LF�!�}ǎ&Q �ڕ0��d�s
�O`1r�B�09�0ǎ����`j�s�j��*���"��2{��k�3[�d`RW���g���íL��sc���L˗�O���$<`�\ߌ���nZrZ�B S:?���3� �D3F �;�_:r�,���~`d}��%�d��������K���U�A�'�Y丼�"9�	��� �(�7�b.�~���x�[���B�������T���&ڟ9sƜ:u���Ǐ�o��F�,s���gϞ��U���k-k;SY�X�L�ȣ�eJb�&e����k�,� �YYV�^3�'#.1�'	@?��h����߯�S���K��	��&NpŊժ��W������"�O[�\M1�f�۵d�cO<e�zV��������<�܋���&��fӖmf���Z ����5Zg��'֯�dn�T�C)s:�y��`�C���<,O0�oe�G�	�����t]y.7�~����;4���vh��#O<i�p�r��?_T��E��#������\Q&`6�����*����6��u^� P��[偨�O/��N/|��n�t�fe��ֺi��m�t��])}�HO�_(�O����[��e�FM�92o%�d���CP�'O~�LI/L���@�IjG��S�2t��<5_ "_�/״n�N�w���0��*�|�i7f�8� :���DQXTW5������0�t��n��T���q��X:խ.�7.o��8e��ئ�R�\ S�M-�r�����4�����L�N]��5�D���G�6���RB�*�e�,r����9b�X3u:	;�Z��VYYz��9s(��Z#���,si�E
����g��N�����~i8<?��r��s۔>��2 �8.r s�if��%�}�2�G�8��9�%8E�_��+s��$�CBR�gOb.YG�9I?�$˶�ͷ)S�]M eAa��ꫯ��Ç��l���g�|�M��k��W^~ټ��+���_7o���y��w���o>�:z��Z �k'����0��(7�u�
/)��K��s'٪y\�Z���}̉�%��7|�VL������9���̭X����-��Ń��,K6F��I+\��
n�v��%z�ɧ.������z��e��]O����ܶu�Y�i��u��f�������ؼu=�� i���v_�����,T���
�?j�<P����Yf}�6��5< /^&�9G s��X�.7ܶE��|�^�����mw�mw�g�p'���'�V���>��S��SC���f�/���L�K:v�,��N�>��63u��6�.���������n��ORy�Q  E�@�m�n�tæ8�M7pZ�UY�4��M�^��@a �����vٻ^����i��Ⱥ�2J4[�g��u�M>��CP��N0��[夦g��S�Ē`���z?8 s��#���C:Z���zΰa�� !F����o-MzF+�;����>�~�3V�o*��w�F������8Y�}0�-u)�
p��{А\�7Y G ��\��� ��h�] ��tL���3����X&L�� ���cʹ��2���s3�� �&W�h��[Dk���h�ƌ�=�L�9C;��^�t��`N��	6��׶�f,�e����=���~���j���� "��x�%`I�o �B&1�
��{�l�?�Z���Yp���ｧ����{��x�s���f����M������ڵk͚5�~W�o��x���r��^%���z�ٸa��ߺe������'�T�2�����G��z_��0���8X`��ܼx�Ř��|7��D����C�Z9B�Ę�硁�-���_�^>��I8� �1�����Mͪ[֪V�h%���D�n���n3w�A��#f��Ϫ���^4��s��Y�0'����D@9 t�����5�[)׹�W�{L9��3�?07ܶ�l�|�^��j���o��)�����Ji�DX/w>�� �N�qu0��'KS��3�Ԫ]��E �w�����o������N�k�,xz���U  u[@�����X9����@��nZ�t�6��i���V��nZXt��n���ݯ�2s9�!9�3r��\y�Z*��y/���-��I�0SR��l�Z�s��X�Xs*���T�_��`R�0�u3�F�T+fB�oԘq:�x��o�	�F���i�$"�������r��Fί��q�N]�u�|�=�@yMleRr���7p��%����f&N�.O��L_���M�'VT��ē��V8��y���i��=t�LR�$�S΍U*�e��9��D,�|V&�U�\�`3s�<s3����7+oY'�է�f��p�
h5R�{�v�0u�% �]_�,�����=�o}������R"��G��MJ^�~7�1	 �g��:I>�дd�r���Ǵ�*�
*�JGX��5��3��!w*���X����p�1OfY�����/Q ��7C*�|#�\�P���
�g�~j^�׿&�CJ�P��o_��S������F�R�?�տo_CR��,׌��&.��x�����iѢE���n3�	�RB�رc�Խ��~��»�-S�Y ��BC�{$�G�_I��s����m���g�����W��^�|�Z�S�֡!�z\�S~�[��DC`r��nV��J �/t���k)���&yŧ[HF��v���{����>/p��<�¿,� "�"0q�R���F�i�n��`@��,O�V��9	E���l��CI(�>���������K��������KA�]��f�|�X��@�\����6o�[�� ��Gv=m�YK� ;�S|��h,Y*����1ã�A�m�
`�=�ILSS�VM�k�l~��_�������7�)S �WF˒F(�Bhy���Y���m�t�4-l2/˪�4��Y�uӂ��F�,Lz����9�k2@�J�3Z��.Ht�/�����0Y�l�*+'#3kgzF��X%0�5T���*4Dsڌ��;W_�=`v�#5t��*`
0Μ3O�4��B �qƻu�)�J��P�Af��qf��|�<�,8����v����Os�@�t���9C0��� ��r���n&N�� KMM �8P � &�#O�Ӥ��ڣ�0q��U-�N����/�y��*��5����g�{\�f�Y�a�Y�n���6���'m 3w�p3e�4���s�f��S̛�+l;��i[���U�T�5
��0�f�3]2 ��>�+�`��T���&��77��; �d��uZ����ɿk��:�VJ,����ŋս�HCX�ΒQjV:@�̗���2=X*)HN"5 SSR�=��H��ٳ�T9&#�0T&pI)��r�YO�)�&��u/���^���}W[�d?�g�]�&�G�$s�� 0c�3L$V�;v����6m�`��Ĳ[(��Gl�ص�l��2{�}���۷������=�;�����r��\�$�<W	 ��?逦�$�䴗ߜ��n�( ���y�}��7O<��L�mX�n��N ��P��Ŝv"<���k�+`Α��Z����30�o�X�.k��+��z������	H�@%�L^�lDo�x���hI@��ݴ��^�����`���U��+�4��կ� �կ��
���g kh ׻<˳t�A3lZ�tge��n�t�ۚ�M��M7T��n��˹
�<Do����2�SG��̃e����~)m/Z4�SH��mڴ���n�3�U�Q�)+[ ����a
�X���9k�\3j�X�bq�B�;r���H�<,���2z�M���ޢ���SR0�7���Vț*�?q��~Vxs /W�9�6���Cg̞c���jg����VTk]�7`�0�V�p�ڴ��� &P�86㍏�s�[�H�u��ֳ�&n�Q�H!XޏL� ^>��}��+n�U�U��nY��/��i��E�. �f�R�V��/�@`���� cY�h���9�<��6�^A��6yO+��7��̝?W�����3fh@>7�kJ�8b�ek��u�߲~��&�پ]{K �Mv�&�h��O���G��t��I�W+�Xè�Y�,��N$���e�:�d�s~����X"�M �'�0�ڽ[��>��#��$������/�hV�^m���H�nݪ�O?�D��I�&1�;w�4[�ȸ�<q�Z5���3��I��[�}�ݿ2��>/`b��)72Bx�\1������{�;`D%b.�k	L����/�0��{�ɖ�w�^���)P��+���n�M���r�O�n��;��F�e��
��n�!�[�W,���m����P�|��Ju���IDA�v"`��-p�"x�O ��:������s��/����9���'8��|J�t�t�J9��
����m>����f�:2���^L��y�C���G�Kp�l߲�.�>�-\���
�;qjݦ��.E5�6U�U5���o�/~�������T�D�vˮ�ꪫTn ��AiY 굆��Y;���VM�K��^�6��ia�,�t[3+cѴ�B&
�V޶�/�)��)9�Q9竢e�jY)�t���r��˵�3��T
0۴��>
�QR�K s�f��0qQ�Ԥ$��&��#Gi�f_�Qc��<%��-������q� �?x�!�7%���'i��ctb0L�"�`
��	`b]�� ������n�2$����0)��6������$� ��;E ��0q��2�n �J�rC"}���r�C����w����g��������6�������ݳM^;VN02����* s�<B	&)`N�9SoBX�Ԋ)�YZ�+O���# p�&��v�X*���;kl_jr��ə���[�yzZ��cN7N��Xע+�E^фP�ZI�Gb:��!9Y�$�p�5���׿��X�}����e��	L�H�\��\c~oX��̐�-��| .PG��9փ;v����5�O����ɾ��>ֹc0� V�Z�&M��-��3�H�� �5rS%>�ŲJ�8K��_'7�Zr���ny/���[o�g��2H6�+7`R�ae����6�Y�u��ʒ�ͭ�D��vs���UMc��<-PI��.] 	x�}�W��t,"�X
�*�@�I�<[>'j���_��E��_����� &�>��O��w]`Z&0��+&q� %�!b�Dy��֮3s,��x��S��ٺ�<�����(sS�*��yW\q����~�s@�<������VF�P>���ϲ��^+gY��M7p���n��Ί@�,˦ۚ4���0��U��K�}BtP�����/��5�6���8�m
�ȳ���dfe��;���ʴ�lm:� k�`3 +�L�*���)t`2z ֯� ���f� s��E|K��0�%�S s�/�lk� .�΍K7��if�,LG
��LH4m4 �\9�f�0M�$7����;���`Ε DQy2���L�j��L�|�Ϝ��	�RF)E����_ s�0����`�n-[�V�Ar3�p!���Sҹ;*�����7�~>���&P��������.;�B�_�0m�<Ơ0�g�27�Zm��P�ZY�����`Ir ���o���:F��1��˼FM|� M`O�����M  �^IDATaa���)o$����N�� �gj8b%p��I%ֻmwܡEé�<�_���v
�c�˚��b!|@��y�����r�ĕ��(m���c�=o��7�55S��2Q+�c���hBPyq��r·zHc@i��K.`y���2�����G�1�v�2�C�*(��P�'�|R�0��o
`�9T�f[���4��#����<?�HC�4@���$>�ڌ�ę[�֥ �Z��u�ua���yȱ|ީ�
`.\�L�gΞ�%¬w����?�չ��
X��;�>�N�h�a�w����Lkɴ��gȜe���8^���hi9��i�0���m��N3Q���*7���.��rs�e��2D�
���H˂ϲ��nk�<˳rVƺ�M��iA��fe,����^����^)�$7<z�K��O�Y,�8+�c�s��|X�E3G�D˶�	�\�����,�`f� �"�`�r��:̤�T�^n�d�0����ƛY��ka�Ν���-Z���dE�LBL2�)9A����$#�����̉���<����1>���J"��n�H���Q@���d�RH:� LΣ���Ԫ�6c�0S�� &V[,�$�Xn��8���58{��+p:K�mX8�97g�p�r=G����� L�U8:�����w:yG�ez���߶��w\��A۳ΞǑ=m�qKd۔���Ϸ�o�L�3*'L������z�|@&7@70VFĴZ��^>gj�R��yl�B��2g=.s����sJv(SL�X� JYc�۩<�
�)`��3$�`5Ed@/�7��{������?T�ĽM�QO��1�6����Ʃ哲D$���<xP3�?��cu������={����ژީH����?0��}�a�EF1���}bY%��渱c5.W=%����3�~&e�ȉo�^)�͵�}�-m����rs����S����r���{��!@NAv��8��^?g������r3s��݀I�P�����������EkAt�s�wk��w�U��E���1��d�|E #��@�i+��:9��dZ�ye�>\#I>/�>r�h��/���I������>����m%�y� L��N�6�L�fb�9?�车��B�u�[д�p����H��̹�&1��]��T/V��h0%�3�Ʋ ˦W�6^���"�,<-t�����fY��@VN�u�t�۝�M �mݴ��ܐ�M/p��Bf ��.[x�e�=����>,󽲼]�+��6����J��b���0� fdf�N��:�9v��L�HJb� 0\I)���ܸ)Q4l$�@9
�#G�33f�ӡ%-`�LHh�ঀ��Q�?i�#㉧	`R߲[�rΡ�N��J�"�͓+��-��B�� ?`��(�.m)�n��J �����#�JS�� S��Woh@��P����Nw �U�I��.7��r$�7
'f˱T,X�L�Ry��,|e��s�6���,Թ���߶��w\��A۳η]�c�ud�[� m�d�=��f�F�Lꅎ�&��̭r�ͷ����Hb	0)MD�	<X�(I�:-O$d/S��E�L�0t�0*�}�\����'�6e��5�� �'�"h����/�T�ܴq�Z8�����&����L�鬜�F&�@(I0�O���Y�uX�g�yV��މu/���fe#�9m����|.$;���Ռt���
b�t�o�k�rYI>X��'띸�'�)�����-70����P��}���RK�ubT�g%�����@��q���E`b���p�<�h�@�Y��s�wk��mf��{0��.#�������8y͑�3������H����
9ּ��ʹ�3���|��\��%�[�G�������o9�,`N�2Ɍ��2l�H�^Se���ZaK@����W�0�(>���~Q`�pӍ�W]}u�@c� f���9b�W�m�fY
�V�k�t[9���N���m��Nw���p�A��֢ia�"��Ͳ,�^д��i�HT`"{9�iѻ��M�5V^3�y�\�Mr�������`�E�����ty����VG���9J,�j����I��<��LLxk��������ӓl3|�X3=���7E-���[������U $�'G l�#��k�M�&q���)�ާ�@�QǼIr�z:���-4������s� ��	&�p���Bg�K��#�3�eW���LLТ��{���� &I=\+e��&O��0��]W�҉������d�[�@4o�3D�+�1��
`.V��ӡ��ep���F�����ח��9������� ����:���g�Y�[.���������O���:<�y�yp#��M������$,���{�P$A��*FR�iƠ"�p� �M���M[���L�tP@o�Ci�6��E7=���,o:}������	�&'n��gX_|����X>_�e�H��{�*��s��۷m7�|�����I���o��s�L�/VP���dt�<H@Z"�(6Ԃ�0y�v��&Ʋ��\Դ$֒ly@1�ys�PnB������k0���3�p��`,��'��,�>۪�ל���&���m�⸓�YY+�{�{�[ �wޫ���q���b���~��Uf��+�m��\�����U�	��h��f9Μ�u(��S��>��g�r|�c��p��u�#��_<<�<D��0i�=n��=�����{M���p9�M�����+�)1ً�-�J"����m�UN6#�"O_�_\���	\���K
<1�K��E$�����E��VN�A��4˒:�[�<�t�f �f �fY��@VM+�U3����6�VM��N�^��,����}9ף���r��rd�_'�������������u0[��I��ؙ��� fF+�i9j�s 3W]�'O�$L�7���Z��f��W�)�'�Nn���XE-`>��Q
�b��(�C�N�&ǚ4e��S�l��dfekawL�KDRO��d�\[ˤd�%�(wd�k�>s�s���T�LIV�)CWZ�$4`����z0p����;u��W:=b� m�3V���i�h7�Qrc]�����n���:Ã����W���ao��/T��$M�w �[��f��� %&��
����"HXF Ty���
�`��X�vؾ��K-=\�?`�1q��ݻWᱲ��_}������]���g��R>�#RR��j��l#A�'���3�Z�Pą�,r���� N�����RSղ�q��~��WK}&�xVv�u ��ϟ�A��WJ�+��}��( ��Ɗ��I�"̀�x�P����m��0����G�"���@t�vp��d6c�$ShK?�`��f��e*^��^O�6���ueE{ u����9�"ir�@:�Kܷ������ns�_��K+����cՒ����x��2��C'�o`�>��g=��������[� �̬��ũii'��6��j��������!�v���=�{��=����e����wFt�,	Hzu��m�$�4�r[8-t�eY9Y6�r�[yA��Bw[4�V��,�^��4+�^Ld���R?���'D��9���F��rM��5�\��5��9�Z��IO/�`�4��6#G�Q�%��<9ҁ_$�$ o��,4C�S��7P`s�h3qJ��F��й���l�`:v��-�;\䃇�ln�7����3�[�Νd;@8D r��=.��M��.q�LL\�ٻ_�[΍��G�d_�2>1ɴ�n���K�ļ� �f�Ow2ػt몀���$�Vw葎�\ +�	�8Q�T��I:w1�����A��Z���������Y0V��Q���m��� �9pYo*ڲ��ᗶ��B�}J��9���^��������^��Kn>���ѣu�u��p��
���Z,���ɶE�������T:w�(�5Q-x�U֔��+pC	��5����e�%�DI�L/D1a�{i�n#j,1�+W�0��}7`dE�$�^Jr���ƽO�!��e|����J��p�ϝ;�lܸQ�Jb�����%���˛H"">�υqۃ���"��r��/o:�E.p��	�qS�ϝe��zr�aq����^ֱ��<0��f�~�?Ǳ�yu`� s�|N���������XJ[�ߙ[n�"�L��^�h3r>�����9�x]��L��@�VM�A�2�-�.^�B��H�K�3{�翹9�_ۿ�D����;}��J�].�+�o�,Sĝ�v�HF'������}��_7l����w�g	��k�\�,)A�A�� �I�SFf�)�'|ڲe£QQ��ԯ?T����Xo�����Qo��9�\r�ly}��U��OD��>�J �c�D�Oe�sQ)�8���H^��¦��iA�,W�4g �ۢ�j�-�egE�iUl"/P�%d�������]�?,Z-�0A�f݋E���SY��G�V��0���:v�D��;���d��%�׿���-`�%�6Uڏ3�*-`R���r���r|,�0��v;�p S �����7I]�0)ԫo_�#�A[ �rI�\#�3[�5-�o��}�(;��3G�q�d$Z��TQ
��L2�9��q4&�dd�������1{�"�A�b����i����7@��̕뛷�qY�܁5�c�w��ɗ�����ع��챐{��*}N���׾��m�������F��?2ȇ��7!�u$�p��2A&��+���(ET%��oQŠC�&-5����M]��ñ�@b����d�?���g�Z氐Uv�H\̌K�7c����/+d�'��f?����9>D�6{|�+�A�}�T�����(�cy%х�jj_�(�;е۩��\+�@khH�~.�;�OY�T`Z`(y?�"�G/`�Vv�ԇnN"�V��8�)m+�m>�X,$+���"m���f�h X��@4	K&��}8���uE��-S��0�?�fR��;LF���y�ƬwCH���s��y��"q�0F@'�	h�nw,�����/mI��5w��%�%����0�O>�����ܿV�nݮc�N�gddU�"�XMT�Ѧ��e����'-��6����m�J q� �f�d��r����)PtZ�z�����ɂ�6��Y�e�ge��@�¦ײYh�����o�VG��E��-9�"F�%�z���k�4//��>�8}_����L-q�Sߒ�6���p�cZ@"�!H�I��ѻ�8�qQ�8��)08Y`�Ijޢ����C}I��"�C��h]�#��LL2m�&޷__�y�#��*VDF��c㚛T��$�2�-`8\�I�ev�v�Է�Ң�l'i7�jfN�jƎo:T�-�u\r�_�Y丹G���N��Z�zf�m'`;��ϙg��p�t���l.Yn&M�a�Զ� �04G:�9�q[ +ݙ�:zn�u^�;��Bm[��_[߲����'�1�ף7$���<�4q	7����4�'w�0�Ü�p��k��7��r��yڰY�R�0t��� �=w��(p߬i���R�z��a��~ 'E�z��jN{�v�&�I>�V+J� ���l�Ȱ0�#@Wv�C ��ۚ�H� ����iZ�#��C�thGb�J^C:o,�$�u�Z���XVdU���J�w"���y�åM��Zg�)���1�.r OS:��>�l����y��)�lx�L�Z��~��'H���}�F�땸�=���լd��ٗ�2ıb�^�~�݌6s�>`Z��2�-Z�w���3Y�X��,��M����P����~���h������+��e7���d΁Cr̈́��������uWF�5����` ��*@	���� <i��?���j�N�ܥkw��zz��Դ�0g�o߹Y^����ٳ�Ҭ�,���e��n�B�;���)����������?�yi�Y@+�T0��l{G��O�e�~i�OĜuD�"�L;$i�r[6�M�e3�u�t�f 7zy�Y^��6���@��Mkɴr�#
�^ٶr�"�I9ח"
���yO���n
�=�)������J 3=G��`Rl��������&��I\%VG���0� s��If�'��m�B�e�h;u0}��;bT	`�f�14;�w�ց�~��z���fqq��oJ���hK�J��@L�SNo�58����/@�l�1c�IG��`"�-�*�;�L�^�͈>��`6��$�͘m�X��Y�s}��)�Mמ�L�m����g)���& =z��.�������L�|��.� $�ܐ5�K���&
�&�I�s,��(AO�(tʫ����x����1kK�I]M��y�s&����}X���>�Ql��QRh�[{�NҖ%����\���w����h�0�J���$��h>����,�m�&-�D�$N�7��>�wb[ �T`�?*2Ҥ&%ib ���f�{�>�w �e (��N�C��������`�m"�fk�6�O����P��+g����
�æ����dA�Q�r	d^������#��ڄ6M�6��+K��e��N�T"7`.^�L�u���Q7q��P�^SE�z���:�LJ�Q��q�oV����>|Vx��{��G�fH�����O̩��YY�.xt��_�]#�x���x���E��%�\RS�1�>����e�ާ[�x��|�lPֿ!�B^�N�ztRtZ���x����e�4��sk�,4��ݮs�U��4�L�n��� ӊ��9�2E��<���k�Y��V����?��_.����5������EN&w��,g�F�P�1��yr$�qH�0u��h�@^��ӱQ&�̑���&*`l�[�6�΀lo:)�%�V���P���G�PR�=+;[�q��nm���zڧ_�TC\�̻`����S?79%���M&^��i���%�`j�̼I�uN�e�����ɨ?�8�89@ 7�(�r=i5q-Z�VYY�$?D��čb�<ߍC^��DS�&Kn��(�>s�t�K�pY
��HD�~%��1���,�]a��'�5���;�_7�h���Zd}Ĩ��V�dH�[70Ğ�nw����<.r7pu, � ��$^����I$dkcu'��%�"븡��"g�(�{�gu�@q�S(���.r��ǎU��u+_{�5�֛oi|�7ǿ��e�N$	=��;`��G�g~W�U[���;U�<��f�34#�\������^����QS�a�e�JF"$i|'i��:� ����O��-�����\+��L�|���:v;�8V@{���,S�(�l����2.�$� h��Z�X1	�%�p��0��03��+��s9�����3�����/^�Iu$a���O��L��H\�r��O��)W��+�g���X���h�R-��Hj��c&L��9�T��[G\;�)A����չ�0�����g5%�+}6��P���nݖ:���g�3--cZZZVDVVַ>��6�s]��LF�����:������}�F�e�뎢�U�]��U��%�T�X:��k���sM�e���M/h"���<�tæۢ(F�kմ��u�[�2�ʴhz��K�-ǒ㟐c�=&�$��uͫV��gi�wxq��'?`��䤤��L��`�ɍ��"�/��᦭��Iɞ�ݺj�f	`��SK�����6���3��x�4=z��c� �s 3F��0�n�d?`
� �I))���[0)g4zL	`��ƥ=8Gރ0s���݀ټ��h�� <i�43{�B�˅f��,�a̔���&�N�zh�j/n�Ӧj1rk��o��f�{���fԘ�
������M�9�~��63}�LJ�ߔ��=k�&� *X��H'F#��{| �����Hl& U^9 ���LMN6ե�$!gӦM���v����pg���#�� &�j���m]��d����kF8�@��(��#��y��N\�� ���>&���Ϭ]�V��$?�E�)�Y�K��@#���MVx~~�3������NIY�$m�c}u��=��p�-�~�]w�hH��?VV��غU���H��a�����$E�`���(���>�X�t�ߞ�b���6��H�q��E��I>���c�:c���܅X2}�<$˺�'��_��g� �<�}恻{���J p�V>�,0ȹ&N���}4������.2�q��1��%r.F�Z)-�|��N���z9qj�%���8z�i��i�^HMO����%�y����p��A ��_<�����et�%�����K�	<.-C�7�6�vI��eݗ"b:dY%���8�e�¦N�U��:��j��>d�t�f �2���LdV4�%r���;���r��_կ_��А�kS�w�?�����< \���	�LNnU')!)'99egjj�����(@��Ḿm9·	�"�[ ��fK���h:v�I9��)x��;A�!�w����q[��\�`� �y��*�8S|�-32[IG�Cz ̾�d.R���<�c�l�,F�3�t����� �t|�fd!��̖:\$u=����L\���O�2L]�E�(玗}ڪ�;1���(�В?-#����J��&��_;�Y�D��!�J1_�vvpMk��L�专+U �]���U,{�}�råo�}?Xh�5��<Y��n��t�X*�^���'b�M�z�FOL0��8e�$M~�%7T����{�`hÝ>r�p3s�L�( WmEL&��ւYC:K�+�En���� ���6��XR�&����G��{c))s�����b�AN��w9�g���\�� ���[3�L`]-��<��\��L>o �Ϝ��{�G��%>w��t �~7jy��'b�!
��M��ׄ#&|}���͑�0n9a���A�}�l�'�1��}#��yX�z��G�#�I� Hl�w
��4E�cP��<�X� �#��Y�P`
O��B�������c�XEy��,�Y�.��o��
�jnh�H�ƭV�����_��%aB$Jr��{������|� �2s]��r�����h��
��%NL��IS͈�㵏'i�c�.&+����SR3^HIM����	�L�[��ze�c��d�?��O#[���b��;�|��v�ѧ(_�������Eef���¦�lz��4�E�2�A��ע	hV�>d�dͬhzaӂd �t/7h��ԩ[�d���_j�p��^�޸?���[�{�8}�S �L�L�L���8A �$�\A�*@T�l�q��;v�_
0)�>Tn
�:t4q�M0�0{� s�s��*劜,r ��Io�!p۽`1J�=V�\�� &Y�ݻ�L�s��.{̖�I f�R�9pP�^#V��]H�0[�6��*��O S-��k�[�o 3%-Ua*o�d`:n1:��l�^`(��_	�rC�>#_��A���6�G��2E��n��vI���D���X��
�:#�hٞNut@���  1{@d��C��8@�Cj.��Cˊb0���a�#���t��G�J`��9\>��S��g�Q�������=,$ǠT�� ^��G�Cҋ��]ׅL�ˎD,&�K�(�P�#�	�b�E\e�ʳ�L���)���n�pwci���P�)	�<0̛7O��|�ī��t��Q�v��	���I,��Q��xh ��5�E���o�£��Ů��+��2q�{����K�F�7s���?@���wT��s�2�L��0ȅ����0���c�/eO��P��`���4��D+t��f��k��{��cz�o���h���L �2�f���R�S��X.�O�fFO���,�J=�~�Ѡ0�^HJI�! fe'ܲW��J����74F˼�М-��d�"Y�E�/ʜD!,��ȶ�3"?`ڹۢ�M/d�����MkѴ�L/h��>w[4+�6��Y`z!��(]��
\~հa��u�?wc��S���a�Ę��q�����29���Ly
<�,��Rn��{�Vo�2@['��� ���~��p�c��yĈ�j��]�0�� L�����]z�Tp�k'ǹ�
`0�2}2�H�̹���e� �������� �1s,�M�@�`CL'u+)��8��}�>�0p	w��YA9�Es٧���́Z&i��aZ���-�L �QzKg˸�6�j��9�)�Q�d�"�����A@H����)��R��j�,$ڄ��o�/��� ��6�e�v�1=��%ﱼۜ:y˵�:�q,ϔeb$�k�	ޮ7^w��@�My�&O�#F_"�G�	�a�8H��4����$ ��3q��
1zX�b�*�E��Qz���U+#����%�p,��X	�^����78��d�ۺ� ��o�]���G���}ypw�Ǵ�˸�MK/�(�y�2]_�ľ�,�|?�Pb����^���X���:���\$a��Y&Y�ڜ��y������U`�8X�#ßc�@nFmڴ5S���og�Y��yH�>� � h��Mrl���M��;�=N�F� !6�:��Y� ���
�+<�� ����S�����L�s(�F��:�1\�o����t��[^�,Y�٬\%��b�?�{/yH�~o���r����\���B&�ۊ�3�?�s$��lu�F��$�>^��)׽G/M %5%5�xrJ�f�`ډ��VX9�p��ġ�������D$5���K�d�S�q����2R����+��?3�-�n��6������MkѴn��I��+�^�t�"K�-�^�~�S�58�<tw��ѫGh��zf��|��o���ҘW�L����>��d3!))'19ygrJ�Ѥ�4��{	��� ��d���� 2��X� L��6H������!6֤�8D���*�Ab&qA����v3I�)&�y�@�Ev�����;���$ `r���qA f/�J��x�^��h��-�[ٮ�&-��#"V��v�;�+=VΝݦ�Z��5j�9�A>k+L�g��f&)%����K:��
��������pf�� L��χ�y��9.��@[��Yz�/(�a�n�����:�g��J�����͋�Qd�o�~�k�nj�憷|��r�vF���ȷ7�u�nW&��5�,p������kF�iƌ��0����Qi ��s��vF���2c��	�a�F�I�MF����p}��Cr��di����o��O?��y-�	x%���:��N�e;�������\X箃hֹ�8N��O�x/����mذA���g�o��͚t����k[\�d��J'a���Xv���O��|�a�#�'}�F��۪֭e��Κ��C�}�q�� H2y�!TÁL2�K&�<-_�g�4v���\����L\�(���9s��ƙ��9ЪH�)	>�I	!��gfH;��e�H���e9q�K}:w��r���3X��ȃvo3j�8���
�z硙>�e�=��>����{˛2Ռ�&�h���Ǜ�#F�} W]�|�T2i��-��� f�$`�5���+�_ ^�� �YM�1Q@����
@N��B�;E��L��d����"Fz �D2-hڹ4-lZ�fy1�eY4�.s/d��n�t��}�f�5l�H���Lxh�χ�i����ǎ�����&#��MS�A���'�/�xf�ӟ-nd���jc>��|���������l����=�~Q��?7�~�3�w1�RS� f� f|RBN��ĝ��)G��2׹K��!
����O��zk�
@��_�}���uK&q2@^�܌�6kf�22e]_V�$��ƕ��16.N���:w�m��w G�F:��I�i�Tx:v�l��*P)�iC�&�;��-}$7�����79�YG�O�����Yj�"7,�pm�29v�N�����Q�|��֣�-��3͔��1��k\_| �Vٙ�k�"�"W��A�
`�A�`W�r@]�1�m���uo����S�+n��Ijѥh=�3�fAm��r����{$�7z����g�����V���6��CI�p,Z�Ӧ)���C�4c[c�d_ॢ2En�"�q�9F��r�֭S�	�*����" �+&�s@�?p�;x���杷��[9�w�˂I����K�k�I9!>3����`�d+@�Ϙ��\�N�����g��b�O>����{�
�]�j�~��5 �Xs9���e��a΃�>>���l�-�Q��q�:u�ᡑ��nc&N����U�:)���0�ɂ(�i]� ��dZ��x&Mђh�7oӶ�<ܖ����zU���)�4�L�����)��|!�:ړ̄��{���<��4�̖υ2C�V�"��ƬX����r�j�F�V���������{���C�R
j���F�k+%i�W����~���&��9.�Q�ƛcƙa�ƚ��͠���AB( �g���EՓ��}�Y�t���/��:2��pL�����b��Ge�S�/��SYG��"Y_d�A�¦ۢ��@�@	Ae���Mk��Z4�gV�nMD�e��d�F�e\�Y:%��O������Q����h���>����C_>�N�i'�vH;�N���wz��4/�hN�3��jq�˧���řo�hV|���뽿�}���������0�sZ$���21�hBB�Z�p?w��Q`q�!���A
\ Y��]�K71d�����d}o����MlczF��1��i�� Ӽo?�*�4J,`�Ln��V�XE���#��峛��.�i��j�� !���`��y�m�,�']:~k�似2_��m&��JA	7y�>���ֳ���5�i������S�]ntꏟ<ٌ�8I��'i��Б�L{��y/t�}���8E�r�*���+%7���l󃞯���i{���c�ڟ����\�i�q�׮�'��L ��K��&�o|&�(pӣ���[�k-;;zǅ�=�NJ�09�xٙ�4��� �
�>�FF��uN�&q�X?�,��L@w8e{(��{�2<XO�p~o�~_��M����|�@ Eթ�H)%V�8�*��}�*�ȂQ��.��g��q��yz�8Q�@��s��j�u���7�'<��L�߭��j�ܾ]3�	3 ��%#��|G����:rc!N�$�2Y� NU � H����a=��{VVk�=~;+nqR��1n�bʒQ Wy��q�oَ5�)QD��v:	��iG޲�P�<X�<N���@��MQѿ�&N�*wS�xٟ~�����d�w@?�5���G*p�v�@�K�V�u�@���f���`׻O_Ӧ]{y��U6�ƉS���l��,���u�����0���,B�ʜ��!�#����}����]{���ޥ�瘔�r<!9������	))��Ʉ���_��H��@c]�tQ?���<Ap> zS��l;"�\D̦ߪ�N�n�t���Mo�fe,�偦۲�L�n�.M?\���:����>+�ܾ8�|�構�ir�����W��?Řm��7�L���_+|%���b�(|�����v�y�N�o���om/.>�M��J?8��̑f��i͋SY���u���rZ�l�3�e�Q�}�HLb����_!�B��� 7x�tl*@�<V;�����Y.G`�4�H��cJj��ڵ�X�
p�M��yi�K�UT�� -�Ա�����$Z��6��ZB����- ����a%32��q{#����6�I%�����Nk��q��H��8o�.��<M*׈�_ �mۡ��3D��#D�G�� ��q�P+�с f���0��hS����V�z��]�ge��ש|ǐ��fiyS����;���z�7N��ϊ��Ē��mw�l�'�pr^q�_-7�)r0�C,��B"�>��Gl��%F�m$��	�،e@d�f�*��pw?p��z.�k��L�e�j�|ƥ\^Y���̧�|R�� /�X�H"֓����p	����+u�sn���g���zJ��	 &��K����f�L�`⢒N�ϙ�G�,�.���	/X�`�Y!�+F"��$��7	���#�1M�;��w"ˬ�5@i�9Y�������۲0�w�}�)K�#�L��$�Q2��;�v�y۝�vY��#��<^�Ǎo���=��:D�a+�N<=��He *��!���K ���/hK�%�`jz�IJI҇d��
÷Q��D���&ijϮ�t���?K����1��������$_R]�"y��ީ8BI<[���zb�Im� ���������_:%�2�r�eb�	I�3�y���?��
��
$�`�/@* ɈD���\�w��%�^���"Ja�,�n׹ךYhzc4��	dzA���L7hZk��L/hZ+�ے	`֫�ES���pӽc��7�}��K��(������:�R��^�{���oξ�̜z=Ҝ�WP񉗂�
^�)*|�]���F��lYљc�z�H����ԑ}�o-~�۟}��)��ryL|L���f9�[4�ټE��8-�� պMk��z+\�t0)��B@�I��22��\��3 �e0+���bS�K,��XvH.�X�؆�K'�f42����r�IMu`0J S�r��S��Ʈ�zjlc�����@�+������ 0m�xF�,���,�b����7/Ŋ���l�b���4��s�C���k��M�Ib.b�	@7>�Ĕ�Fƥl3 $� ��m *$*�90� ��M��c��X=m�Y�� �'� r�y�k�)�e��#:M�. �T��M�gW�hS� ��k��+$I:��H����!��
��0Ɉ&��C��B���<_�<+�Fٝ�e\� "�v�l�ԩ:�Ӂ ��j�~�:�b ����ڽ{�fuW�\ˮ]��C=�V���_�a�ƍj�M��'%���/��6���l)�0=����hJXj��e��V.�07mب��lp�1ׯ_��o���W�ԇ���d?dZw��u������58K�(��Z�&�5�����W99�cnܼE��`:�m�Vs��U��H_�T��f��ѯ�ëK�C�q-��Ƀ.Ɇ$2���*�W�f��F�HxD E�i��c��䁞>��)Ӧ�����o۬�,�-'�~�m[͚�Lޤir�=LFF��K��ys�	J�GR$�ue�{F�Va���K���W9����xХ+�]�^ �3Ї��0S�G�)::����Ժ)��'�� Q���%�A�c�5u7��"�R��4�r�{A�<�9�	d�e�t�f ��u�[�t���M/h֗~�~}b2��+�ީ�ۛ���������T�f��ovybo��'�������1�6f_c�	��~g݁>�m̉e���oN���3���9�/���p�����_����f͚�4�m�3&.�hL�t�r��(xN,c�s;��;�%���&r���pi��Xx�x���F�h�	�ؾ}'A�ͱ�Y yd{nX:�sgi <�խ+� q�@��Li� ������8=���#9����:-ز>��=w�>��vg$�={i;:3,�\#�q�7����VZʉ�"�ڸ�n�o� 6.u,�7�S:�� e���eA�
0}�����|G
��r̤�3���9�%�'_�  sҔi�� &�C\�m��5�.q��	<�B���L@�'�O@����|�NX��p�S���&�H%q�����rE$�����^�p�I�v�@)��[�n��$�\� VO��Tܽ����P��1����4Vq� �O�f$7cpB�b�N�c}4y#���\��R0��"�gR�D3u�ds��e� k2���$��|^�������L�8Qa><4T��XH�ղ1s,�"7`2�,CZP�>�R��2�b2�̆�I�!����X������(0a�#�T�ѥd��X9�Sy�uC��~���x������x���S�.:��3"Yp��y�A�lo��9b��s�N6���g�W�l׮�IKk�^n�%������"�3�?�_�G��b���o�~Ѯ]G��I%ƽeR��		��h ��楗^Z��K.��ӟ�4X@2C�r��W�p��."1� �Y7dV4Y5ݠȢ�L+�2�.s/hZ�tC��A}SO �A�F�M����ܮ�m+�>�j�fŧ��.>:���O��<�yܙ���5��s�1�&�� c>�d�YƼ�d̻�Ƽa��8c>�h
���u�>��~�����:�=$���������^L �.򈘘:M�6�i�$f����h�h@���!.O��S�n
ydeZ@#m�ҵi�N;�zh@��Ш&ҙ
Ҏ�l���cm�x����xM4n��杻vӺ�X��z✑�Qz���iӭ{/?�6�]�`�ӧ#��i��j�,V��b+IZ��x��Xy/X9��}c�%��� �s��~u�kJ'��E���I�"��[8��f��v�A�m>ht/��R�9���д*},{=����9ǲ˴u Pft"�0H�ۋ��%6�Q8�M�����o# �̛4Enpm.��fڭK�V����d����OWk#nt`�!�Y�$�nfr�f���5�p�ԩ?�����?$�H�v��䠁���Ν:i=M ��#]��@IBLd��A�W@���A�I��	Ԓ��&��ɲ���'��*�S�����u�cI�R�[�snڸQ�Ur�Ī��}XoI&Z*�,��⚟1c�f��N纟{�Y��O���q��{�.xJ�(U�:�~}�L�F��`��o�B"���3��3V��M$�P�h��׷n�d,^� H�((�5Q5����d���%w?�k]����K����������d}�uzh\���#�҉w�|54w���sո�ъ��t��_���G�E��~�T�,{��_�q���n�1�i�LBJ�i���<ȿ���0=!�"`���1Z��_
H�E�2L౭��0y�B�=.b�����u�[ش�YY�&��M�뼲�nK�2�ܐ�M̺��4h�識���۷�27/9�=��..�{��a�}�o����k��O^1�+��J�ǘSOJ�Řcs(�~� f�1{�N�9�j��ך(~7����;�����K-|���ůt��y�3���I3"�NttӜ��蝢�����@�c��`1t:: ׎�Ua�d���m��$ �X#�#0i�zb)��<�"�M�]$ ���s>:0ίn��TQ�1<R:g�F�؉����׈%6"*�D
�b��R��8v�ٶ��Ҥ��B�I����C��5�?�����x���dn�����`:q���YN��ys�ܐi�MNaO^�T
(�\�? ��'N���<�9�8�L�4U- ��<�2��o# �$!�f��L)���&���r&.�r?��ļ<श"�^(`���QT�� M`� ,� '���^@1@�����S��	w<�0S�LQHH�VO@�ښXJ�R:�v;v�Pw4��R���f(Y��OY^�zE��0� V�RE?[`�Z�X]L����C���rS!k�$.{��X7�G��r�ࡁNXp�T�K1�ي �Ź�۱)�/T��x�Y}+%�6*PZ����uf���
@c��L��A����R��μQP�Z4yx�K� W?�ko�△���}}���l��Q�C�M6*9C����LJNU ���ྦʈ~�-�;�Ȝeڸ�;�,�A�m%��5�H��W�E�E�<�I��W�9�V6�B#s,�;(���B�OyJ�����n��6��ϧ��ۚi!��YխC�Lq��uׯ�/8$趸��۶m��=�׾��Ӟ�?����;���gVJ��/��EE���>���o^}�̑;_>��̗���J�i��x5v_��M�����D�E��ts��'�J]w����������j��*c�\j��pI#0#�DDG�DDG파�:�P&7C 
WKfV��^ 3����)���$�7t��v���m���rS�-0Gg�qH��ɔ�F�-2
ב�΁�d�Xm;�k��"����ұxN�s��
�a��m�V��,F���}/r�0�M\��bJk���Q
�D!�R�)X7�����s}%�'l�)���͚�E����h��~+�9<�Y�c��M��`�^_F[��׻��}J���*�("��j�����'2�&��0��9��v����	`�%kX��(�]2������s1�X)���-��=��q�lp��.���B�Ue&�?�����ڈe�z�X�Hp᜸v�^\�dnc�|��ԒD��9z��*�60�����e� .�Q��|饗4Β�o�Y�ZK*np`�B�CV�4��5�"�G�|�%$Uf������������]�w����ٳ5C��Nn,@!�O��I-L,�@(�H�a�H����ϛ)�<���1�*9�J^7j�d������m��o�B��-�'�C�[X1q�����Yd�S�h�j�Z��o�2CT��A�N]�EW�٬{.�-��Joޢ�>�m@T龤lQ����ׄ㤷j��<�F�C}hx�	3AXLC�cQ�*X��1B����@��z����n���||V~��6�W�zSM|b��u���{0+;1�������U�2\�E�"W�����
`��~��9���L@�9r��hr�{!�2�@e�fZ��2k�T�V��jhѨ����ѭ;4��9�W?����}�������->{�[��/�������^�s��}N��W�����|�ǐ·������½�-ؓ���כ�0�Ę�M̩ף�x���o�]T���g����gk�����q���X�0â#r"�"v
8 
� �<E�K�"0��thX�pt������=i'0���б��:�q<:D�ɹq��� ��Ģ��
��r< �vXEqExN[���Z 0$,L-��n�ܤ���:.�%�I3%�v`����ԓ�����p����q�
�rn����ڧG��y/jh%�sҔ��V&��?0�>{�3b�H�"�A	`N��|����)Ƽ�[ɹ�߬�I�Y�X�H�`�FH�u�o�n�#!�R7�e���� �=O��[oi�Fj;�>'	i����gF`o� Eǉ9\�z�ٰ~����CdhJ@�����Z~���q���}�6���[���2>��)S�XiK�6�O��װ�y�m�/��=�x��&/`��P�dy�X-�ɐ���}b�廻An �峠&&��m�������y<��C�Y̙5K��d�x�G��0G`��o�"L��@P�QtJ4o��%� �5k2W�B�#��o1�W�@��L˟���W֬UG ���f�z��z���7P��_�a�O�+�yٲ�>x7	6u��5�k�2�jԔ���V�m�Lu����e�jX�j�4��&4c VL��@�Q�fG�g+�����s |�-�T�����^���{���LII�f�E�<��������& �Д9�@,W�6��-�B����E���(6�,��M��<PI#��\�N�ڦ^��C��ؗ�`Ø�f�n���Z��8��
����0�O'�ι���c�9���?������ć3�\x`��O�?7���3;�z��w��=�F֮{R?8�V\�y+��Ҹ��f��z;���t[|r�Ȝ3/I����n����m^�a9��;��P��1Z�\�9�$�
�Xq%���N�L�ҡ�Tc�ot$װ��#F�����΄d�W�Qj��*
�1�Y�jEP�va�a�&C<95M��\c�S��8$D��7n+:%�x�DF5�X�y��ܼ���N\�@5�P"O�!a�X˹5��3R����Q�¥S�Ɗ2���ǎ1�I`�d�@��فOw����, :�%.r߲O�6Gv[ɱ��k�R���D;�L-��Q�![���0��� L\��=d��X(��,�:�,lZ��=@
�T����j��$��.�M�s��!#����<��DY����{�쩮ug]��d{�2���q�q)3BѸq��rIf��5k4{�c�iu���$�e��X�i&/`yԯ�'!�䪉ŀ���K�S<q����0��2�<X2��X&�}Պf֌��]���"�q������dHA�~{���0�8Z$Z�D{KWP̀�E %�CT? 9h�Y�d�ְ$9$4\�V�:���v�Ҫ��<y-���<"R�[0�m��#�x郀-����
D�0U�&\�ZUS�z�����UU}:w���In洯S����aSO�Vb���Uf����Фd*��C�����`2yjz+u���6���?a�#V�
\����-(�8;�k��n=)zC��y���g��mn����&�A�l
h�Ȍ�Y��V�y&�z����l�3%�gqNލ�+1��|� �����'���_|�N���������&����̾>o�I**z+ڜ|-���7�>/x��'�{�?y���O}��s�4(>r7uK�w&���&L����G�C�"+nf��X-��t<��>����ȓ-���ΠN&	C�		�j}��mx���y8/�k�t,��
��""&P��h�q�F ��tJ���5fi��6
��Bk��x�l���v\�}/��{Z㤔T�UbK� �Ar����y?@3��
W0���N91A}rr������M�ͧ��`b��2}���(G����� S�+`P����E�-�nt~��Y������oԂH�$V�{�WK�P��=3��N���ԃT�k֩d��(�$�^�DD�6S�b�X?x��9YX�PzY���_��~^��e� L
����R��Ě

(SK,��GyX��w�P+-�d�Ӗ0�|w��,:�h��+/`�$�9��+,�tb:������|����56U�VS+a�Z��Y�;+�M���p�#�}���PǗH������):pY��j�$7�rS$n֨d�jr��L��Aҧ���� �s;e���@�����:�f�¶��u ��x<���"Δ�&��O$%%�~zF||R�E����O��X�� �|�����e9O�r��QY�O�?�����������,����h�L�7T�b�.�����R��ɫ^�̫��ؖИg�N�_�ol��1S�1��u9!�5���O��������>|G�ɃsN���S���ġ��e�[A�൸�3���)��߽�{�M-x�o����j�V����������[�jU�i�f9���;�C��Q��?v��&�⇵���!:Q�y�FK�xuq ��8�����c:@�S(� 8�h8�ŭ��ΈH�|h�!@H�",��fr� 9��$F7��k��b��t��r�A��
��N;{�������Vk��'���s�T6j���{��*2Z�"���80�t�rӐ�P�5��x��a�W��JÛ_em� ���+� �����/��싽\���	�0Lg;`�I;v�D�yz�=H\�č�k�Ēeӂ���eT`~�D΅5W:�a]$��$���V%��{���,u,�,�{�]�޾}���b%I��M;�9	5$�|����Z[��ϼ�<Xa������p ����D�-�2J� ��&uB�/J{��RJ$(�X�9O��XS^� &'�"�,Oi�􊶎LU�}��L�r���Pi����:#��@�;�F�+
tke#�L2��;ס�8��;��#��#���ʪr��������m.�{�m\k����a�Z��m�{ĥ�K0Y�RL�ɶ�}�>�~�����R��D�]�VB�D'�ǽ�".?.!.*6����;��⑤�B@�F�h��$���% �G��,�!�m�2-hz-���hVT����M7��l6�Z�L���<S'��Y�Qh��G��=t�m��L<ھ�_��:'�|'��k����2����}��ҳ��2�Uc��Ř���n�9���9�f���}-��x-���7�g�c��w��/�3���,��ʹ�����#����yJެ��8C�\���J���;������k&x�~N��/����s�U�)@FI\,��p���;�.���O�Z)EA�:c��N;kI�6�|V�L����hS����B���N�K�U�M{�CC�}�r���w�x�B��#P�ۉ��&��Z�PE,���Q�^c��^'"ó[���	�������|�h�k��H�����rz�;�\bA0��.�?Cэ?��8���`~W�9{~���/
��;�w深���M�fM��'��?q��l(�Ι��;��" N�3���f����+W�T79q����ev֬Y��`O�u0������b�\$ He&Z��c�.���Ϟ�O�1[�9���6�647T��T�r�����@[5S�Fu���8}F��˒�c�����<H��A�V�ھsy�9w`��Z���[��%���$���,���c����D�0�]v���k���}Hw�Zl}�Z�Lx�0:4�i�MӘ��4m�tb\�&����W�nq��v�T`���׉B&;	DN�$)������@�ۚ�v�WƢ�u���i~�@�u7�`�v���j��rsH��G�Z�4�̩�̱���D'=| &m��͏{��#g\�~�wSJ�}�n**�?����1�G<hL��+ͩ�sͩ�mΚ��8�M�kQo�������KO��3��g�}�+�k3�q��2����PT�&G (��B	*ļ`�LNI�?;�JCn�
o�%����[&&)�Q��:��>zSS���	��oY��-��Ab�Ī�ő����t�<k8'�C�kZ�UԹ�4� iS�a9?�Vy/�yq�X&�F�y���4l$�G�-�l]�<%�>���X��֗��y�Z�R��>��L>�s: ��t���cƍ��> �2��d�mH�O�R^�]��0��'����o�9�g�0�,]jf̚iF����"o��I�)̹r3^��8k���V	`��\,��L sR)��ɲ�n{0����|�dy�1�ՑxQjn"Mt���k�H))5x� 3b�p��|͇��Xi�ڻW�/'��]�`
���[�J��G���B$�ŲT6���C�s�i3瘩�Se>%��45_�M���4��n�rc� �f�ښQp[��i���Dl'F�������C=�=����L�2�"}�S���}����d�XشPZl�����eT�袨�O��Fo�e����$F��8}ӏ
�p�"��ES�r� �z��}�G����F�2��L�Ve�ͽ�L7h�M@�o�__|�76���������]'��뛰��_Տ9u�N���#?=P/���-�%��| �K�)�k|���R��0}������ߧ���2G_h~St��oΞx��3���Ʃ&�P�'��/��<�j�����/ڗu���O~0|��'�~ozp�����޽������f�mH=ݴ�a ��t�@T�@��8e�I��+C�@YCǒ�X�}�1������q<�1�8L2�:����t����S ӱ�6�LA�?�X8r<έ�(�.m��o"����mPO�ˍp����5Lp��Aau����	��RC�XN�9��-�D��DA*��0�fRs���3��>������X�������2T
B�:�y��e�׿���S�M3C�3=��ع�i��"�� �-n��,5��&*Ȑ���@�x� ۀ�`~���wN\w�L�X���s�dT<	̑<x��[GS�<p�J���J�䘌 t��A��3ϘI�2E��T"����>�d$�Ys��;Y��r~��#,�����3ͤi3�$�O�?i��*�0o�z��5���>-��̺���Ai��F����-�ΦSWS�Mಁ<(ci$γݰ(R�,�v��D�M�8q�A���c�����[���˶��:�<i��g�Ð44@�S�x�2�I�1�g��j5=*&*.&&�6��Q�@�5j\*�_	`^+
��$w�嗯�����G0�M/dr��4���[����@���ɚ7��A�M5v,i9wr��g:��u��k?o��_����:Z+���*��Ԋx�`h܃c�Hn��XZ��C	Y�s� .h2�G������ƜU\T�T����+�O}����KSN�|��7;.(x��}����q���B�i�9�V�9�N�+ş���Gs�~���W���w����fV���R��v	`~N�PC���P*�X�2 ���~�<:vM���� EvVI�� �X�a}�`��QG�9���#��7@��W_C-N\�t��-�0�����
��h9o��u�=��E7yS�[� �/A�Z2�k���'d�:Q 8d����6�t�n�h�z����rE=z�4y�&�S��B�r���v9
�nˤ��輾��?`.\���M�hb����L���?P��˟=Go� �L��aEb��q�L��.��U
@"d�R�m�0/N%S �����K�O�'����1>5@�˷M���k���!�t��c���z�Z:���;�e�����G���)�~W����4m�l�f���
��'O��3F���Q�K����o��Ƣ*ժ	������ZuY�^��F�ZEu(�%�xQ�Xa٬�
�"�C�%0<Z�Ƚ�d�L+�%��(Z��k��������-���1�UN��j�������������E5m�-*6���������$�xM��p�l���2_'ˏ��Y��Q��en��^�ye�2�ȼ�o����ox��M5g<V3<�8&��鼙�N.^����٫��q��m/�Ed��,>P+������l���H��GR�7;Թ��+��ߍ1�~a���*�>и���O��q���0�72�`o��{�g��d��GO�^tjOtQ��N�7��̧��(�(����U�Z�;����/KOO����=955uo�f1'L=G 
77�H��,�(��F�	`�#�q(nr����G�%�/*8֧�[=�Q�ɀ�ʱ��	9 �8f,��$�$��
��+�6ں��\#��-�wJ#՗6u�֖�����qx�c�Y��Z�Ȝ�tr��ss\��,Y��/�a�-���/�����J���k��uhoF��I2+W�2�W������ʐn��]��^J�6��ZW��m L�x���:c$w��[��M�Z��q�ǌ/7�Yzs��l~��2Ǎ�� ��"W�tÆO
�l�׸�˫�i��e�^��y�������c�c�d��N;��A77�mne�Q�������n����k���>��<��Z���^�ڦ�|�����]�̴�4��;�L�1���>k���T9��V��*'�1y���H���0���j׭{솛n8 `�Y�5>�Z��K5>���F�Z�լU���u��,(�⡘��Qjf�TRKS�yT ��`i�^��%��5һ��E�g�6 &��ó�)�g���t��yi��D��-����V [~K�{9��7�=$��S��S��M�l�L 3%4.���[�����t��3�p{� %1�cDk����_~�!�W���4���֚�g�?]sͧ7������W���:����������Ǟ�Y��?�<���ś�6g��7Ǜ���j��CU��l�����{�uu���Ǘ����=\�dL�O��xY�E?����^|tÕ���v�ݡ)�ou�y����N�����#����O;��OzS�n��N~�7䛃����eWsߡ�3'\	��233��+`�Z��3#���"@F#��MgD��0�?��(�p[��L�,�M��&86��
�q^u/�y9&@���ȵ��S�ktJ��\RH:='�G�D�X 2Xc|H�i*�$Q��I�>-��Y�n]=���8��^�,w�Di�u���[��3�&��rА�:l�"`.]��̚3ی=���;@�Gvf���u������hrs�6Rw�@��q�/�w<}��_�$>���a�q��Ϛ9S��Dsf��d�k֑)N]PDzJQ�驧�ҡ2iӡ}{��2�fcBZ�w���-`J&��3i�t3%�9�y�ʛ2Ռ�8ٌV��3#ƌW�9f�>jLq�CN��n�ApX�3�j׾�v�:w֨Uk� ڝV�wV�Uk{��u�תS�n���0����9��ٺ��ME娤�]G���{��L��z����u���E�s�v�:������<����/�^C#�p*
;�jTT�y�QQqA͚��wk�8����p� �M�!�mE��554d��e�5�mѴ��M�.�<��?���k���7�t�̠�U[D���������yˮ?s����'
��۟x֜�2�d�4��I�h�s�a��5I��`J��G�j�ʹ0{�\j�n�έ��U���v������7��ַ���ȉW���u���Ģ�73�N�����[|��g���|��of���L�ftt�O̬���i��'�o&@V �ȩ �' *D@X$Y��xz%�x�+&IA�/��ML ���2@N�M�p�`Ci#��D���7{L2�3���S��|� ��i0%VTkNʹy��/!�7PW>��c�#�D��'�ٔN��v�zǥ�;a�r���k&�e!�^#s:\�� x+,��\;�l��gT�0���Lo��W��~�e?���>��#_��@��u�^'3����Z�[F73�u�/6��G�4���ӱ݉�lӶ���%놏�7��r3�&?q�rE���v s�@�hW\�n���� ��ᓅ�l���0�-����k����jús,�.�d�	��k9.n�aR�Ȋe��@(�Iqu���͸�c�}Fz���9.	>��Yv�&��������'��M�<�5~�d3fB����cͰQcL��Qf�h���1�sG��������v�4'!)ePLLL���u�V�Z�*U��`^�f���jժӭf�:}�&�جY�λ5k�-���Z���K�-�,��l�S�����~���>�r �t�u�:�	�vDH�F�^#�Z���G�k�IMP$�&�A���_�=��ҟ�E����ϡ��!!'BBB��(�)���|����c"F�]v���9"\�{*`��Z3-dZ�dn!��e�t�k�y�v�����!93�b�~+;�ڳ���/*.>���SƼ��1�n5E}��¨s�vd��~���q��������߰�O�s�\�;�w6I_yY��+�R�H�w�?�N��'��]S�Z�?N��y��Xs��f_�}������?}���N�D��?�P���ѿ�hˏ��k�^'�K}Y�S4_mڬ�'\{.�h�&$,��Ò蔃`\���H`��<Pc���IgP,:-O���#"���$هLo /J +�<���wE�xȞ[t6"*�+9����4l�_�f��Z�k�-�!�QQ�z�O7h�� K&9�	�yd�&���� �ɐ��O�_�װ���Cr� G��{�x�9�trg�7j��.�sD������%�c�+f�n]��S�rEX�]> }�oG�6eB#��.0�:�^��䦛�;��l'�٣W�3|��7�L�;7�q'�+ڔ%��X���a�2��1���O�9YmX0���|qy����w9#?_G/��%#8P�3��ypY�f�Y�v���%�E���Ӵ��W+5�ܖK�Kd3))����ߌ?A��!�/L�ͨ��,�*�A�o|�0����]0f���'M�_>-V��3�5��ɹ�Y�f�רQ��믿���ի�n�Y󆚢�rw�Q�vJ͚��kԪ�l�����QS��f#�M��ү O�H��:@�� L�B̹6F,�_���w��-��~���U�M�2���N�|��ƍw��6��=�Ü.�Af�W\1Z`r�������@�?��B�M;��L��"���|�^�z+���;:��tE��}6p���~�qǳ�N=P\T���S������
�}�/���s,���G���~����ၚ�|�,}�Acz_}[�G����_^-��NK��3����|���77>�霶o^pbO�K'^�:m�2fc�3�>�Wp���;�~~����{��ꍄ��5[�.��ܹ��222�	dv�\,O�����j�,f{ll�+�_V@%nb@+,2�TpX�!Y���#��iK]�fq�M��^�g��4="��~bR��q-�	�	�j�5��+Z@�9V�А���e��VL��,�hwdT���+.�
�"P�%@h��>���l�(������"��8��T���TL����4�yP�g� �-��?*��gi�0����e���l{_�wX�S�W|�N�N�s��E��E�M���a#�7u�p����%��I��-�A���6�N^������׶d^�o�y�����=N�K\�^�d�n�{�A9C�M>Zn����[JaU`sp�M�`�AL@�^��~�1nye �;�Y��jc'��۾�c�O[;���4��9c��gNLu�ز�<����M�t�q���'#�!0�v颮�;�n5O<�y�����O?m��>��RF$�pl+�w�~������hz���XG�Ņm���h$r�� ce4t�H3$w�<4�/~�s����f�Б�G���=qz��y��nٱ�w{�카W�^��m��I������^��j�k=V�z�c�^�q��K���:�x��w��u��Ze��9��.[�,&�I>�O�k(��P͹t�l#������:���B��fj�����nШ���4j4�Q�Fa���b��z�L �/���m&��V\�C �d" �¦Nk������Y�:uv=f̘F���9��&/�ғ{�V;{�X���?�w��o�>th@�?v��j��!_�_v���}'�{����~Z��O�D=$���������;�|����7��[�!��I��ܳ�Rc����WO�t�ŝ�͹���v棖��6�S���)|�����׼U\�����O7�����ů��w���S�����̴�����M�f����OJJZ����	\�X�""
0��{X�)4,�ΐ���`y޴o����LKO?�E��E��32�Ƿl�OQ�L'�Q�k�a9�?L�����.ˏ��}2/��*mO5�m�j\���1��=£�2BB��h��{�'0d�G����Pppئ�����_mҸ8H��T���f��;b�7�%�٦QH�ɍ�=ްQ�c�z����"9�!��a!ۃ��
l�u�1O�;�� K����M��\��,'�\ -_I��H���S_�6�]'��:��%m/m���V����׶d^��Ｒ�xQ s��|3|�HuA�.]��~�\�)c��7��{5r�8�&4H 3�DX�,.�3�O[;���4��� ^�j���LrϚU��믿��h���i� �t�����}fL�n��q�y��͎;4*��#{�1W �mdD����g��@�ٲeKӵ{w3$g�Z���Z"J�/HI�b��o~��!"gy�h���f���\_3n´I�&E.ٺ��n��	جZ�jm����j<R�Z�cU�_5��O�J��C74Z�w &�x��:U�}K�}ޒ���K,���ge�F�~Ȭ]������W�A�mu6ڠq�H��{��-��}"6�W��	T6�l/@���G�u��M7d�,_{�E�pv@X呴���={�^�z�/�� 2KY��,ް�������[���ܛ�9�x��}�߬��Ŵy�:���N̩�6�H�fgG&<ھ�+G��z����cC�z����}/��帗�?��ѻן:��؜^f̧]���CL��u�ٷ��b�t�;̙c<���E��lZ���`��9�����Bfrr�11�ĥ���]�v�RRRz
x�h|]@豈�i���6�������_��8{�QP�a,�@UdT���}��bcc'��lѲ���f1+$_��P����>6G����6V�us�Аw�xg)��it�&wF�D�k����Ш��vhPH��U��'�		Y>R ��� �_ 0������y�{*`��4znd�&-b�}GFF^�8�q�@�2y/�5n|+�\�a�GC"�f���swm4�~��[�I��Zu뜴���	;��L��<�L�1�e��=�\�0W�Y��9C2:q����n+m��OJ+������rD^�D�:w5���WϐaÝ���G��� !�r�E��'W��$,`�
�>���.����&����;;Uf���B��k7`�dS�J-E4L�ׇ
�_�q��,'IlӺ�Y�t���?�i^ �&`9~�x�&;�d�je&O�����>M�a��͛��:���7 ��I��N����-
��7�|�c��:����s�^�������c���ˋ���f˜�o��Z�j�q �� f5L�/ z �6�����f3��n���w�@m��8.�G�VK�e��k$�5��v�W`ZU��Xh彝���]��6��D
l�����?j��r��j��d�@���U�OD�b3��_�� ���j��<@�Y�f͵���#���޽{׀c�=˹�U �n��f����^vK��y7�9>m���Cƙͳ͑��Ň�bO��02i����9_�X��޽߹%�N'��QT�鼳�}e��4��bsjo[s�0S�F�1�s��)�7��`���O�7j���Ʒ8���k����p�Pӷ����ܟ��C�zDTԭa�a/	�"�Y`���eXTp�M2�% �.�-@���9�4&� �{Tw7i�dhӦM��bc�G��DFFG��_��Ihx�����hK	
�,ǔ�A!!�4��8����C#�v�EF,�M�����CB��Z@7=84�f��W�����5�
֘�ލ��p<�����������o���68 @��@��r�U�x�����qF6j��A9Ƨ�����B���%��5�D�V�v���$��n�z���)�cwF�p��y��I
��^�M>l�p�i� ��K��� �ʿ쓻ͿA���|�7A]��X��ٺM;Ӿcg���Zp]�>�v�2%7�2�Wn��*Pn������H�����L�PV�ZUA��y��N7�������!�0@������x�y��O���#�m^��M�j�t�\�f�{�i�fB˖��^`���w��'�S*���J�w_�KԳW��1�zY>>('g����ǎ�k2��
N��OWԨQ�^�5r.��%�q.��kҿ~!���F��w֪S'�N�:����g_��#�+�
H��F
T.�{�W0�9ڏ�\�3��믿�Lrr��ҥ�	?!�^m���Ԥ���ݻw���˫�~�����_�T��˿�v��ko�]8}��oZ�x�H�f�|Y;�|Q3����@Lڶc��j���/#��ݾs������K?�^�����g?���S�,���3�p7c>�5f_�9�'���r���}�=��-�'�?���?��5u���i�i�7o�3�IԬ���!�!���B#""�&��,� �YX!��Dߛ���hFf�mY�[��HI�p%6���֭��&,<|aXD؎���D3�Ã3��Ʊ8� �X9�0���;��B7	��4
���4�7..����(�����	�@$�����*{�!��76
n�((h^����6
jt���s7ʨV��q������c�)��844�~h�u�e�kQD��������S�V�Sեc���8%\�N���B�V���:VL���2m��Q>q�����?�>�<�`b��=�ݺ�i+7v���|�7s2̑{������8��!9��6#=�0(�2 �|��0��@�,`�*�����6�޽1������$'&���Ʃ���_6O>���K���m�4&���/��㎏5�$
<�PG���s�5�<�yO���'��1���Ԃ�I߯O0cc��a�x���o�-֣�P�n=LW����M��N���4hw����#G�m��W�l�̪�j��>������"��������q�B�U	���i[�Ԗs���__zGe���cW�U󘼯7k֪�T��56T�S}X�z���4��E�{q[^���ӥ�$�* �.@9X��fY�)P���; ˧���?%P�~���?�8#ŗ]v�����\y��6h�`[jj�6m�t樝��S����;��b����g,j�U�]��Ⱥ�`�Å�a�<{(����q�[&���4:-�fi�y),�+���Ǯ=]�N��/�K?��c���z���G�?[tt�ٓof�Zt��FE���)ڟYp�^�������Y߼6�?#&�;u���W|Y��MZDEE%�F��

*���iڴ����I�	�3��Fu�ҥ[�^�"���*�2���iG������[6�l�w���L'��9$2lx����4n�\��J+ц}$�N
$p9L ���� ��&��g�BB�5ؠQ�����իmc��(bC��;7��6($$�,}�t�R��o#�F��{ϑcn��[�n�#�_���y"�YlE�)�#P��+��L^�*�n�Z���m�N����m�.պmc�3nC�� 7Y7`bɤ&7d��u��������K��gO�L�nݺ���T�Le�.��׉��L>_��䓒��c���ն\�n�%���s�i�%e��Q�(-M�y>���]��[�rFy��kL�w�?���w�R�Fu�L��V��jY�ܥ��>QW�X�:Yu���lG�-����Y��:���ew߱��>޻_�݃sr�ssGV0�W�^�j����v	P}Xy�Z���t�UMy���kR`��`P_����s�R�k�2m}L9O��5M�j�L�j%���t�\�=f�m��6w��B9�1���d��j�^]�v͉��w�V�Zȍ�J�^��+�_}��W]~���L֕y��~����]w��?���]u�U/��'[�ly�pŭ��ُ�=����_���	i��ܓ�Y�j��ꘒ�Rc׮]�A����(g��G�����5MY}<,a���x�uP�9�ާ�ہ̃��B?I����[ݽ�G���z�U�>U���Ag�������[
��`O��_�~�����m~�|�ڜ����7[o+x�kۂ�3�j>�}�����'O�C��'��_RR�aaaH���/�1J�k�ڵ��ݾ}H��ݫw�ޝ��Rm�����0j���i�ndd�,0z�����FaaU��4nҠQd�^2#�6
m��Z��اs���\c�ƍ�ҨQ���#M��׮� �n�������\cc��r������_ZZ�o#�Cj׮�&8$�����O%&$=����'11�H�Ĥ���-�U�L��p;�H@��v��m��D�*u��$���0=z�2��P#����Z1�57e���-{���葫mY�ҥ�@fo��w�4Z�H޷.}@�I�2m|�E�~ߵ��***2gϞ���\$��� �|�	`Z7vlL�f��S�LQ`\�j��̉�����͸1c����Սp2�O�MVf���t��r��;,�}�IhZz���u�hڵ�.s��]{Gm�ц�����5u^�M��.�q�	��٫��������;?f�j�
��h��.{��z+<���v��}��y_��}*qi;� q�Sט�@fY�h��r���0��W�Y�پK����	5k�lS�v�(�c�^�������ݔ�ĄE�_�U���4�N�:����?M��_�:�y��]���ҳg��[���iӦ_�x�g.��������K.�d� �2��t�%@Z��U�+_
�l�w�i��C��
C[jc����[���yZǈ�2	�����N��sY�����W���9��i�{Ú���/����C�$�+x���Ŝ)z�y���N�����.�
���)x�gt���O�Q��7�2��������I�5?�Jپ}�+)�[�~ܰa�+Ȯ�q�~A7�ٍҶ�@�.��z�RX��6vʒ��y9HH&�sϟ���xc|��u��*�ƶm��V��8((�1�))i��S[M������$$%m�"������I9%���)йb	(�*���VUU�馪��m,����ߗn�r����M�ڵ��i��m�������df�ֹ�){o���#��6����w��C೓I�t�||�	px`����m��0-L�Uv�ۘjǏ�q�?��#����[��Kh���Me�}��'z�_�������>��J/`�S�W7�ɑ#G��+W�;��l��vs��%1�v4���erjeb�ܺe�ٰ~���d4 B"8ID���~�.����M���T�ڇ�r e�v��M����=��4nw~�^ m׾��n�z��ݷ~���MW0C�r��E^m� �]U�W�'�e ��V��r���N��Q��c�kV?V�V�o0�Y1K �R�����>>�ZΧ���l$@���H��U����8��9����w��kv��l�\U��aY�^�jU��kX#� �y�*5jDT�^���������C�]�*;�$66��޽{_WO��f7�tST�fͪ�=�w�����}�v��$������?��ϰd��~���׿����\sM�אu��ɴ��Y���8>;�`���'���W�d��/�,��{��l;��~ȱ�n��&����v���O?ڒy��C[Q���ߝzL�S{;�8�'}}�Io�~7��y�	���N�{���)��>���˵��|���3�w�����`d�#o��g�~yh׏~����]/����3���ߐ��P/--��<i�����KLLڐ���v\��0���s�4鴑���rcP�rT]��wd-�eG�[�D��5|�e���S�N�]��YǍGnzN��lѲ�iߡ�Ƣ��qF�,.J{cvߤ�G��q��w��M��I"	���� ��S�̧�~j^|�E�${������v�ڥ�l�O����L�|���z����y��3�-�y�g���۵�%����d�_�?}���i�F���ޭ���r�ؿ�Z1�΁L�?7X��w9?�&��F�&==Ӥg|;���R��#�	h"�mڴ?ޥK��={���?�r��q�*U�^�F�L�řU�W�S@��*ի=.��G��eK��^�������e�C��JR\�n�@dE��CE�?	P7mڴ@������<�b���v֫_'�#���,�T��>��`�|�U��V>�,�G��ߞ:t��s���1""�w�0��;��K�.ɲ}RLL��k����%�\R�����F�/
h�,�;���?�y^�L�>Llw����͏Ʒ^y(&�����Íb���Ƥn=��v衬�X<�~��o�5 ���A�ֻ��Ak�n����'O�V\�J��F�>�^�SEG�:uh��g�[vꣅ�Oؐx�����_��`
�mb
߾^��r���дbŊK,����E������Ą���r�{96��	�"�&5E�3��(7��}C�I'���H�1��O
�ڦ���0u�[�QV�Zm[����:@��pndȧed��� L �f���nR�2T�}!JMCzc';�}�&U �aÂ��CZ��Z��,\�o�"['

4S���W�6�V��i~�bd�~�z��={��'N��͹SY�ɺRY��5Z�Côn�E��/��z��w�;|�|�ݻuӘJJ������Вd��;VA�E�LJQ�Qb�{W<�w`����k}�hl�"�L�-Mrr���T��WRr����&���<�w��yw�=�{���d���S��P�J�*un�Z�U����	��d��P^�'1i[}�@!���Z��J��>':"�ճ �t��*i����'g��n�t��z��}�G�������	l,@���Z��MU��"��A7U�֩jժM�X����ˋ�t3?y=��G�ǐ!Cb۴i39,,�a��|JI#٦�L�K"�d��ѣ��U�e�����_}��1�PR��4���T�4�Mp��ςb�;���`f�!�:��4���j�tO�G^y����O<����'�?����O�M-0o��?Ę���9�ǜ}�9�n��N�7��S������/�W|�������+2f�|�3�l����4�6lxUL��3[�L�W��8?`��]2������o�+X��� h�D?<:�R��mʶq@��R��Ll�jű�h &7\�21)�/{���Bb�B&�jӦ�IIN��faa�y����:�{ �v�?XQ������w�=�5z�L�s����4��:d�y��G͗_~e�޻�L�<�4k���@��.���H�a�m *�~}��%�رc歷�R7:I@�BZ`FFDj&y|���L-��7�~h�5�w���m�u�ݥK��޽+�:	T�R�7��ZU�T�s�M7�e^�p��p�5y}S����׬޷z���	$�[�Z�S�%`J?U,��B��=r�[��_PPP����qqq�PDD�|5�^kY�"ދ��M����^b�.N�u��u��隮]���СC^xx�C���o>��gE@�qы�����v2���8�����;���ݚI��P��ÅѩEG77G����Ԏ�����(��k���d����?�����=N�f��k�<����>.5�Ћ � );����fӳɦwi���{5*Blؐ��XTP��Wl�5*(ҤBzRHB�|�{vf3;ل���y���i�����3�ԝ~�89=���񄜌#�`B���Q��	���
r��mBj~���Ic]Q}cÅU�7�w7*�׷[hh�!,"buhX�O �0��q�X�	�`�����7��cK�������J|���?��/p��ks0_������5y����F���ѣ��>�X��_)c�;�F6����!�Zg�$�-a���%r��9Ә� k�?����b���<|����6�a�[+��A̱y����444�s�ṷ�xm?߻���1�6��=s>�:�pNND`�@���3e��d��q6��fb�:�mEx�>���8��f���%��LB�"n���#��?v�&�R\�	�Y5zLJ޸q��feM��}UM��\�}2����XˇK��`�B�����~����&Pl��&�4Y�) %5¦��:��S2��p���`w8��ا�ܣ���:c�v�1^���|z�LW,l6_�l٠%K�D�����۷�},�d�����}2�j5p�8�����
k2��G�č�x.&���$r�'�!�;�xaD�;�c'�.=��f���X�]wc�N�K%N�T�ŗ��s���B�$�T1ԓ�}��������)�MH�*��!��'����� ���nT�^�+(,(�rMPh��A!!�`:�9N��_b
�� �����
�Ѻ���������dR�D�ė0��CBï��!aV`F����D ؘ�;0�����D�sŧ��яv����ďvpn�̌�exb|<� (~�Hj�>�������3O=E���i����!K/�5��L>����~�C@����Z���a|4�jֱV��٬JH���:.73+��z5dȐ^Nry(��29��ԯZ�I<^`V���g�8�~J&��.�o��O<18,,,
~������pA���/�i�!�8�����I�&�����۷o��3Ǔ�{�&e�%en��I=[Oʼ#IY��c�Q��)IȜ_6n��餬[V�I��w�/���XW����,�h<v��x��������S����j~��z_�Er2�� �DRw4�\<:���_C�k�y�k���k������s����_c�ncٿ��s������F䶷���H��h��j���"�^��l4
�,���b��t��:�Y�J��Mn�ҲB�2��&+]T�^�qq.��!_��B�����YK`�>�AB��(>>��DG� S�D.�#�x�!�& �� S�G)DJ�g��_lA�.Lwl��{H�´O>��|��俟~J�豟꺧��}2sW���?��tآ�^{��޽�|��0������?*�9�#�S�=�g_����a|�9���Hk�ᙯ���7:%%7-3�&6���ϙ���
 �<&�����E�0�%P6�O��q�H��qV:��01�����3޽�����(�ʳ8�$$S��8����?������s��>r�L��+�������WĦ�iK&�}��|"�F��k2��nm�����y�'/�u�|����rg�Ξ^{(if��	/��_H�f�rԇ��@j�������5xo���5F�9�����{��O}f,�u��o�)�x&ǹ&�}M��!�O�8<cXž�a�!0�jYL�{���i��xuw'`�Ő�/z�2>!)�󂀉/^|��f���^lq��t���F،p9r�[(���-�ŀ��?���r� ���J�_�G;8���]�(4���+d��E`�ơ���sǎ��>�����s�rx�k.�p�6�sQ���7��������#���}��`㳈����B�9���@fU숸�Ĥѹiii�0����ŅsRp� ��  O�녿S��5��&��%D����t���/�8n)��=`2�i����._�|�U�",X�����cA׮]0y��%�a�رcg�7N��갆�T�ֽ4%+�h�čU#��Y4�T�Fњ̂���|Mf%�dޢ���vE�s��O?6�X���X�����Ge5G'�]�c�k�?3��t$����A'j~-���p�`1
"��l<M��!��I��/#�*�ԝXT^wd����95b���_\s`�Қ�Q�j�.�w�t�������s`pP5�����! ia
� r"��y�,Aޢ�{�ح���d"0c�lTt��kt�e,���/l!Nli�`o?���Kk�"\G����Qc�m"oJa]�dj�>W2yKP�wSk�'>ky0�`
��������K�,!?�Y��cd���tLa,�5^�r%�чx�ޛ���ɨ�#��m�~��-5�{zoxn����3$�%kn-��Y�B�C�R��!4���WEF�捌O�ML��yk�n�N��T���@�g �� �FӰdM5�M5���L�SN�(+t�d��v��9��~���aM�+���}2��N��"..�x^mll��O�>8��j??�0H���ȱ�h�Ĉ���/UĦ�ׇ%�J������E1c�.=qatn���2�O+7c�t��c���#SC/����E5GƿPsd�C����>�Tͯ�g�����|�����5��(�x(���H&�G�H�!e5��OT��?V�/ l8V���8�9���V���&�4T����%A�.L|���y�y�����W�X��/c|1{z�X}i_�����7�A���Ǝ`�y�������Z�� L���D�����ҡ��ΞMX���|�&q�_�����M��8�X{�y�F�	k4_z��\���K/�M��Ѵ��b�u���R�: �'<7���K��ϙ�Y�f|Ő)�ځ?��� 2��"�rcbF��y��^�C2�9s�ew@&�*e
y�LN]m�5 '5�CC~���V�,�}�,��8.���i�t�\&�;E999m?���as��}8&&�g�?�w���T~�C�;�odzJJ�����Ǚ��ZX����Y4:ksu\����xr�/��bMfx���	�ʲ�T��i6�᭖q�L��G��;r%w�ǣ/�ʙS}l�ڋ�'<Ws �Ś���U�{`����"^���IͯaGjD���-��p0�� �������������L�Cz�����p@p�CP��~��j���&`� E�)��Z�(ġ�L��[���ܜ�h��ڰvC!'.����Ϗ6a㗵�l����Rv�����������=��=$,���So`"l`m� t�[�>�B���t$�?�IM��j-�8�Zzk����m�����E�����Z0>�ww�}/���7�a��?ؽ�6��<����o�%�~��9r��믾�M�����5�����I<�����c6����SS��ai^��9�<�\}2q)t����W������!!���������/8�Y�x�	g������r�O�,[4��OΜ�g4����=r��i�B�
 ��7ӝ-�_	��=eʔ��i4ұcG�������볧O��iӦk�LZ�9fRxER���ش���$R�q��7�xql��┬�E���s鷼&Ӫ����?X}l�{��yaU��F_<6#��𤨪�Y��L��;6)��h֒���[ ��L�W{(�`������������o��VK�����������g/�jX�����}0�&zR��3�����4��4�.*K���Ee$y���ÛOC�4}� �^$,, pm>D D@���E�E_��8������P��M�1 �f���!b�4�f�l����倫���Ҥ�B���W��5I��]��&\_Fk0#""��8[�Xb�$6��]��6��>h����T�ܳ����w�}����������9���ӹ�����s�0=��g��R��qn}����Aڜ.ش|�y Ӣ�0<�_��������gT��0��Z�T: D�t��q�����5 ���̲�Μ�'{���p�t ̑2�J��^2�M�9s���iӦ��4h�ܹs-� ���
�9	k2!OO���4���잟2-�d�čG��N �� ��Yߨ�����E#���[��΀LlF?�l{������3��܏������m}/l�_���}�_���N�J�9������rk��ZS}(����bWW�������տ���7�t����{�z�kt�5Z���n������7��fp����!Ƌ��d��h[�A��_�����B~3�R��闧r9����#"�i�4|��K�22���X^����Р�PC�"#� �mbC�@1�rM�b�[�8�Z�X-�k-��t�|bKe-�raA-�E���! ���u�#���tIJ�.�u06�G����<:'~Q��jhpp��������� 0����uӁ�L�]��<��&��d��~����U�y�����m�	j��� dz�d�@Z�	���+��L Ǽ�3��K��F����֯_?hƌ�QQQ�U*Uu�����ڵk�ر�oC�����v��c
:�5�T��2��i�uᣍ���B���|W���q��N�W�<ٛ/r�E������ʏo�q��*��3�|jO>T�������cfP�S�j����o��V�`�������qQ�~v�j�q�q���Ʋ	0��Z��x���G��z��Mq�xsX���������e������h����K����/e�CxIӗ��˫5 ��^ ���� ���h"G��R !lϯ_+`
�Z:ZPK���ak�b�ӥy�i����I�bI�qݢ&\_�	���FCT��+������T	a��gl�ɉζ4i�D���W��N�z�-�`�<z�q��m�j��"�}��G���h�9έ�v�yt���ԯ~���:�=<��ݽ���=su^^���<�6���������k5����5�i&��NYYY�����5;�RԡC�CX۷o���ћ~���%K�8C�5}�V���#������M5	����Cy��r>'N����7��-K��s��'��c	��h<:�{�%�*O�������a�+�������n��*K�Ti�����0y��,`
�ײ�$�`i�&����m4���G��� ��U��cb�x���@���?��_�Wf,�
����ۍ��l0ai��|5�)H�)��j-�Zzki��&]�G'�g-^��<���m�+r\�{����"c�����!�ýA(�{���H�,ZD����s���`�Ԓ�=���-�9������wG�4[���Z��C�u#dbM&v�0��`I�r���W��=��dbb�Ԗ-[���'���=z��jӦM���m����'N̽������Y?>�U���%�J�V�>mCIbfq]Ę�"�`R��;~�հ=?p���)�gV����YK ӵ	?�qumLWU5¥y�"�f���L	�Q�k������el0E�6A�)o�� �h<7�@?:ߺ��D�`�B�Jcy�v�7H�%�����7�#PHmJiL�`�\�#k0%���ŉ-Vki��4ݚ.WFjA�0J�O���b��k��I�;�� H�p_�|����'���ceT\��g�$'+����U�-�vpAk(����3�?���h<<c��C�
,@&�d��x��菡*��.���=W�c���t'jٲe###3���޳���o۶-��Y���-999s����5�x�윞�S�G�dL�T���g}t*���x��9~�%`Ga��9E�&���Kj2��@aӒ0&��Z����z�u_)`^�M�!���b����-�%�����M_��/��� �؇5 �?i	0)���@�҄0�Z�%]ii>!�Z��˥_���[�4���¸����,�����2t�S��(���3Ԣ]��ִ`!�d�&S�Lk��yRk�U���պ�պ@lZ��;`bb���e˖�1113������ 4k{���@�Ë/���{�m��%����=K�慕N���d�Ē�豍%X�?v�5�����ҳi�L��r��ꄀ� �T�����@�Z�
0	������Q�a����B��L�0o���|M��kr>^��@Da: �\N�`�#Ǆc~
�2!Z}�_�(Gx�����p�LooZ�E�C dX��v.rk`u#$�6i�Zt-۸��b9���Kk!�kn�4�����R��7��6��{D�5C'_���q��`��îE�LV��-YEk@�v�T�Ik�� �u��Z��Vks�j5L&�;T��̈́	�����'}��%mڴ9eoo�#>>~�E���m�v]5�X�Y<cQT��Y�Ҧ�j1�\��l8�y�8��k23g��b��d�:�Skq:LL\���^�-��kC�f4<<�� �3���������D
5��t!�Ey�x
����s%n�/��3�ϯ�v]�e�U��T��y���d���t�}FF�����_LIIɗ�dFc�=�(��7���gM�4� �Ǽ澒�ً{M�^2y�ƊqS�kbR�e������YW�w
G�/C��y���={l�SV��ty� S̹(� �0Vm�2�]�
�͌ (�Z����`a�b:O�5hb|�b_Il&����B#Z|=��',q��z?��؄��� �Dn��<l���$��5�j��	��G*!�4�����Z�+)��<-}�c��R�B�n-|���į�]U�f�j���v��t�-����g��H�K�<#�*���c,s�%� ���ּy��>���iii/k4�|����1{��uH.��b0�=<<����;�E�I����.��,�b��3��i�I�{E֟�y��^�4�b�����rEk�pt�
���e�� �e��$��D�İ�&��a�P3$��u,�5�29G���χ��&����#��������o�!{��%����>��|*2�1���>#_~�%�����A*��-�km?R	y�����T��\I9�S�-�Q�yBK��G�0OS�4���)M�o�_ � ���.Ѷm�z�3&���۰a�Nw�С��{�������# �������׮ҙ9�+�,/��tsU��ӵq�k2���+��+KZY<s�Ĳ�_�*}�}������+s&�B�t&���r�2K��r�+��ˈ_�-_���.��Jb�KM[}�_��t�dV�}�IHh����h����Ν��~㔅s��!Ə'������I�H6��1�6�:y2y��ȶ�_�p����o�I-�\K�bY�#�	���Z�K��R^�k�#�u�j�w��|���t?>�R�%.��'6>Ohi<�q4�4�K�h|6�7_��'W�seJY��ڞ&���K�ޛ���0�z׮]�!� h��ׯ�fx��9r�`S���}�W�#�#.,xh}E������I�gx�Yg�3�n!�W4f���䮭x�_Y�ϼ�A�����`��:`b�K\���e.͇n���6XO��^�>�0�JKɧ�|B��a�386c�ĉ$8���ii4A(&*��x�Q��w�њP�Z�7k�bY�#�	���Z�K��R^��G&�g�����`21݅Z�v�}TT�R�V�א!CH�N�΃�><���/0,,���`h�g�f���^���9�j�->Q;f�1�$����"}왢�	?eL�<}���ݍ{����S���h� S��45�㋨e��~���&K�^MY��3�"E/Xi>4��?�������Z}����Ԧa���º3� ��[L�.��נ@D�<t�"]�s�[SiI	���ɬ�3M��v���u�Ȯ��'�����?�~w�NZӉ5����$$8��<����oo`������I�mk����6���=�|?D�Iz߄�-����(`²%�4���k�MϪ)l���>`	�y'������j{�LLw�p���̬���_I�޽�mڴ9ݷo�w�r�B///
�|��R�{W�	���ڗ*>\X�9�T�Ɛb��]Hm�gء���%IYS+Y�A��z�E��L�'&~��:`b��/}��9_k$LO̐` �0:��-L�ș3f�� ��C>H���+�|^]]MΟ?O]ZZJ~��#�V���n�ᘗ����!�O0���n�:-X��oѢE����4h6��.]��<x� ��cbb<}}}�����۸���^�S����uK��2i�_%��)q�����?���,c���Ցd25I� &,�J�K0mZ��fk�hN�ċ�
�4��Y��i� Q����[h��pi%](��F��|p�q��/k�`ia0��Nr�Wlz

$a�!$�`0O)@��`X
.>$�}���Y?���ys� ������/'�4^�t��eRmm-ٿ?Ll&��G~������������-}�LM�p}i�0����'�8�{c�� -ڎ4�b9����o%}�4����q\5��	��&�]�6��^Ϝ���|v�С���^j߾}}�^��pqq������s��e�K��l��j�s5k^XT���׊Ge�^�Z�ş `^*�8T���d���*���(]��5�3�d�
 L9��"�3��C�yK��y-ʃi���(���@)�q��6����]� �@SW,"�| �ΟO�oll�qɺ@��g
��8�&��ܹc)((0*�f�ٳ䣏>��� ��(��ڵ��~�y�n:z�Y��$u�Xz��}0��E��4qX�S�9`�ϘMa0� ��C�M�`s���!�]�|��9n f�ڞ}E��t7�����z��q��:t�8p��J�r����Orr��)���"����Ж?�Ҹ�Is�B?���,���"��B򵁇���JF�O)��Dwa���%��m�.���{��>�Lw����0��g�<,ZM��j򢛠�@�5S�}0[L떦�u3dr����m_
mX��#LF�1�ǋ�i�8+LK�7	#8�8q�lذ�$%&�m 8._���ܹ��d�߷�6������G!�F��ǚ>nye�r�رf��w��M�x����!lq?$iB؜.)#K�<�7�0( �%6f�3h2�a<<b05�Y���dU����2���&�ݦ���>���q�����Ʀ�]�v��ϡA�����JLKK��l7l@��M���{|�SْU>�c�fE�}�0p��Z�Xc�[pc�{�"���K��,,˘<�l����?R��[~�o�H�q:��BY����� S~9�(3�E����	�`����61�)�-j&�x���.N�0,q�"L|��x����`��01ʹ���h4��ˋ���R#�`M$~pC���qR��i��t�o���)�=s�TVV���RRRRB]�/�e����ɓd���d�E$*2����DG�I'����/'K�,�C���#�2"& t9ٳgԒؾhw��***�ؠ�|�d��5$9)�^s5 &N��t?���9����i-�[�'^��^4�����g0Ep(}��qV�Mi�q3��6k`���� `>�T*�t�u���]���P��V�<xpmϞ=�?湾}�����sill���`��72�l�H��T笶+H��\�x���	��cRI�Odc���t�&�B��=%c�߽�a�;����G旿�S�w�=�M1���#�.R�D����]=`��b~�R0D_`Z�|=�)us�4��p�� Lxx (���Vka�+0� ��ׇ��CV�ZE�������M��]�����>���/�L�H&&&P�u�s�j�D���m��PM�0���K�.%���
����-��n2��G ���>ya��d欙$"2��x����ޛ[a��Zx��4��웞+)\�d�I1PJ�M�@*�7�8�~ ���~����Y��s�2���R��u��;`bb�� i8�����A�j 0�ݺu;?�����9܈a��)�~%�U:}�[%㦖UE��.�6��y�]�ƒ�ƆG�h�ޱ�����|~~��IE��G��T����0��E��5�sq�g���k F��C�4�6�7�+�#؜�������De�M�a�t�ʖ�q���76c�&r7�&r�e%۠�<�G�eD�i*k���VȈ�Fc���,��0���#�q#HZ�82~��q&��l������C�t2*!� �*���H�F�J������>�8:;�i��z����A�O̢��o}t�bK��ǵ�Z��xi�4�q���ɉ$$,��{���C����5�Z�&�o-^[s�<��;}��gH��D���#�C>,#
��aڎ`xk.���aX��3ǭw��9q\
�q:p���bbb�����Ǐ�GFF>9dȐ}m۶ml׮]M�~���P(x$%%u��pm�2�x�ʔ��K6UM��Uq���m������ᄤd���HŲ��+r�r����O>�.]�/�����,���8�#�0`6����k����^� �ti��6�1�1���_J��i��+��ߴoY���s@a����Uc��̙�Hi�kK~�r�vd���`��>e�}g���>�i�<Ұ�8<v�>o���i����8�v�BX��y��;��&�Wz-赕�1]�GH��`s<oqY��e,����#�?t]���0<���s��2g��7x>�@�F'�i)�e�������������?x6��]����)))1...�0��k׮�T~�O�> @�333�8p�#����x�c+sք�/_��|�C��M�W�0n��J!� �� 8�c/����}q����g�)͚�P8}�O��e�N?�dg���a/!����۞䀓�Y��A�� � �k�*��
U5�m� f��@��--o��
E�/��^�fK���(`��չ{xk��O�j5'UZ�	���$�I ǓN`\
�?�8� ��2*Wד��,�.���p}M��Tg�ײ���Ru�� r ��p��'|���N�gƥh}��!'�Nr�W	e\���K��Rk�1��
6�R��2���'�rr�`;��_�a{�x�Ri��A��x7������A\�nڞ\ ��N�N�~)]\,�ss�v�����/N��+����±�}��-�&<R��p�?�� .O X���ɰ��%�L��Tc��p9��
�p\21�����1b�f��p�����k��@��Crell�+V#��4�H�]<y@��7����3d�'�<���M*�zR�����s���
�F�.�M{�d���%��GVdN�T.X�P�b�=���Us�,�?�+�y��U�*�6��	��>p���F �Z���O7��s����n���|E�s�
0�U�ɶ:�dtٚ1�-�qs�
ۣK�n7�j�z+\�� [eNtIǂK�%�U��<<����2����Sl�n_ǭ������q�ۿnsWl�w��?��fG~��5��f:G����=�c���h���$<Spn�y�0Z��3�M&��
��E'�l��L��M�����t�K&&���BCC�̘1c�رc����w�ؑ�iӦ�W�^����|||b"""���0�}���}���י׍�����򛿔���K���b����8R�K
�C�=��?��y�0(~nidJf��	i�f��M_�znɣ��>��_����o:�:�:ErG?�M�u��4K��t��כ  i-��/*WM�J�&JW�Ț`��[~���� �@���O�ծ�괓6S5:]���5E�P����X �l�B,`0V�ј�"����tt)M�Z�h�1��S�������dO�XO4��|t���o�n���܈{p��ј��s��e��K(��P��r����kWx�כLLS8vz��<Ǎ�(���Խ{wҾ}�pa�Ν�ݣG�E��|=	!7���sO[�w��5�#����7n�\2m����윲���-M�jlL�@ʽ#I�*��@P���W��Q�G�[E��o�ĥ�Qz���e�?]����K+_��Z</ǹ2c�Cq@���gt��z��<�!2�j���'P�R�R���h�j�:A��L
�7�b��%�5��:���J�z�E�2^�*��?{l>tpp<|��!�*c�������l���x�b[˧Ӊ�k���m,9�;�V��*��2�j/��aC�011ݹھ};�Ō���y�)���m�h�{��ڵ� �d��70��sO���G���i��zi���^V�箛^����/���uYX��u�2ȹ�Ѥ�;�*_X^�	,-�**M8];v_Q\�{ű��K�RgǥN*K�*�GM*�{�O*t�T�6L*T雬�8H�<������)�n!���1�ja, LO�R�P��~���Y���i|m	��&mL�H�����<M��x�	F �8��l�y��t{����r�A��*�H������|c��v��$�KN�5�<�2��Y��7�_|,����,�)�=b[+�Ƽ�����6o��n����N6=����vXK&��rrr:M�8Q����000p�εi�?�)�ׯ߇���s��ݵ7�rk¾��/n^�|Ud͔��s)_����?L�瑒�$R�j�W��@c�.���#�.�3�l�g�����{
��w��/���U����3l@�|W�]�.�&C\�G�G�*��]��Q>��Ca����Jej�P �D���%/o�^^����(���!�,�Ei����\^'����8.��ٹ/9�������:�t�s�����q��ݛt���,urrz���;k1!�-�2c�9��tNN��^v���k+�z����+>*K���0hԗ���_��cN�����J!#F�b���'�b�WD�#8�d������@�_Sࢇ%�1NTS��)t�-����<��mP��:]'�B��j�zzy�v�����U��
��M�i��H�f@(2��D[K�b�~x�E��!`*�X�Ʊ-�������F��l���;t̘1Y �_>�����hccSfgg�_��%>>>���m�����M��*s�
�Z�hl�Y���S2KӲ��dL�R6q�OegUU���X��PWW�	�Z`YW�������͇]�
4�uEn!ue^���]3�.q7�U뚠��Wk5���Tu�́m�+3�5� S�»9`"HZ����v��{��@ǅ�~�=�,w���5'21111��Z�n�MFF��#��T��:w�\�8>�NNN�CBB�-[6Д��	��>0-���-=�_zm`E��ʇV�)[��ъŏ�ra��ec��)���84~�Yߘ� �;
�A;
T;
\��q]�;�5�;�=�vz�����v	Ѹh]|�*�"�J��B�,�4ZLM�x�n�?4"\^0!�jy�m�-�C�E����R
��) �"�Lv[�111111�Hmٲ�ӂ4���9���?���k׮�gϞ��nޔ)S�6l����-�y޶r���E9����4�d���y!%f�&f��&�zD�jC
Uz��4p�64�TZK~L�K��upT9�9�声��m�B��R�(�LS�QT�f�i�K�,<��7M�@@��K
}R��&�4�Ӽ|:5��ô���q0aد�����4 模C��c?T�2011111����믻%$$����}����}���0`čKKKS<���|�;B$9�#��>�������]Ξ=k2�c\lv����+�@,uwH�ceoo�I�T��a�0� ���:`6��҄ZF�P(��"�����\���x{M�29W��-�Ӝ�K�����gbbbbb�[�*�4iRxzz�{AAA���o���:t�~����GFF��7o�M�Ϻ�1�|ѩ��D���E � n���jbp�R�Oq5�QC9�2)�YX�y��8�ٶ�a�:=n#@j ��2��\�
�P��������wR[�"r���S���>���{�A��Y1`����z��iiiq���v؂IK01�L�/� _�r�|!��' g� ��(�� y7 &��FN./���\��OgggwK�cbbbbb��"�t�6m�����a�������ؘ�,��������0=rrrX32���U�vr��d>�)� <^@H���G�G
�&K��y�M ��צ>�&���|ؔ�di��iszS9��%���p9 Ӟ?]&&&&&���  �GFF&��}����)����~������x&555v۶ml,h�[#�@����\�[��"@*U�w`�er���s{er�28=�7�&�s������wV%e	�'N���}��W߹sgҩS���Ç�JLL�������ɱ��e�n������r��% �� j�Z@Nl3��I?����fy��"��2��8Q�V� ��2����L.� ���J�`�߄������� �},X
0���ã|��������;�y���Y3g�Ԯ[��;_��馩��� Ȝ�)�� ��L6 P�����\�i6�V�y�����9�.X���m5�RR�t�se �������� ���	�?F���˗/<y������=�ߥK��*GG����ћ�͛7�駟�Y���1�<%ߓ��e�˽�R.W��+��1A_�Q ɛ� ���Is�V�T&�2�;�ɹ�e2E*�!9`S��������ڰaC���zj������^�zU�k׎t�֭�?eee=�x�����v���'�n�ưI�)9 ��p
�i��s��W�Kj��dNjQ�[`<�j��s�r�4����-�8�J�N��1abbbb�ǉ�n֬Y������޽�E��ׯ_���߮Q�F�HJJR!��J01�D!d�ؘ �Q
�C�R�����9�3.!� z��b��	�y�0ߑ���|�2��>8�v��bbbbbb�ǩmBB���)SR_�<��t�ر�[�n�;88�	


�>}z>?�MW;'�z�R��)d�X�)�����m ����\�E���
�qP:�c�ȟ�?Qm���� �� L���������4h�,ooo���Tl�cb�%j��h��d2����8���N�pLx�x������If5�LLLLLL��s���`���9s�lNII)wss3���m۶=�׆6#,,�+;;�_����g��/����{����1��z����������[�zuҌ3�EDD�:t(�ڵk����{�����������������tY�ټys��S���������ή�S�N�=z6l�6��Ok2	!l�"&&&&&&&&��?�8qb|tt4e>���ڵk}��ݏ<��^?-++�s۶m�&����������ʄs��������l>|xY�^�H�.]��<��������̤�$ϧ�~�'!���dbbbbbbbb���.]�/888^��l6lXѽ��Klmm/h�|��i����5k�8�ԓ���l�L&&&&&&&&�֕��� s����6�\^��iccc��C�;w~����ѣGg̛7/���wںukWS�;W���l&&&&&&&�۩)S���WU*U�}��Gڵk�3���ҥ�g:�nkff���;w�z��L%�<0w�S����������n�6n��;55udXX����g���p:I�ZX�rss�&44tSTT��q�Ʃ�o�����ӝ���c�7���)���D*���6�u��ټ��۝W�Z�g�ԩ�����|>&&&&&&&&�۩����OJJ�=z�+#F�(��� ݺu#:th����0`��� �����s����������999��M�4�t� ���# �=j�(9�_���05<<�)>;��@b�y�捚4i�Ƙ��O����,���!�۷��ر�o}��y���q���ۜ���)iii�f̘�b�
�-[��ܽ{wl��͡�H=p��.���]6l�@���M� �԰�NXC�����;���u8z����ŋ{ @:!H�3���NW��Ӈ6����aǐ!C~��011111111�)�>����~cǎ 7K.��(��ѣ���ܹ�7}������¶&&&�=ztژ1c�a]��驆�؜V�.]�hP�>>>����t���⼽���B|PP�N�����+����Z�v����[[�O:u���i0�N���������t��}NN�mnn�p �L�]~~~� {D&��pF��y=@�y �SÆ����a����# �a}~�~� �-l۶�B؞��\اO�!C�, ]2@r!@�����xyy=�P(���ۯ�����]�2`���`�<����U]�v��СCl����O����������!�mLL̠�cǦ,X�`�i��GGG_�͎;����Ν;���]�^�� ����C��mڴ���Ll��@��gϞ�q�?ww�O�Z�^77���ju	�U4��{�� � �a{G`�,	��o@���ھ}�֪T��U�&&&&&&&&�;Y�6m��g�I}����|E�P������Gggg���#�ӧ�j�q4�p��K �հ�- �@�y(_٣G\'8�֒�k�k#�Fi<�2�0����O����qppx��������͐����������N�dFGG k����������Q�F-T	�Y	PX�X`X	`y\�����8��ِk"�]�vmD�DPŦn�#}���(qlN�k<x�y�FS���wB������^���{��`��>��#G���211111111�%�9�;�F�C�u{��G�S�N����𔗗��C�}@p=��F ���K�Qp�\�/�-�,suu-p-ONNn��� S�L!˖-#O>�$Y�d	1b�O��ί���?��@r�1c�ϟo�gϞ�8fNNN'�N�z����������n ]G��A�G�vIIIѦ�����ǻ�T*�;��s�/�w�?�ضm[�mmm?T(�;����܏֯_�����So���ٽ{��9x�������H�V���W��p�M65$��P؄� x˖-��u���ph��$�4�t��iݻw�֯_?j;;�i^^^S��ӧ�Z�jګ������{��>[���G���sΜ93姟~r����i*;�8�hX��3111111111��ۃ9������+�J::  @�)`T�2++K�q�F��o�)P�֯_�����8p� %�=8���`GGG��3g��<�h�K���`0pN,��߬��������������������������������������������������������������������������������������������������������������������������������������I�{��6E�w���Z    IEND�B`�PK
     �8�Z���1�_ �_ /   images/fce5a045-7211-4fa3-86b3-f57a3d8041ae.png�PNG

   IHDR  �     G!��   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx��Y��y.��jOgH΃8i�'�R_$��<p�v^ �p:A���p^h=$�vұu(7}e'���$���0ҷ3�#���-������{������jU����CQ�'���ګV�ZU�ַ�*)'N�8q�ĉ'N�Q�t�ĉ'N�8q��� �'N�8q�ĉ�m0�8q�ĉ'N�l�8��ĉ'N�8q�d[�L'N�8q�ĉ'�*`:q�ĉ'N�8�Vq Ӊ'N�8q��ɶ���9{�l�>J��㞺O�ڵk]��}1}t�}�ٖr�ĉ'N��/���������}�	�`buu5�}ߋ�(��v�L���xԮ8$�v� �I sQ9q�ĉ'N�w� �},q{������V���O���y^�6�@}���\�S����gG���ע���v�_���J�r��fG9q�ĉ'N�7� ��+������&��8����'���J���@�Ve#uJYj f@q6h��}�K�R���
�}�~�q�Չ'N�8qro���T���/��t:��{� ڏӮ�����D���їC
�D��,؏6���v�Q�i�ߢ�����sM�@��8q�ĉ'�^����3��L��c��P{��>M@�ijg��#�Y2lᎶ��4��f4���S��J�r��k�����r�ĉ'N�<�� �}$gϞ�	��n�ZGQ�Qh�� ����R/`�SR0�6����tvӮCT���@��=TN�8q�ĉ�^��O�V�M�<M ��\>I?��C �0�R������F�>V��vR�k�y�����c�ӭ�}�s���O����8q�ĉ'�8�y��������ҡr��8}}��0;pi���`
��0��1�[Q���
ȴT�#`/i{��/�������O��O\����U�ĉ'N�<�� �}"�Vk��%�,OEQt���� �1���Y&`�8J��y�>[pL�k�>��7���n���~�]�'N�8q�d(q �>��gϖD��� X?e���{���SfR��SP1����D��r�]�������b�T���SO5`�6؉'N�8q�0wX^|��ॗ^���jG��P�[|��/�<�c�	�
�����]������<����8q�ĉ'�8���r�ܹ0�Q��O��0'L:ȡ�Ф#l �9Pڋ�,b4{������m��dN�v���:{���[._�'N�8q�`��;,�Je�>A�����ō�d˝��)"��lN����S���n������K��ʝ8q�ĉ�L��A���>W& 6kl/�'�.:��A���{`��Z�;��7�>���}����OѮ���������L'N�8q��0wH .��߿i;��a���A̖J�����m2����+���j����������)��G������@0�ĉ'N�8y��;$�N�������N,;I ��	�� E�b���qR��nB3>h܌���0&�	�S���v��	S 'N�8q����.`��,��"��/��},'5��)�2�=�K���D��<U�ߍ�D��Ù�O��A[9��Q�}�Z��g &�x�;wn�ڎ��MNN���e�X�?���Ř�������J9q�ĉ���8��C�lּj���[-�T5=_���,f�ǂq�3�q��S�F-�8��l�Y�S���{��٥/~Q5��b<(����JƢ�c���[�v�`��	��v��j�ږ�޻���~x������2@��+��r��^X��_�ED0k�"^V%_��L��Svs��
p���n�1'N�8٢�s��V�`�#D]*�ix��Tvފ�ڼx���f2{������CZ!���),���vч	W�#��hP�,�J����r3���&���o�fO�A���^�5����T{��Ukkk�k��O��O���ו+<� ?��?�Μ9�*���>��S��T��&��8�'�s��]i�8R=$�[�̮kK��>�f� f��j�\ZZ�H���o~��ϵ����O��Pǭ��v\�,����?�~�~��%�N�D�-ct_��8��L���������N����<���_�e�/�➣6<;xn6.�+;���P�ҹY;��	!=��g�}v]9q����P��A�	8��H�Gk̔*ҶB����s��^�s�+/:L��8�ĝNg���vج�[�V�2Kx�G�j6��ƍ��ŋ&i}eE��u�)Q�N��9$�˟˷o�W~��~422�]�z���SO�ݷo��j�z� �n�o ��}}�~���d+wi��p�0O��&�כt�]�|���/�ܘ�<ám��N�����?�G|G辀-~��w�w�����z�-]���J�+��JRR��͛7U����M�.\P���ZRO���[��@�Xݺ�D�X[ݾ�yAP�� nNNN.<���Wgff�?��t��ŉ'Ntq s�djJ�F�W	\�&�h��l
+j���uL�y�j/�;J��}]o�h�3
�)��(��d�Y��N+�	lǱ��"3��Xߌ��l7��ҒZ_]������*��~ �7������a�	����J)f?��;x��!/c�v+0��u#���ʠ���q����u��;���ś�o�_��^[]�U��<�Qʺ�>u�!]�e�F��vդ�"�����Z/�o<�"�,�'�& $�g�ꡅ׃�bqq�����i�gnNU�Ƿ�"o�t��W�T���Ju����\���ܼ�o|{�[���������ʉ'N�� �} ې��=!:G9�2?���N��c�5�݈(&���ɇ��J[?y	 �:!���Z��sy< +��U`�Ӥ�E �M�wJ�`�ƍ�z�1;666�f����,��&E�E� �~;zG�� Wq�:�?l�}tn�`G@o�@�v����/޹p�K�~�h�A�D,�P/��`Di�w,*To$m#��T�\�� ���j�N�X�S:�zw~^��3����|�?B��Ž��h�$# fl��X�y~X*�W;q|u}}���.z��|�>�Ο���}��G�|򓟼[&�N�8qr_��;(P�u:L�%�-���n睬l��`z���c�Y� C��N8J�+���w;�O[\&:�Q`[�B*���NYsט7O��Z��{�n522¬�Ҧ� �^�m�i�_l�:՟���L0��۷o�<��j��z}]�Z-U�B�.>� �X`�����`4	���:�^�1������c�0G����*}|���������+W���y<s.�c�7U����Cv>�Bz8�(�C�@�l����CT�j˅Z��ʍ7.Ёʉ'N`q s���K����h�ՠ ����Pq��/T���R�_�V�0�V�Дnh��y>��~p0:�ެ���v�
�T[��A𞉮t_�!XE�7��q	�@O�oI��Կ�*�)s_ˆ�ʆ�cY�:J��YQ�#P2��}(v��/c������a2���`׾�:r��!`)b�y�z�� �k���Y��`��S^����X��_x�6��~��.t�'NHq s�d��1���L_la�4�:���^�U�\yw���<GfK�tn�u-h���nےnO�N6/lQl=HNOM�={v��]�j||B����	�- 	[���( �`?���j4��A� �p�*��f���Ne 0W�w7��.�ݭ^��8��q[��$�uN�ŏ���e�d��M׷/�o0,u6�N�8y �����|��W�ߏ�e� �[Q�<3�pBq��8���ql��&���R�>�JP�~�ڎ��ķZ�15�BV�>�Ӄ'O�#G��ܥfgf���,�L ���5�+���Kw�pT�[7o��n޺Ŏ;Ԡ�.��`�9 �jX�L���a��{fS��d�^�L'+ӹ�"�=��i{sbbb^9��ĉ�T��1�R�-�%Z�{\l0��>8I�,�Fmˤ�Ᏻ=q�9Nl����:61�4��'�b�%��U�ԝq���A��������w��A6���k{���m�������܎�ˁ�Ȅ�$B��r�x�6	(..-�[�K �%��жx���}�63� �-Q�ù`��y�����2���z|K*r���'�w�`���(��4]OP�R�B[��l�l/��ĉ'��8����x�}�l8��S&u�������Ocԛ_�� �.0hP�r� E�܌D�& 	{�} �n�SK�>�%DwY��*d�JuK��!{`���U�Z��sLWXJ�y��N���`�H����jue���v�h���503�v�!�.frjJ�#ޥ���{)�r�^�,/3`M�����z+ϡ �Ԇ���;���6&���]A�<�MMM+'N�8yP���Hl��ٳٚ���*��:m6j+@lX�fl�0�] �d�g���;\����Ӌ����J ��'��E���֪_����� J��Vߨ|q> ��=!�Ђ��Չ�<�=-���X�2hsѽG] x�=�k͗�)i�Y3�U����J�k�W�\Q׮_O�o���q� ��ǜ4�_991��rrr��O |f<�M&XO����;�$�ӎ	l+�p	p��&��9<���&�P�ޔ'N�<�� ��F&���;�ʝqoę� s; &D +@�ݼj��`���@E?M�`Gb;J8#� ��,Q�B��@�B��! T���|,T�8 ���0��D�ǥ�e�E�>�V�dN����۷o3�D��33IF#���i�+�X�u�����C�Qg��3u�K;I����Y��苹={Ԯ]�i�����!�9ɿ�`�]S�
S�6&@�ZP��0=�_J�[�L��*�h��N�8y_��;,�����s7f?����04�	 �m�%��[��Ma��þ0���aˈ�Z8��⢺z�*�_~ �X��N�xOMO1�U�I[�����z��%����m�U/�!�υi�F��^���|vS{&	���*wVMS��� ��>:6�0�b�i9�i���Qݢ���&p�ݧE}�}B})!�����I"�l%6�&v�����1��7���c���H�Kl ��3I-)���p��0.S�Y�L���>^TN�8q����VO�Ɵ��L��F)�J�R��m�����WWI�]
{�] S�UJ ��>V)���^}m;�^E�{ �p�	��jTi �6������E�l Fb�X�V���,�Y��+��lq.�y�8@�)l��ۧv��Ŭj��m��rE-HF$֧���Q�G�0� &�n�΅��6�(}����C���'N0��%�� mx�HJ�D*O���T��clYy3!�����f��{'��Rsc��`b�TDE���3��l����ĉ'�8���bg���};�����o���ɠ3j���Y�$E��n���l�`��޻���uÖ	���&N� ��>��
�"����6Q��SS3��N���`
ep^��333�'�8r���r�����0����s��P.�B	L|vv�*i��$�{�G=]nh��Fݸ��ǎ�2ٌ �m��%��[��d @6�Vx��q�A�$�0�y�X�J�&�0����=�}����[��;��ĉ�W��A�$([~����幸�b��us�j��>;\��X���8��/*�2O�`普��E���B�;*	#�O�u{� ��0�0����Ph�J�Rl��9Ѵ��4���1c�c'D�i[㲣���l�K�_��ػw/��]�VX<4��B��
��(K����@��s�����8@�F���4f�e��܏`���"��}Q�O\[� L0�+F��J�K�L�b"�x��I+�|Þ���������x���0�ZEf�R).6�8q��A0���p٢�{%���@6	ĽqIA���aӺ���K ���4�#<�9v�8�X�D�F��1�D,� MX� �"�"���M%�ْ�+Y���X�_8�ӌ,\<�, lF���(!�D��O �۷n1����v0� �pĩ�Q��۔#����ŋj~~^{�S��h�'�ͥ�锴�Pi3�j��]�*q�%�4~���>x�/��C6���/��u6�� S�l� �^b�9��Չ'N���F�L���:F��������K=��8kW��|Ȝ"I�@WdE��VTK�r �$6k���m�7��/ �f�sN5�a4U{'e`��e�j�������ۿ��J�������� c߾}�z���"76� B��0�N���xCW#�5 I�#<n�
&�3�F];j�� q i����������x�Tu��	�m3l��i���*!����:Y���;ڂ>��*6I0N]��O׀{�L@\�NB�;j������ft�<�Z��E/r/QW�AI;)� SL`�!�vF�N�8y����l���s$������p�^m�V��`�
_\Ya 05���ر(�ea����=.R�C��ʉ'�
� J�I/;I[p.0� ���ce�O�1 �)��9�k�s�&6�������2�'\ڋPH��G�H�y�s���=��8��㈢-�/d
��A�cw��O�B ȐE���&�3�h��I_g��0�`���-̔��f⡊�\G����1�N�8y�ōr;%KK��,T6E&�Ai�l��- ��ٛє��[�37��  6�ZU$ 3u��ߦ���|/��9$Ϥ�h���/�T�r������}���L�7������M n C�dv���m�'ϊ�n�#�Nǌ�fb�h~��3R��R�/�M D�b���L-[��-�&�o�*�Q��q��s�v>����(�E8�  �
`����������jj��9�ę3j�޽� �×_Vo��63��	��NN��>97�*(��Hi��h�̹05sYMT��̄bj@��N�8y�ōr;,-I��60���4���1��*�DB�=�mLۓ���"��,�	��eb0n&E�0�9Υa=�~H�u��q�)jw�� ����Iptd���-��~�!8��WQ%�N>��]�z��F��cN��� ���C�"v�vF�aDT�hL>���������K��>g��X���au��cG�r�/����N�������Ǿu��������V���j����GyH�NA��؊b�L��-�m0}��3��L��O|�D�������d��϶�'N�q s�6�;� ��	��TJ�VZ�0bZ�}���i(��Ol;H���]'�N���0ag�Z��x<w����fk1��)��y��dz|����~/N> 1`9Τa� �\r���~
��Ku,`R<�YnlT� <0v`� �����|;m/�]_D�h�_���� s��GH a3�����-$ ����gJ%i2��<�]���s�q��_�;�k���s�Կ��&�)8���yF�:}�Y�%���|�ט�<B ����̙3�ƍ����˜�Hy<`���\*S_T��>*��ر�k�{��J�� �� ^a0w���~�ת�����Y�"�X��ϳ3���%(�ϙ�����~����_���P��9N�8��� �N�as0"�0������X�35��)W�g/�.0g�,�	<�r`�-�A�0x>WSP�l2���1J �J�Jv42l�������?:Ee�S�8��r��)âe.�{Fmh�X��&mf�� �Je8VΎ�	�J�u��q����1��W��������|�j��Uuca�ۅ�1�G��1�u�W��˒��!�8�|!�,f.� S�&�/�]��U)�����/y��(O�v��;F��g��ei��+�C}������]$�z��_�zS9q��}-`�L�Lְ������{J�W�K?�n1sZ�v5�0�ƑI[D%Z*卷Y�VI
��e~�=�j����՞�`����$6;�C#dXH0sy�i���{ ,x�#v�8�$�����{Ƅʷ�V�����$60�p�aU�q�
M�`��C���vT�[`�D�666#Tyɳ�y/r��W�[o���=�z�!���;��s�?G �8?�;��*��Or'O�d�y�悺h�I�t��~F=v�g0���`�>� S�>lP)�����x��RΞ=;J�������=D��70�Q��y'}}1(�I7����9>;;�2�?������p���-`�,Y���`c�S:�c�5�1��zyd
�/��l�SQQ�5`�p�	ֶY`v�1  ,bK��v_L
�WST<N������8� سؔ�: &�n,1����{m��e�6� q@��@�E�(�����H�U6�*�Q��NT��)Hǚ���s���E8���S�T19�{���D���?��¢�M�G�8s�G���	��.S��_�C]x�z�7����,z�7N�. �F�Ǧ<���k�3�v�,���N>��)#e�F��B�o�>�P�>H��qj߇�� ��~��a0=s�`0��*m{�� �r�o:�"���J'N��8��C��c0�<{1q�f^�})��ߺ��R�L�?&�q���-Xe0i�$N!�F|o`
he� f�`r9�vU��Mx���=�mVK�k�Dr��&`8>� �d�o�4XGxU�xA��|@s��	52�*�ioiV�C�m�X� �tx��2�DPNr����2g�M�m8���{��H�a80�}��C��IcK
f���k���bQP��,�s��jɧ����=JT�`��3(��ANT��%�`�� L].�PE����{*t��o��o��9B�{�>?F�Gh���9�i�x��a���� ���6}^����"`��;�����T��!���.����@��P�m�zɰ��W@������I�iv�)���I_��E s+©'���� �S�kI�WQ��R��T��Q�ԫ�b���(��,�a��L,L ) (,@�����	6��q<CP5�Iu�� ��Z��n�m��E;!|���<Pr_o�k ��� �����Ģ��%�V9��	�.v��#�yv�U�F�C�f��y��%u��wl�cդ��k��]1��gp����%�S�����ō�"R �}��ԓ���_���*�L쥶>B_?Fmz��r��)io�3To��3|Z�Ҿ}t�.�=z������ԉ';"`�0cؚ����V�V;̽�h�����m�΢�8n`�)��	���d[ ���ð�q5�nT\tPϖo���KLKl�+0$���>�mdbiX���
s�rH����#t��¦&W:�L�\T�6����s��2��M���"��i��@0�<�pB�<�L����"Q� ��a� .����/���ǿK` }�8��	�/*�2gH��k�7l]X_ۦX�S��E�X_��	A�}���6<Bm:N۴8\�ڍ������X���^���ĉ�� `�`��$�����,q9n�a9�6�Wcy=����Kҹ&{��ƳW{<>&��4^�<��"�Rӊ�l��M�C?U㚲F�nk��h�^g#ҫO��I��l���'�Ǒf�s��, 8�0@�$kM�,g W8��-��:����[�1�ϻ�s�g�0�rG�ՙ�Ly�b��Uц1����l_�A}�E�=�8opH���ܛ��,�(�� G�B͏����׏��D�oH�ST��ӊ7�&�0D�R�	��+��Q����cz��Ԗ	�@�禮M؋�����Ǚc}���}��qz6�K��ĉ�R��Ait*l���6�P�!�	�Cj��A��epȕ�e���/u�<m��<��R�wy�wו�]�d �����a���)N.�Ad&����S�B�  P�6���~�:�����D�0v#	�����b��4�o����{]�|�X4I,�~`E�"q-HWy��9��#_8RB"����عЏ~�^��6��M�`���[&����.MӠ����է�e?һ߅�����f�d��vD��bj�@3��EvD��
��&���t��4���gϮ8G'Nޟ� ��8�Da���� ��@���(�q|-�&�Vc���z�V���Dؠ;��@��l�,9�6���Z6��^�E��~lϤ�0K�R�6��QKÉGT���F� �# "X= �U�}e���\��A�߸���U氿$`hb�pq�J�\�O � Dql��d]����ԯ�6 ���	�����ko�����?�p���Z�J���E����z���D�:�Yo)����.c���z�r�w>�� Lapm��5x�=������=����{'6�9�͊�/S��$?I���v�·�ʉ'�;q s�d~~=����#�!F��qj=f1KU,�����0�n\}������&��CN��!Gl� "|?(��t�,``����@�����nI(�� ���4m��	�3!����CH�w��D���ˁ�K�<����i#�Dl@7$�^� |��WX��� �0�4�ĩˉÏ�� 4�,��%��A NC�ű%a-/z[��] �T
�Y����0��u�o�)?��O���?��gff&޿����W�\��3U�6��,%�.�*�D�I�u���L�Wמ{�:�/{�����vj/>��cɾ���������?}��^��8qrߊ�;&�4��(�ه����v�Z�uo�x��C�dk,��8�۱C��YmX�ԹGT㉭�q��L���"���LJ�Zպ��J�a&�d/{�Z�~��j����	u (A�"��a� �e�5� �hX>�t��9��L/�]3�5��mY%��xx#�5�r��)V���k��A8�K�D����Y��X�T1?�~�m�r Ϣ�o�(aQ���\��70�UL�%�<��b���q9~q�>D`��7oN_�pa�رc~>�c��JL�я~�#ħ����B�M�x��E�$r� M�_�9�ӽ9J��]ZD@5_GY:�P+?��3��� Y���qoϟ+�K�_|q���r���})�����mo���24Ld�۸��Ѽ���x�؋K�3h���WL�ʫ��Ϧ�)3�o䀭����b.m������f-P`n����$�&�P�T�a�I����۝$o9&׹={�� ��B2�,p� ��x�v�\����B ; x��g��X_#8��>�t��A�]�!j7ڈE�|�'�,�L/ '_ Ɇ�n��'� ���}Ŏ>`����u� L0�҅y�`���_
�Α���O�5B�u���8��v��[��,f9\YYAy�����(���9cZ{�*r�;�j�X:@��Q:���0=k� ��2��K�S�+j�V�:�צ�ݡ{��w���\��]��c��쳟t��N��G�a�����c����o���3?�3�[m���?_���M�1M��b~������瞫�}������K���?��?�x�"�Whռe���O��pW����(�a~����0�[͚�a��ډ-f:g�m!�'�ALZ/����n����&֙T�nNiuyl���]��^���ڔC$��v�X�z�������0-��vO���1'sNc>�5f`�')@L2�A`��@�}$�N��{��ȕ�O����uQ݃�3�?�?o�������>�N>h�s��+/���߸������ڷo�w�]S��/��~���38��SOq~�cǎ��T���&�l{H[��ro��P�E���|��8���]?�1������{�������wQ��c>B��S����}����3<xx����	�&�6� ��.�׌�\V�|`J��j��-G��g'���)ME���J�k5�Z�wZT�j��f�����g���������'?�PN�8�/dh�	�Uj�����J�h|�������7/޼S�s�s��\��X�����7��M��t�dRG����; eզ��[_��s?��z�,V�4�T�>oyy�]D����i@���X>7�j���߾�߮^Y��X�F\��Ko��v����Yt��g6A��\�26��tµ7���_����w�,�7��j�6����k���W^9���|����1z���d���U��84@�FL`2�-ذ��G� �3�	7�툿=C���D&b���b�3�7� ��Ϥ�{"qm���H���0��J�����^6�v�i�*ܿ&�㞹9��#��G��������7���޽{as�N;P�/�|��y������v"���O?Ͷz �P���*v4h��˳��2�(Úh��w� ��R�s،A��v�Pi�c����݈]�G*����.��8�z��q:�|��9�8�c�y��	 ۱������Hb�L<X�x8*a\]��Q�ik�3>>q��
ޢ9��SO=���8q��2,��hB��P��[����(�
�N�V;w�ȑ�T�K�K_����4`L��&0v�+_��M�t�����VW�O��W�ay=22~qee�?��?~�������//����7�xcW@A�^�:��5��/����f���Z��v�=U��oG��N���x�.�[��[TқM�D����p��[6���j�u�]�?�j�G��(*W�k��+���T�e�-}�_�M+�ِ�l���/��/v_Y\|�������8�N���fA��`���E�F�W�#c5V�i�ejl�nq>I��nn}��5%��Q���Xl�S��b���,�H.S��m�s�3�K���RH�]���ٶ#�Xk���`�i�e�@<�qo�w0��1�Q�@��G�aB�͎;����De;Ϲaq]m`���~V�����vǆ=5Ɔ��w�˪��n]Q���ER���G�4��OFil��z�"�x�E�k8�E�'�i��R�Vן�N��G�9��F䙔�Rb�6z`Hg�(�G��z��x��i�[[[{�������?=���'N����80Q��������ӄ��62r� �X=�?��?��ʯ�������7/]:=Ҏ��
s���A�|�K_���[���=�|���G:�f�^����lu��T9T�������@����W�rhqu��V�qd�6V���{z����.���/+8���??J�#�F���K�?֬��LLL^�����f��������A�;����?�O�y��ɶ�Y���R#o�}WT��ݎ�G���X^]y����+�{&��G�v>�⋗�Mea��������[��Õ�V�V.����/�M�2�r���W_}����ՏѤ�� ����G{).�̱1�����r��*���m�0��ޗ�PmE��)�x�k�m�P���x��.��*j;K����i���pz1Yn��@�׆aۺ���w�e.9��N<���MNQ���܈l�����`�
?��f�;�'N�PDt��@�����O�l��=z�����_���[��7�d�����s���×�@ױ&����tcM���P	�9��7�ۇ���WĖ���;�+�_@�oN6�;k�9k� ﳾ��<a�}��L��sei�(���T)��Z��K�}�C���N����.��l]�c�kk�.//}��h�!�f45ɡ.�Ju���赉�����k�ꫫϬ�՟�Ib?��^��������Wx��痦�ҾN������3X?����p)(Ǔ��v�Ӊ�Q����?��?��˿��]+�����G���j�V�!r�F�]��������/�U_���=~�u|ee履��Q�{+��B�Ռ��������Ͽ~���x~a�t�>So5��a{o\��)�t�Z�j�o�	d� ����z�}zuu����'i���'&G�0n^Xh�/���Ϳ�˿��Zk}���T�Q?����\-U�Yh��{��ٳ�r����֖��^]Yy��O�o���8f�a=�M�HQ��<��n���G�vKb{iX�V�m#��ԭP�w��a���N�2�dRL�i������QA���U�[�{$ ����nQ}��Ζ�ArmE�3���7�6��V�.��u �?4�� ��GЈ����S2@��;��^�<yR���i[N���~���o���^��9�KVJ��˰��;�j�~`�o�aYLاS_A#`��a�1~�/}��8�>)��|f��ISl���>�߽�2�Q�L4[��V�1M}Z�Z^���_������?���ʉ';"G�cǎ�7o.��Y[ٽ����@�����W�¨u8]'�VGW��]o<�xg��VW�ϔ+��##�m�(?����7��^�4��olyi�a�$�T���<�h6�JP"`P�_~���4�6Z��i�x��֓ 3ht�J~<Taӿ����?�^o�ZZ^<���t��������(�6���q�/uv�[����Z��v��c�V�ri&��]ϜG��j��^�q�G#�Z�z���w�,..3H)G�#�V�@\������Buv7ꭧ���3a':{JoP[G	<���\�u����^�c46~���	�ơJB�;0-z<Ӷ����'Y���Z��33˓�^w������̶~��|V=>���VD΅>hk��W�A��(æ&�Ui�I]YļHx���f�0o�.Y{t��b�#��� �Q�yV}�B���@���든��}N�ۆ�.\� j����J_���c���V�wB�>2��=ߗ`�oܸ�v�Ⱦ��n��� �Ď������$&l3�]��޹|���x�K�e���8�7�A���J�Y�W�����c�����e,�mX;N���#XW��=E��=���}�f��\J
�RgɘP�E84�#�k������iv"d���w�{�tL�';!��?�-,�����R][Y�4��HՐ]#�@y��b��{~��jF����=111>��*�j�h�ʯ����Qo<���tzmey
6�(GS����%?�jA0��tnݼ}{jiy�1��a����yS���ڡjMu��:�əՕ���w�Ͷ?:��-�[�ÝJ�.������k���������v�8]\m�BF���T�G�`c��^Y��X�s����ʸ��(LEg;��a���u�EQ���������c4Y>L��>\�	�4�Su���h�Ꜣ)�	��Q+�&�b^4@�1�$E`�m�1�K��^����N�2��=�c`=.8���QC�����f���s����n�#Ƚ6/��< ��:Q� `L�����o[�[V_���~���ˡ�<��VK�E��1+�k^db��|���>,��z�? �8�C�a�F�༃����8 �\X�b�"c����88I�,3V�O!�*h��l݇����{����>��S�^����x��Sk�l��g�xi���)��u�꽚��I����"�P0��y[V������H�+�qP�=/��%�,-��;^_[�L����_|�ܹs+E��N�8�{2`"�H|�;��	#5���	;!X�z���?�n6���90��N{TO�Xq�{i���F*�G��t��~�Y��4��N̄��Mu=�{�)B�K���9D�,bBTUA�4J�qG4`{�(\��d��j>�^�����5�U����{�f�C����}������~D�N��Eh�;�1�M�{����f�9M���׬i��T����i�^^[_� �y��l�a���D�Q���6Ka�Cm��Q{�z��*��X� C��c�x�����ԶL�Q���쩡ۥ%΍�c~�Ք�y���v3)��{��v��G�u�i9p*A0b�J�K��&��}+�X�H�X�r���]�-�hb� p�M&a����ԁ����.�C��`�"p����)>;�h�M�MI 2X�mp�M��aD��Dm�ݵK�߿��Q�o~~ h�N���P_!w=��Y	m�{���P�����"��`=�ܳE�|#�[`��C��k�N���{��W^���O���?}��??c�^o��=@*F�f'1�P*�@��{%����]Uls)�y�0����~���Y�*�*oe�?^�_^��5�<1���z���MA���[T�r���=�� ��������
<?�M�k9x��(0B��aA���k����D���YPB� f}�G!�m�����F}m��b�"(�V��� ��l6k4��i�����M@������h�S�'°=�j6W��F�j5g:a{֋=�����Z<���A�7'h�[Ѫ���/�@4�Ϩ��Xl�u�P�M�)S3�/��7�����V������Z�7���,�	�3Iͨ�u�j�[A��>�l��-f��e_��W<�i
������/��3�h�a#���6G�聍�!��m2\����If!Q�i[��v���|��fW*B��Ȩ�ц�:w#}�$�7�kq��f����N�h�Y�����y�����:�9�IU��^�`������M��6����6��!Ё���o��Ȁ���/�K� @z��QΗ���� i2��ƥ�+Q�4 �tm��>6��Dt��;w�^xa���F�'�'yТO�^��/_�;>>v�^;E�Y꛲�9����}��6Z���,��=�wMX6sZT�kα�)�,�Y��|�d�i9٪����DkG��V��;��Ș_�{�֯�꯮)���`����P����/�BR@�G]iOg�5���@Y"8���vi��2ƆA�^z/�SP_��V=L���"��"�r[k��/-/����~b�g1t:����[���F}7&}������;�"`W����"u^���L\5�J����3K�8�G`y5 k�ۨ�%����T�Y_�6���b<cK��<�J�B����VY}�Y�>�8Q��$]1i9Ӎ������+(Qdy�ߕc>=q��כ-�߰h�0
����z�^V�߿�W Ą!x�m  !�0mS��"e��X� �RCCPv� 6-��҄��g�%$P�L<x�Ă�CYL���c	��1!Qgĉ�,�*m`py��I��+�9fQ��S��ӪK��4 Di���G������S���iFqdɼi��³��F�t�U���~ǹ����%� ����|D=��3�R?x�ڽg�[Q�~){�`�=��O^��^emu>��@��������8�]�vm�GYB�\���ܹse��I�	��L�R~�Z�!�DBagO��1�6q���|Z��T۽9���V��Z0{�\����w 0�<l��ؤ�͢��8Nl�Y��6Bs��V�E�f�36V[��v��ٳW�}�Y�݉�{ &���(Mfx�S0$��؏�1�yl�%޵��c��4�<L�`���L'@���jM��#�p(	�@�O�(���6����M�L�~Yqh���a!�D|]\B!�]�ྶ� +N�	ZV}����|^S�dD$SUm��5a��������r���M�x/E�Xje�0Mbd'DX����-�&�?�s��1�����t��5�tn�105�Z�L	���m%@ځ�:�6c;���,�{�*���L}� �ǀ����mF��C��.lhc,mK<�[\΁L9�Ȩ�%TXA�EZFxo�g7=���f�Lɓ�*�('���qN�/*}71��П�w�z��E�D$���(��i�Φ��O��cBmG�O��%Ww�sq����A��#bSW�b��U�7Ӵ��TjO��x��ڬ���ʘ�%���o�v�m�=c��e��R��e��q�����l La/�]��b_���,�b��4�6�#�J��z�z���z��1�Cv Ӊ�{ C� ����S����.�@@����^`1�8j �'KN���%_�3F��f8j �f��z�-U�0�Q3�[��sn���^bw��r˜��v��%��qT��G��zSpFU�ύ�&��¡����NԆ�̢�|c�\a�)�t�\�uc�2��W��c�Zʮ�/�:��[����C����n�a�x8��h���%6�����S�z�z�*滭�F*Ea3���~��!����,����:��e` � b8~jz:c���ۭ[�؋�l�B�����D} ��>0�6��$�2 [ }��D������``qwn���6�P���%� '�F��}�v��Pq<�qͨ��wo����������J��,� ���K/����ϫ:�K�d��k�8�z��S���i�����u�Q�୷�B�w��qڎұ�@����e�'�ypdd��Ǚ��}ok_� @�(�IS sZ#y�&?��Ӥ�&���3*l.ޅ�D1�1�ș�G�i�}�r�)'�RR���+�@�2{��	L�GV�V�P���M��H�9�r'N�0M�9�0H�*+Y<�(�Ͷ3�4l\�0�z�0�x2�g��N��+mZ��s����lԲ6x��w3��=����Ԃ��E)Ꝣ�����*3�%m�ίY2���H�bP���K�C������ӓ���
b�������@H@�x�BM56���UML���f3���^6���V6���֨d}�I�] �MjGvz1a���u2q�ʟ������H��g(?U���:���$��ȋ�V2�c\E�o3��lD��mۙ,v�8�!i��믽ƀ�eL�~ڔ��-�L�}@�	�s�y�O�]eN�|d 44#��D��	ϛM��n���ůx�c���55��|`�E�X�a��`���䬩R�n?Y싓���z��-��m҃����Q��F�1�nu�5��J��y��sUj8q����P S��ӣ�̠0R �6(�J<��T�f�S6x��/ԓq�&�9Z+V�Ꜿ�� =�T|/vIp�H���� ���6+7�P�5�V������̊��$��g�'�U���]��(`z�	��8^ f,?�$ٕg��Fe���3iU6k�;i1���ɶYX1���C���&pj8����{����O⊎�Ka��^���\ ��|���x���CI�h3�C�3�h�̄`҄� ���Fy�E��L�P�f���C�=�v��B�.,�0x�~D����'��v��@�G}�s���~��k	M�y��*���o�����f�9/���Ye���w}m-�/5���z�3�-�>W�:,�5g�uс�A�4e��1�jV�X�N�A �D�8��<�g�q/�X�R� �� m��3���0��~X���O)Y�'㼹���4��T����o"�P�ٚ���CaܙW�s��u�����au�ĉ��&�s��T��1��/PJ@�g�*����~�Qٖ�֪s0�IJ���a`�T+�	�2�Nԉz*�m��!(m����mƑ�|#�A1V�.]l��Ф�G���R�fXm���ä� �������S`��K#u�{QDUV*|o$a��@��0ѱ��,���a���昜v�$`w/O�q���8�;�&�=�!@�	^T����H ֈ�����`f<<G�s��)	�����i�y�m�����Q�]���U3i5KF�.�>�1�։�꾗H?I�9/7�v�C��~�%�{�h�W���x/ީ��gs����f���/� �eouƩ���e�c�60cel��Ĵ��;[�/ms߄���.��H��!�-Q{�J|o�=�����K$��w�l�ޅ]T�P'��Ɋ޳y�ĉ��* �zbf%��:�v�)Cl��i�7v��v�&+rF%��L���p,[��SXQ߬����W��6	̊�2��.�<߀V�Np��CxI}���è�+X'u�z���̵hu16��1����b�S���kr���֎^!����.ӣ��"�z=c�sH����q�d����8l�?� {�!�wn�'<_5�a����`� �8ޢ<�Y'h�v~�l9 	 i"�L@29� ��w�=	3��ձR���/�`d<����z[���S�ۦTҶ�*es�	6��o��KZ1^����*�d�e?0d��K��<g+������dQQ E�{=_]��V�l&4a��dݘ�������Zm��&�"� 0G���q>f3&�E�̶�͖�+ڇ\_��z�P�ݩm��Y��0SM�<�v�,�9M�̻e۹��u�}
h�V�J�
�~T.\���=r��%�b0��R�mw��� G����(yZ�i����� {h3qj0**rZ�V+I�3���"q
ЫW� �@h�$����6�t�NQOu�%��Lk$�\�L��*u�v�W7��V��ʞ���B���$8pv"I�3~AF$e2't�����r}nj<D���d:�S�)�-L`�yq���F �m��9�!��ذz�CT����o�ԃp|�[����v������Po�I�8��tN�������-�����9K͐�k��p~Y�$m�}+�> j~�m����(���`�	h�	ԟ�/"�.`�tQ��F����8f���j7݃q�#U��̃�.�B��-n?��i.�CP��1�̡"�/�6��+�}+�94���K��wX�7e�3�-�s
���͑5�lo�6{s^3���Y+<�1��W0�d"'D:rBd��h1�(z������^ԛ�	�.��w+�A�&,e��}�A+�x]:qr�es S�̃2��|.��Iզ���7�<9T�&^ɴa�4��1x��4�'쏬j�v3NS&�n�	����n#�D0��ء�=?�d� фe����H$kP��?ub�%9�u�c `0��xti�n9o�%i3$]�ݒ�����@���֑=Q�3kif���(�,5x24��/b8�� �)T� �#ƹ��[���+<;��c�������wl3++	���8!�0�����0v0S��k�,���8p@ǓB��T�`q~�����mA;p� ] �lSJ�%�:���@PB�q*M��K>r1�d��"���|\#����0�yI�+�H�*�f�{L�t��2�#йs�tJN�����,�,�j�yƲ�K����]�,".��_��yv�g��9�	Ѕ1:2�H��&L�	U�!���+�L��v'ed+�:�Ԩ���^�L�iDY�����y�m�}���L�5<ZMa��TS.k�'w[6 0ŋ\�![늓 �`e0a�i@&��a®� �8q�)%y�1��wV�0c�i�j^��I0� ��S��d�8�	���%+{M����x8H��따���&{��Xc\�;)�t0�`kbn�pF)����eY0�R�qW1O�\='��xY��S� ԓ�9V݅R?ۆJ�+�"����̕ũ&&���{��ԉ ��q��8K�;L��	p��l��VŊp� VPV����<�`s	�e�v�</b�����{N�%��
��{��w�| �pB��m�v1�Ƶ�Z��ˮW���V����q(���,NI�����1���-���V:���?Π���K��i�[}%�9�=ssl!��;�/'�����|�������&��12�y� LϨ}�<��O�V;�l���@�q�� ӌGQ��n����ߚ���ƙh	�����N>=3�;mZ����� SL$�m�:
 �g��t�DJ�4��ղC٥�o6m���AL`Z��r���]�3�¶��Tbl�AETr�S��:5��a�0P������F��u��J]��#\�fB�'>�;}�ð�P��Ы�*3e���Aݳ�O�-��J���-20��ᇠ�ĵhe�1FM#�Xz��ssVʄ��NRz"���!^��q�b�̓^�c�D�)p���d6���( E�Cż�>�Uc�����q.�	���`�L��"vL΋����`��ofL[-V%Ë��������<���v�E׀v�� a�� ���[ ^p,�P	i/[����3�6������>,�0Ib�,�BT^lM�\���.�r��f\��r$�/NA����������.6����*3�8��̦o���q��Or�sx�g�涠�%Äf�Ș�H�6�;���0R��I��^����b�*�J�g�)��Ѥ��s#�|ؓ�R�f�����.0�ڕ�ͽԩI���q:��ơ���B)���;�ڧڡ�t��Y��v�K��`&�pO�='N�l�0a�(�"{v��f2�T��E�3;	��O�J<��g�G�(���I�tZF=�%�) 8�{�4h�����AF�,�笶�B Imfm�o��T���j0QiW��o%�:����e����~
�F�V��d2�U`
S*}����4�W��'Q�b%sh�H��03rބxȟ'=N&V�3�>(ϔ^��l,�^*rLx X�	� P8���<`�L;Bc�Y1a���3	�jl�71�@P�)f �J a�&�Z�[�@��à���A��I�I��s�<�v�p~Q�L��R	�Ơ���;	,q5����ء��>�U�Pl�z9Iyy���B��y�C�ox�ӻ�멚L-��-�~a;��hq ���<A��㞚m����er�{=�E�)NU�ɴ����� ��e��l�c�W�E�Y�Y��z���m2|��<�5������M�'�I�����ۢfu/�N�����t���j�JbXB�� GrudOXcI��.�����V�ۑR�"Q��܋F��$��욝8q�9�\�"�UR6� ����1��eB1`�0�`�j&V���jS�bZ,"Tϣ�#����L���ι��������$JQaYQ^�ICFb�jA Ū���`������`�5� j"-���]R���|4ò�*�҇V�����Yd��T˜�^�Sl0���'��QOji�x����c Dq��9�"�9[�jہ��Y�{Y��[D�*����ve%�@��e��n_`��r�E"y��v�~L�, $nc?�w)/�g�.�`J����ŋ��!����ǹh�dh�;��ơRG_ F'lO�|���l����LH$[e��6J�01^�X����L��2��͌����бcI��4�ף���8����5��6��f���6aqU�%���7\f������]��)�����4ˉ'w_�� M�Ķ�*�D�	�&϶3�Xv�����\��*'�D!�0R�C����*�'bYA����z�m�ƾ�픨,X"e��D�F *A��\L��\&�f��Z�L�=��m%�n��̤.v�FaS�z\�i�
(�l���^�wӐ�kV%+��P��F�L&{J��r����@/�,Q{�$�\L�zč�viX�hP����Ym��9�=[&���3 ���  bۄ���y��*;�f�-Lj�8���@���B���^�v_I�LQ_��e�}�s� p��N�3ز��|�BywV����a_�d�O�g3�q����}�y$d����|��L>��cj]�;Ｃ���׹>f�i��S��1N8�`��&�)qP�ڒ�~���"�3
�L�{�O�&-�gRI��k
L}^`k��ު�a�v�8�.�W�i���8��)����.���˗���9�'��Z�k�����0�v�� �<����z܉�{%��)�ި��GX��d�0�x�ݢ	�x�%�3�(�eR1.3^�F���u�X���bT�,� ].���e㐣c8�&X{�:�F�s�X���/GԦ�<99��Q��=�Y��Xn�$ ��޻����=LN�VB]��3Uf�u�Rf����(+^Ѱ!�j���Z�����p�C�s��a�� I��d�T*aQ��Tʳ�O-u�8�wh#�;�|��^md3�L�ۜ�sv���� ���TqF�o����BN/���C����}�? � �X,��c�Z:'�k��! ��ʊz��79W�믿����6�;'̬}�HSj���Y�f!�`b<�ź�^�(�!�p_{�Z���5��f,ݦ��a�o]e�e�orD��$p���]���#�lJ�q�1�A���%�*��l��JV�+J�/�q�эf����h���k���tN��,�oɵ�S&�6��H}�˪*	�΁��4�4D���{
T��JԘ�-�u;/غ>�����VSS|Qp����v?G�eмJ�~0R��w����S�I�5�m	%VR��6���^��)�W7	�Ud����zq�7f4F��-�����-���ʠ	)
�EX�Q΂2�vzb�JPtB�:	�#�� 0" ǵ�����$�R1�>7�퉺cʳ�''�%���^}�׈t��W�����Xv�2�# �mkl��Ye�t�-=U�r��~�?�,�B��WϝS7���984��������k�����`����hUtd-P���@���)��Z S��ɱnM|�
�~���EmI�>Xd�� V5�V�^
�(�Ӷ*�"]�%��*�� �׼:�������!��a��0^x�8qrwe�6��9�Ӹv d���D%� ������s�� ��ldx"���*	�R
dd1��ί�Bג����Q����m�N"6�\Φ&�`F�S������̸Ф�I��#n430=3�����Q��ՕU��n�Wν�@�ͩۂ�z�A�x'���y�&Ol�t�f!!{���<ʞ���l�'?���W���J'�@l�</�8
�
�P��aluŖ�*/��0���y��A�gv׎K�k��<�P��2�#��Y@ޓ��Ifk�QG�F��H�=��A�9g����� E�)�jv�1�X���'��v�.Yhj[k������Ӷ c��8�޴Mo��O	����M����発 �ᤵbR�z����FD�4��3ԡ�L'N�0i<�hl0c&vR<0�l���*\]�6���%+ wܭ��Q�R��xf�*�a,� �pt��$L�iu��S�XeU�A�3�ѵ7��&f�6�&;&{0�̎h[<0L��0�/�yB��6K�/]���@�lp��HmX��7���R�E��v�b6��O�p��f2;�8_4�ó�3���R8vɗXv�<nڈ:SX���p;&΢�B� ��x1�n�c�}ý_7�VO�`&� ꒔��@\�Z$~���Lx:�'�d��x�g�Ί�M
�,��{�~�g��*u�*f����H�S�j_0� �6�� ű�Մ��)	�n����1�}6��h<�n�d�m��vD�Gږ�kN����]�瑇�Ȁ�(�_]1�4Ygth6�I�:��<�ö�We�l�E�*��ƭ�m0Ve��3�w�$KVf�͵��]��ӫL�Ҡ��e�rsͺM�'N��� ���k��+��L���-�R�(P#Nm29n��)����jN�.Q���A��0�<���^T&4������0�_e�LC��I&��A9��%Z8P4b��E�C���f���&�Ѥ�D���L�	����5����y>�ԟ�$���%vt�'�xh'v�8g�7�f�;���X@��ԋ�`��,�p��l�%jj�ե�+��\7`�-�dV�^����;S��-�v�YA�|��"J'��K���u����bV�8�W9BB�"�)l-%�|�W�[X�1E�/	�.,td��Z�(0� �mI$���( �`����u--%6��GuO$o��ĉ��C��-�W
K�=�#^TXۏ�@�c�b��0a@��F��'�c�զ���������������%1���"º��e���a)�s��	6l����!|��Cc�9���M�P��_f���|6[����,I�,�(LCf��7cyY;O��M��,��jY��6���%dg�0��ɠ�-\IL1e#���jd�-~� l��v���j�(m���q�A� ����⹞^b
�l#FM�rP�;?�����$����mg��v���"��jl�)ǝyj�$��:l��pP�(�ə�
���酮�U���v�J��'r�092����̙3��c�Y�b�}�k�`�&Nc�y�;_���a&��z�C����b��B���� CĮd[�M4<Kx$Ԕ^Dz	�n�����e�/�c{|�<�=� ui"�8��1/�Ȩ�-ո�F�j�W9ae��k�V�����`{2bo�$��V'q+d �V����=�n)Pg�8������$�b�K@��N�v��D����-Sڈ�w,�Y4�v���e�� J�T`�<�����L�~�oe��>(�,$`�g�f����.Q�S�o ]�q��O,�y( ϼ�� l`%��/�uZZ^NT�6��O�bgֱlXT9`2���˩3�ߐ��$�Ax�ؓ���\� �Uً1�c��k��zդ-��e$����yg��}K�K]R0&���I�)zlS3NÐ�9Q�g��[����n��.B��M��m�)c�ޯ��o�EE�+�,�'N6'�LZ�F��u�7 -��Ż��� /��_fG�	��d@��S��4��<���;�YoM$N,�N$Πf�0��j|�j8E�`&+f�Ä����Jv�Ƃ�+y5c�خ����0]�c(n1?�����5e��
J����AN�u�b�UMw�������F'\y�p�;�ؼ����S*�!��,T%��Ӌ"�H��[&��)��;�Y���b�a�������|�97Ά� �p����<� �bYt���"�MǤ��#�"�f��!9�-����8&mm�:�G� .�XD���f��[[*�H��S� ��8s�� ���4��,/2� �����n�I$o��gXV���ޔQ��Q�a�UԎ�0��kK��M�
{�Q���m��F���3��K��Am�M��#��h�Θ�$�\��楘޳8�jX&'N��� ��c~9���`j5V�7���Ab�kj&1N.��=N,���'�ڎ#c��L[�8c��cEU�\���i�V���[���X	�ډ�������.���G�}Ńn���;��]]Z�M�W���tU��NlM��$!��:�H���\;�p� �.`�6}Q��(	FL<C��������=/�/��0Z�� qm�"��x&���˗�]8Ι�Z��������q���S�5t���MH�9I��e�(!����u��8o?G's�Q%�\��}���<x�c�F�%F��zӰ�h/���߄�}��E�#�xe��A��a�Q^���޺fo���~��gj�S�ז�1�;J�UEW+��f�
��H��)��|�a:�i��ubU��ё�x��g����]�� ������[��I����E��,"�ڙAK�'D�W��k0**�$���(��-Ϊ�c��He�3����[�>��t���0V*3`%6K���"��e�Uw��'�1�O�Kf����~M��'fx�2�e�1�4�i�2Q�G�Ԇj�E�L�$�3�!�(��"� ��d���r������8^bj"6t�2�J�[�H'U��
@ ��9f#�x�� �+r,���)���#��P)�bKb����- ۰sD�LQ���%�<2Ô��{r?re��k@?r��:��'Ϝ���3�� t?q�mPi���Wd�]8b���������r�M�l'��Q&����0v��^}��Ŭ�K3�s�d���i��,��p��U9��Aו�a�Q�q���L ��d��v������ɉ'wW�g�yF��M5��;4x�d[�P�?S�ŢR��Uē q�of2M��
 �,%T��%���X%�&��
ö�׌� �3�d�TY��ӔqT�5)��\O`���6�R.k�YF_�Λ�ɏ}�Zw5��:s��<{z�z�M�Jk�͈Hd�>�q�y�����VȜ�j���Y��++�����!�����ȑ#r��]�r����IN�� tX��kۮu�m ��g�͚%9�41��{oխ}/j/�*� 
(��`z�%S�� =�L/2�I��&� ��C�<���$3�ƚԓdݲ����A�b#@־jE�w�����q?��y�- �)�fd���GĉϿ���EP�A��A7�+ՠ�Ջnh"+�V䍄/�Dlk��al�Qɨ�Vf=��s,��hc���mIB���|JEJ��O)���F)Uȴ0E�T^o���y��q�i�f6�_8��%��Ut|�1�F�������'��(�Ԯ]����s�؝<u�����$c'n�E�N�iU]�F�@�λ
�Sn]5����n*�5��X�1<�����RQ���2�ZQ�n����_3xl#U�ȅ<E�\c!B�X�6�F_M���U��*��"+��� ��?���?�ݿ3�o^7w�y�Q+�<���`��ga0��ɇ}n|�l��b�mm���*c0=;���L�Mo�X{%�qP2�W��+�~L���ڌ���0�:��(�&�/e�	�~�a�X���M���)U�X|9ۼF�������꿕�U~v>�_��kd��B����}`=�����}֠f�{!�f>0�����,h��M ��4U̀ak�J��a~`�mhK��sö[�m�L���\A$�dX��2�Nd�����[�E�×����~���O�kn޸���5�	x>��|���D��w�s���������=�y49&M0���� -RX���k?R���r��w�bq���	�`�4]K��p������3�5u�p��������Jb�S�<mip�Nu��R�6г��6�{�����7��/��/�l��Y�?bi�9+\�;�k_EI��9���Gq�gc��(^1��A�~���ɦ�NW���EH� &��+�I#ߥ|�?n���rs�"��թu��|:}_����)���~v��E`*�1n&��]uN��Յ�wjۑ�e�_R��z�5��^L���SU�='R��%���I[#`��_�p~0�"��> �6 -`5�$��۷�`P���W	��W�@��	@�_#̲�`s6|��h��i[�[�f3��\�oh��`bgP����|�.�{8'�p��]"�/qn0%CЦ<�`�%a/e9@�,���TQp@����I��c�n;m�� L�GsMHS��e��~�8A\X�?D��&i�]���V�}x��py�O�9��q�ڨ�6.����5���-��L<�%�ϻ�n�{��fԤN>EK�~�����u-i�	ji��D�0�}}�ѣ��t�������_��_ΙY�Yv	0�9�hެ߰�l�!�o�C��'�%�S*�L�sa�2LRvV�Vj�la%M���i���4.1>h3�vI�;��͍����@�x_9�vz�{h��V[ɽن�����j�"/���M�UH����Y�.��Ԁ:Ec� Ϊ���t�!��S9L�H΍�?)VNٴ�k��]�r�\�� fm��@� :`��An��\�D�M���a��/����(�ю6Bz�ِ�ru�x�{�K�#��5`(�a#�%�����O3 8h�c���r����ƍ��ɓ�O�� ��H`Ԫ`җg�������k�10�/*X����w��3�ҥK��t���_|P}�y�~m��>ر_�&��ٵ�l<)��PUky�V����'M"8���lB|�)��g���USSs��];5աg�^�x��?��?���o�ֽ��;���6OR�`C�p7�����$#�O~�fuv��G�}��p��X=c2���쓀��3
 F1ig �Z����5��Z��U83�����:עM`Њr��G���`�3�/	i��*�)M^�D��f�f���[Y�/zG4d����J\ݶ�[�r����Ě��ϰ���{`L�bN��سm�1�j+���{i~~!2�b.F��J�6R�����Gx3�\�p(�������$�F"r &��!O�s��r�T�6UR%�8s� �K��c0}Ċ��N|�� Ti	���%�y�? ��Bfi��q)C5��|0ۈ�iz�0����_8' J�F\3,��)�+�xB�1�58w����`�?�_L���5 Hc��Ǔ��L��a1�j�;O>z���%���\6yw�����Qp������jt?�O��ܟ��j71���T�c-lRz8�,&�]<�/���гտ��Q�?����>���o�_|�۲�cv�!�I�����z��޽{�ѻ�oVdE��Ҋ�<|�%����)�;���K܃� �:)7$����K��!b����q� 1g�9�E�;�)W��*��ғ����Y�X�HZ�+���o���dk�jC��R)�l枂�Z ̰_?�o����OeL��y���x �F"���HnT����t��p�F���!/�{��`9���LĔ�ER�H��ܓ, �V����r�(f_�0�R$1�`��;,��y��� (���b^B��U��sU��L�hu�5�r�z!R:��V�.@�A(�j��޿w�� D�l�ʿݾu˜�p�|��g\�qB���q<�	�7�� s�Q��d�~��1����P�YV�"��]޶==�Y�8�U����g�{���-��{��{E��G����嗷�\�4e��X������N�!��׳t��t�_|��o_�re�&���;r�H��ȷUZV�7�
s�?�f�6Dsc�������FvФr�6�l�lg����)=l`��&�S�����ɩ�Z0*����m �6�LV3V&R�*���c\M}��20L�:�G���)�.�l�xk��{�5�)��J�����&1���4nj3#�H���o3v[j��{�ENZ?�����C��>W���IL��B���9�9�,��������	�6�� "s;��e}��0��b����/'�]��G\	�a���L�:����� ba>���)��Նj>��r.��&���ux��腾� %@=�%���	 ��0�:|���ٟ5 ����>̹kN�`��8���e]}^mD��i���O�ݢߋ�Rڌ}�6mؿ��t���[*�}M��>\��UV�:&�m���	\b���`�{����D�˽�{��9�q�K��[���h�����-,�.�q7M�Ń��ޣu����>�@����{�+��Yꛣ>WgΜy����.\�0kVdE�e�`���KR��B����pWr�@>���@݃:���d�;]���#�KE�@�Xnu=rà5�v3�-d�o'+5+�����?ex��6V��L�Y�J��"[:J4{9�^����ALv�^��[�j7��,��E/��8�Ѓ�oC�hݸ~�A&@
�d{�k8���GI����|Ԧ?0�`��"X��(�;�MВd�M�	'$��<��p�8��RQ�ܘ����p
�y!��n^}�5���H޹}�[��ƍf�~���_�v5�N c�)�	v�����:]O�;�lٰ�~fy��j]0�Σ��I���e�C���]r�ȱ�dy9�!�!|Z�`�%�X�-�2���x�9b���c���W�i�U4;��y�t��o�P�	-�ʧOyL�]�e�w��{����0������q�~��cǎ�v�F�=K���$��ݳg�kw������?�7+�"�0	0�x|���\��oG?C�GL�F  �b+����.Q~�`�PXi[qd%���]T�0�bm�uv��(��,��<�׉BR�EL��+����}ϲ2��[�D$�^3
�ﱊa��,�L[dC�,��6��6�z��������� LK����������_6��",x��k*uɱ Nꅣ?�`"�]ΪCu~r�(����I�#t���P]P����v�*���0�#w&�q���@)c�@����^#�:�K���{C�K� ��%�B{!���ݻ�[?��9~�8�ſ�m���s� Ͽ��y��7��/�l���Ǡ�4λ#����I������q2�7A2{!7��ImȌ��$Z��̑�^|�UN=�[��t�����6�v��꺒�ʎ�YD:�B���0��wA�������U�L��l4�}����=�^���"WW.�|Z�v�f�Q#}Z��>���3��c�Ӄ��/c�tZ�msl'mw���۷og Ic�nF}��?�яn���w�w�WdE���4��o<cd�Oz�K� *a+=�����L���f�b�f�gZ�?@�`'�t��T*2g;Ŝ���UiG#llP�}�p��g�|�=ì+�*�7�TE.��r��[���Y�F�5�K�zqԯ�$3V�j�"���HBr^� �͛`I�jl6�#�339�z4��F�ͅ�Z������}�J��(���4�C�j���I���4J\m(�N��Yt��5�o%��<x��&��x�~���`�O�:e>��3s��Y��S��NH���E$9"�e�	3�R��I�{�#Z�G$G[x�5��"�[����1�lԏ^�t�1f��@�>�c)�b0�ҡ��vk��ΆEϻ����)�`�b"{m���� �T�M�;��?N���0G���'�qn������_��Ii lgE�!}�MZv�9����OP���;Z�@:�+����$�}� 6��$4av�֭��wzfEV�k�� ��]%���(k����۳y]#�ބ��+�A>�EI�?V:'~��g�$��2s'0�R��Dt���v"�4)��ِ\�$s?3l��"�
���B���^�j��U���R�z���/�cN�nM�*$f%#�E:��Q0�����f�K�N��BQ��W�g��ڍ�z�z�FE�&\x��� ��L���������Pf�ku߼���*���@�|������}���ρuD�J��ٌ@��T���׭3[��8/	�т{��x�<w��D`g^�R��/��$_- +ƣ�X�6�c��ZXS��{>��o9��W�>̀ b�f?�Md8����|�,�\Hׄ�Sț�
?`���t�M��F_?�^�_ړ@P|��Ƙv�1�����&#~~D'���4��tN�`u��a��Ue?F�����Rw~dZ�R��@�A�[��5?i�_���֖$=y�s�$���	��w��
%D��_y�:�[�F. �kGc��ڜ������c�F�fZ����%�+0�`]�i�I�r��<I�_����s�7�u���w�;v�ĉ�͊���(��Vz\�՛#���GvO�	#���Lbv��aGc9�^�h�`�QIE���E��6�*J�C��&O�%
G|y���?���I(0��ɱ�G��?s��ǰ��z3\8�ϙi8=O�W/�h�2�/ux��gc��V[����>�sbb~�L��T�|rMpZ � f�D|?��ql��F�.�Gm_H���2X�� � ~ql�u 5���b���u@�c�tL�?��	��~�Qco��_'{)}ĵ��׿�5�L<t(F�#���Z���擏?f@�{gX\��+����[БS��/�����������,*��k���B�x�> L��f8C�Ntr<��]���~?<G�{��W��Lr�����1�F�Z�qQ�)0�K �hj�V�9�X�ҿ��u����r��֍u��u~��f��Z:�}�&���Ά�d���O�{��y���Jw�s ��i��7�|�K����l�Z �9cVL�+�d<�f�&��!%L_�>���1�Y?7Sk3��I�;1�{�(?c��lm�rJ��zY�do�
 32�.�$$s�*�bI=u��3�P����n�0UUh�O�x/�G����-Jd��MER�g���V���-w	�2�������u�q�S"0��lb=��X6������� X!��/l�"%���x�Lh�� Q��)/� ��� 0��?�	�`!@����:�����Lp8�}�6#�!��,�sX�(Y�� �|&$q�����:�����!��ܤh�����a�G��5�g`��F�"�α�CM_tI�^���.�{�&4��T����~�3TT�Ϟ��@:p6��jb0E��EHq �*��Гy�����q�a��3�a�J���M.�;��%�,��{!����{W%�|9��sJ�e9A����	(�	76�K�[m��6��;���~�& LD�_�m�FP���/$P����N��&�)f�Y�e�V �UɄkREq�6�� 83��ZRK�jo���o' Ǫ�>qU`&�悉�+ka�\ �R���2�Ѿ�hUf��Vm���p�GU(.���~��̢�A=l��^(E�^(0���� N2��Jjv֟��aj��>��zh#�+�݀Պ��g��v��s�Mb���;ؖ���7��  \;�E say ��c���U���X@	� c>��H2r �s+�#Lf)m�Ԩ��Ov�� ��>�� �{�9T�A���h˾S�ԇ���R|K�D�9�Z�TB���#Z�#į\��D`7�� ,�7�@ �S�ǲ��fgg��9����G�)>��7��I��̄ڒ� �)Ѻ��Κ8IŽ55�*�i��i	0E��7_n�{]�^����\JI�*�#�w!�z��39�� �d2yQ>܃)�|#��$�׃��
HG�L�]:�Z����w �9��0/����(�9��M�<K�9���?�H�̽��{3fEVd	Қ��GW�o�Ga�Z^`P6��,���N�TWq�=�	e�sN�C?���;�N{����}�g���B��bX�������bnD�Ǥ�$=R��l%W��L�xwa���ɶ����6��y���WviL点r$��߼��O*۩ئ|w���� 
��,�|��P��z�.y�&fѥ� ����f-4�C�� �8N�C`�V����׽���f>����\�1�h�6�F7����)��=����"��/����C��-����������h�\�j.�?oҵ�;��g�5����9��KB�~	�p\k��n޴�<x�]`.?�Q͵���b�b�;.�,2�-/�0�q˿��`�l����/���l��А����3Yi��;�_J����ͼ��x���Y���(Ɠ�tN�l���0�������& &|7�s=�7h�,�ۯ�;�%mz�ĉ��o�Y���`�/̱"�m'f�hjN�m61�����G]#����l�GX��E=�8��l�uf=H�Lc㨃$��K�UL�T�@���ב�J=�Ft�Ď?�r�ȶ��q�)'aZ?3�8&��ɧ*7�՚������Wg�.7��`�=��U�8`�>���V�77�l�����u�
�'"N! 0`��X8�x��:#�S���%���|L�Mik�	����ӧY��E�3JFvCB�&i2��2���L�f0
���,Q9	��#�s9�ͷ��OQф��`�S�N1 ��A����>�ob�0�@}�����B�%(�3�<M�{��4\����<� ��L�<Jb����LuX��ޏV1��#�D>�'���=]��T�k������d�@��^�+L�>���&e��L&�})��DVa��r����0�X.��9�qFY#t�Mϼ��D��Ӵl�)�������h�~�;�}��? �	���t�]������~둎Z�u�֣ӧOϙY�Ҟ��	X��}o
��ML9!�Qby��v�S4G/Q)��'�AN���9�<x��R�)��	�����\�b�P�p�>΅�L0EaU�/XĔ�A;�s�O����үB���`w�H�� �dnОI��'!�It�"I!4���1 �a?B�J��7ۙ�bP_F$�K0�o��Q�fX�=�e\*�:Jp�9����������K� �v߾}f�SOq���/�l�y���/�������HrNO���}��ӻ�f��6 ���L&F���3�Iqha���ɒ��u$�Rc����C&���
 f���\�?I�#V ���2�8.�,ۍ�Z���K��7S+��a.&_��/�~��'�vA�n���t'}��lN�CZ�>��o���=���|H:���Ǐ_�1���ͽ��;|˛fsEjdqQ������.��<}6G3�(������+�S��90�6�G
xK/��<�̘��%%gra_��kS��8j6�hp���<�8�P�%��.����y��f�"��?� ) ��hs�KbL̃)}�u�I��Z��i,�I�F%��'�dsj��2��~��1M��R�	0e}�&&x1p �m_�|��@*uo�q�i���L����7���a'"����b������uLN���ޜ�@������F�K�I|�h�����.��?��|���Pr% �LM�d�&��i	��B�v�R�t.�Ն'�`�jG[�i���
au���H��ٱĵFo+�]0�K�苲��ow_]:8��[��e��-62Z��+@Sũ���+�kk� ̨;����ɨOu�dB���8M�_�V�9p���V�#~�4~����a��M���Y}�6HۡT�mZw��?E���Ç�^{���r%�抔26���\���_�ߡ�R�BTd��d&���ŀ�Hɦ���C�}!%HƯwQa��go��-
H?d0%�����,�vM��Ux�!*]L^�F)2�p`�)�&����&�A�k 	�$���c�\%<Q� (���ħ��ur=�{ƅWA)�0I	׃�C6�-�i������$M@"�%�g׮]>����{����N��q�N0��KE�y���^  �TEHc$�ݣ�����q<����T|����V�h�9`��[�*L�#�'�@6�~�"��݌�>�[��Yl�M��Ͼz��=C�8��y��1aܣ}�2����mb	��7A�{��T�s��u�����s����uwC@�>z~����wh���K/ݠm�W�V���h�y��y����`&{��,^��g�8r_���筬T$7n螪T��e�/�Y�OJfi�4 'x0u�I��GS.�b�(O)���RS�N{!�ŮJQ�z�.@��D��.g0甹�(�%=M"���,���r0�A�����k�6;����.��
'��ug��S�泶 3~�� ��V���	��߰�YI��!�C�RH�D���؆�~�`ļ���lj�"��j�' =����k39p�|��wa��á=.n�B"}�َ���ʽg�v�a_r�(������;Y0���ͺk���>]az�k����_{�i}H�`�}��*Ɇ*蠤��^��Pȯ9���v�!�A��}?�ޥ�*��wA���B��T sX��7(�I�~��5��ж������VGD:�k�X>��
}?�z�곴���/�|�O>�k��v܊<1i_ɧ'��3�g&����9̹ ��~�k�W�{0��?,n�� �VR�}J�`�`��k�Y��%����Y��H$�7��	��`"w��|��|h3�R s��(�$R}.0��|�œ��F��RN-�Uk��F@$T��}B�Kv�( &|6�b�T9�N�L���
��i�q=���厧�b7D�?
���A|dc0����:�t?m��d��]io����Dxߎa��uЋ�P�e&2h%�,'L���7x�`>�Ɍ�u�ct�t��=\���8���,�Qr��i�_~�.� a1��o2��ז�'0g�߇���Q���)�a���>7�x�d�$��s��t�)��D��7�x�����Э[�*��W'N�?WՊ|�e4�ܳ��m��|9H`+'�/}��"�<�5�$]b���(�7��~��:��f	$Si6W0�c/d�;��*��\P�RXrn��Ƅy����օr<�{F��P�n�Y��tD�~��G��7֨ꎣX� �m*�W:�q�>;Y�žf�-���2chո�k�F��聂���
6_ݹ��<�ԃ?̫��L�3R X�=b�^�Ki��j�35����sW�M._~������s��Q�`��NJ&m���J�i�	 S\G���I[v��Ӿ���:�'�R��s�IU��ώO��l�������i�Q �v*���9Q���eV��,6����/+>֋�����)����.m� S��u���f�(��0���b�)��$��xF��pa���>�Ъ��	&�w`6��}@���g��������gV�FZ3�1-#-Ġ,�ϋ�&a�VRҘ��\Lnnr6A���!w��J%!��o&̢%�Qث�)�k`D�m� W�~pʌ�B���q�+3����X�ԏ��D0��8�j<�i����؉I��Znݲ��)Q�" F�V���7�[�¼
P�fݺ�x�ʕ'E��(�� �c������0qs\}�=s��is��uN��I���5I ���ta�j���N���d++E�{H+�^vl�7��nQ<!͸t%'&�! 3�ϔ���v �뺟K �2�f���� ��:�?WXb K�A/�b�Pi�)}�YAڜWS�G��a��&im�]���H�n�ljz~�y�ͭ��� ��ҕ���`;�>��޽{�z뭋4���޽;���ݗ�&r6{�H�:�N�K��yHa��U��k���P|�c@M��Pc3G�%�
�h�*3�X����w��B��8�M���D)�t�>�GAƌ��	%}"`_o]���>���d��Jq�0��N�Dhb#m��S�Ĕ�wa�-}��}�ۇIA�N�7�a"����>�S"?"ج���3���\I�	��#p�kS��;�SO=�,���4D��a�ô6J��c�>6�L�e'����S�7�.�$ `���A�q]��$�b;�w��.������T��7���</�) �*�n�׋.9�R�w-V;`��j�YF���, M��B�^\<�����k	�����%w����q��Q�p9���K�7� -���}���
��m�Ӥ����-�<M���'''��^��������/���J+��
���ҹ*.�)��S��C��Y��Z]�}����<(�~��}��bP�����&ӓ�/Ǎ�,�H�2��c�d���s�R���Ӕ���^'��˖S#eJ��2j~ik�n�mjs�s�6Cۊ`b��h�dUu�$c)�}�L��^NNM���5f�֭���:֫W�:д��ÿ�� ���z�/�oӋh9E( H0�pI�������<@�~�_YޯhG3��N37L�N8po�Ѐg�Y��6y�=�Ąk��	T�}�	'&oR���a���'�h.���o$l^U���rI]��[ �rln�ӉSl#W�����b�Ǒ�h�;�f' L��
qW�;��&���c9�d�{�I=��&�u�-�5Ǣ���&s��m|]�瓷�m`F�H��K�̟&�	3�C�ɏW�}��%������9%�e&#~u�H
�̠�E�z�!,"���/t�`�o |��߄U�Q��Div��4}�cW9s��\�B��p�������f�~
���Pb�:�_.�>����պ����e���m�Gնf5�>�������6B(�5�IE��_���<������̥K�\"��!`� �τ���'�la��u�A~ƹ��� �eE�^m���a��3�X�{�y3$IG�"���8`Ђ���AMx�a�Ll?���1o½U����W�j0���&�O�y��!?���ˮw� 3��5%�"N=�"*)�M��5>��kH���@Ung1Ѫ�S��I���W2ۃ�z ���X�`�ƒ�R3���QC┎���`�5Y�ۗ7m#�ۀ�aߟ����({.[�O���������'r�C��i�(I��+��r�O>ylF�!+�m�� �2��.���M$�����fL0'0�f�b���:iOC�B�M��8��ά�Mmh)M�aU��Z!�~����;�+��m������I���F��ԑ�٤+�>O�[�� ����o�r��A'��GC�u��n�2O$]�4Y��U��V��1�eD��x����s��L�cQ�/��I��Wq-g\b[ L���0�^�����C�`�}Z���~�my���,�Y��k�w�f�1k�#�姟|�� ����&�Cv��Zݺ�&�y:�`�dqY��dn ���F]�p�D�����l$��q"�S.F#�*tT(��M�\?�iu��~qVk� �eJA�e����D' LZ4�*N�4��) S��JFw��G&z�I���lWj���c�ɿ����4���Is ��B �?M�����o��Z����>}������|p�С�?��O�e�_�o����\0��U)(E���pf%�t�vi�+}�A>՚����J�8�����t(|q����g�L0i��8�A\<��Ze��
�����D��:�/AGّ+�j;�Ar�9g;�"�>�������� ��}�@������*���8�QU5�t�'�����{���qG�\'�z")l�m��"��/�؏��EeNF+�if�=?��l��]G��s�~�Go\��?n<�QRwT���ѝL��� f����
\�"ಛ@< &��5hO���I��<���p�di����|���.�x㲹0��e3}�H럢�o�r����-_^�x�ʱc�nМ#��.ފ|��E��=�t������S����r#u��L�X+�#%����+%���t7���^��l`I����?*6+$����F'��6����#�sk#I/d�#�@p�L0��2P.1��)�ä05TD�X�/�P���n��˒rp���~O��g���F���OwHd���ͦ�[��"��h��GH��G�������ͦM�8���MQ��
��a�@<�lư�,��6J9ą�	$�gL5�"����k#��eWx�	O}�L|�����s-�e7,	`Zf0+0rݞ�Nxs�d<����]4���	���H{�.M
k�Wi���x<� 륁�μ��s�S�~��gX|�O'�OAw�wB�]:g��9�a}Y�6�ȇ1�M��Y�,m�0M���mۯ�3]�	��iYO_	d���'p?O�%�d���gN�>}���^������>����CS[#xE��Ҋ�|�h���Ϙ����,E;�[OS0�����/�G(�J�C[�GS�-^6
��#`��O����U�!�̚�I��}}���-�����$`�m���bCJ�'͔}���2f�5+ֶ"mU��c3����}+����Ht2o�T�AD�#�����-(0���'m&�C
�\0�UTw)J&�`<[ȁ	�9L�m�Y�d��r �N7E8���^��!�ԩ&X�ul�9ր��I٨.���[*�����Ħk��� f$k�+`-;\�q��KHӑ���t�&�;�8P��E��sw�o�v����f��s\�<l�ךq�zFs-`4t����{��U��i�,��G�A���+)��2`"Hb͚�ff���2ȃ0�\iv,Ip3�J&Й?86ؕ����6��� X�6�xS=�`�R����pl�W?�����f S�H�*��3��r���� �_���ƥ��ے�4Z�����_��E���vr��W�.�i��/�\q�=R{V���>`A�X���XI� $��$!|/] �T��~�~��}�����ܰ���Rq�I���ڰ��|����lڮ��m���B ����k#��3 T��k����F(��%��T(i+lys����3?��FIf���	�U�	�^�CI��̻��"�>��l��C.�7j0Yw���묾�>ɱ��oh`�\�K��pJ'�m5ih0�,?�,��� @K]�1�r]������m��O`��S��&��)d\v�N���~���Hྃ��F�i7��i|��[t�Ђ��k�|��~��K/�tid~��y�<z��fK����[6����,oxhdǦr_^�Yn�W��f,[�W��i��_$6&V�bC{�N��N���� I�x����$L�\T���%�>��nF(r�B܂�A4�` oݺſ�E@�S��ֱ=�"������')㴯M�ee]&Oأn�;��Q@�I����
I�i��HJ�Y�f���"���9W&��v9�۩S�b`Z�-������s�:�T S܈x�쌪F����$ �~�Hg��6�&����	^�h��x�Ɩ��l00���.� 2;	�[���2eT��pm*�|]AlX)�q���}� S��uی���i�v\Y�X�'=�	۱���7�<�Hs4K��<�zM�rq�رk���J	�o��N�n��^�������u��':V��F�4ktw�s�o�F%��Lx�����H��.���uR�.C�2�p(�٢��q�A�T�}>��Dv�'���!]�r࡭}�������h?�k�U��m��{E��Ye�'M�P���i�@�O >�[6o�'�-+}���~���v�*G3�[[�F��Uн��~�@���#����9����}G
�)R�S��<����q>)8|cQ"R�X���\�����H�#py��~�@���t�Le/��X��Ā�����~s�|;�-�t��eXm���|��� �J��/��l�������]ct"?T>ݗ�����V(}��ɃUద��n���'L�,b;�h���3�(�lb-]`�%ќJg��N�����m��u�6�3.�Ҧ�Q���%`��i��u���;鳲�%0�0��c]�@��;����ٳ+%(���`r�p(�� /� ��4x�|2M��َ͔Pd\����\t|�a�-��$�*���к遐�l8���X\ ��]�qR}�؜�0�����+�X�c0.'�9�_j����a֜����Nt�/6J�h����D��ojY#�6L�۶m3���}O4��\XBpFc��'(0���#�|����S��l�O�e�%I�� � (��m"�M��Z�׬1ki���FX$���} ��H1C}���P�|�@�� �l��i{�O��s��)s��W�ƍ�;c�-J6t"�X)X�s8�ԠP��>��P�1�]gZ��)s�� �I��I������b�ۀہ���B�v)�)�D�3@8�(� �*��4��]��M�a0G�[����{1U�}���WB� �]�7(pz��N�K���7^|��/���;===��h~s�=�$�2�p��m�o�V�/M�{@dx㙨b�mS��F���A��I�K��v�+����?�2��	��E��4��,J�:�m�HJ�x��G�	�����Z��9M�\��Yj�q��� �j-$�Ɍ��e�#��ҋQ�_��;�����4������^�&\WI��O�wV�p�g�^^&�o���~㖒WpD�#�8��}�6���6	�@��-�7|N(���/�!�GT+�m�B	U�6Dʯ# Vw;�n��"�	�T1j���3��Tw�vz_ _ ˃�Ç��w�f ,��_Z��8W�K KN�O��I/s��EΩ9;���$h]'�.Ĕ�M�� {'�t"s���̊�$�A�~�~�E ��sz	L�M��`�+SiԵ͇$ץz|���eWM��)eV)�� �_�K���V�~���*7pki`׆�{X�ۦ�So״��z��7S� �N)���m u���m�?�h���#��U�<K���i�|���>~�������Y�?���^Y��S	ɝ	`��n\�Ⱥ�o��f0lȦ	�1a����e�8v;���׳�6�������d���#�;�����`j��(��2�J�"}l�g��] �o'�}������{�����{ęQ/&g�{֛⌰�$���H�H���~� 2O?�4�?���3xYn��  Q{�� �������<H��H�]�Hi�/���%��C�K �.�����p�L�O�A48��fO�c��갃�ݎO|0=kY.FW|�&�����KG�p�ȵ��T#�L�C�̡g�1�	c�Ξ>m��}�8�\&�Md�|ӱ�	��JQH:��F�8*��6�@ZMF�SK'��Ȳ�#A/.�>~B"�(z�-��o)�[>�q\�ݟO*h�Y��cɳ��YN�9.�ش~T;m f�[��c�춑�����\��D�G0����L.H�~�����s9F���{��.��~@�ev������J>��ٽ�3'�P���0F���M�n���6F�Bc��8�G�8�hf�W
8*�e:N2�h�gMb@Ebj�N'���ͳa��5YD�����Gl�]�:疸mL�2ӰF��:S���~��R�1h|V��M�H�f����)yy�K�X]l;�������_�:)o���2��0�U�L��2�Ev1U��B�o:�b&��W�^5�O�b�������t!@�~� ���sϙ�}��ܵˬ�;T!��Ь�zH� "B�/���-���~�l~�c#Z�.��nrїy��yj�N�,�?p� �&��0�a��:������~�C�N����͇���Ιk׮1��'��_��,�C����|��'�N��o�e^�����gsSLB?��Ssw�n#;�]$��tn���@�T'}�w*�������>���o�l���q�� ���� +�ݤ�r�6�&W��L�
�>�Z��Ynk�����!�;�^�%o"�<͹.}�૩�{Y�>NU�Q��`����F�W�V��5��Y'�th �������B� �ObмB��h�I��WH��z饗n�^yhV�k��L� n� �`�"js����u
�����^�}�fS^��&�ԀI�=_�%��~����y��qm )��/��4=�r^>�V|�2h�j��6�4��6G����$WM.�2��u3{�A�� ����+��ғ�  )L�`��a�V�|-D�T�={�kf��2�)!
 /KaR��[_��Z�?�����^x�#�KA�B�&��'��+W����|� V��O�:t�<s�0�޻�M�MR�"ҿ�5����~`��� ܿ���H�;	��l�~o$��m)��_���l�k��N��Y�)>��6�e��y�Iz��B��0�gZ'�f�$Y0
������K9�G�ڏ�����v�R��>>u��2����^_�`r�.��;6��M��v��)����9���V	��~����6c3�kk�d��:��|+]G�g������A͋�\���8}�ر�'N��m��F\��e4�D�}g����� Pō��?�͂=��˕�z�[v���n0&*
� ]�!��f~Eq
����=S{���T�G@J�N9B�c���2�wi�;�sU	�7�� �L��X᲏�z%M� ���,�b�:O��v'�$%>���\��4Lߖ��q<����	" S���~��E��j�"o+h���G}�&�_}Ł6 � �`�`��8�?��+W��!�/Olsp��� �<K��	b,@нk�.nw��w�ڗ��?���1�b���=r��y����Q,�4���}���p�>�d������:�pd<�'L� �OQ��t�p�pm1Vҟ�"U��o��%�	<4����h!�z������� La�0�3'l��{_598MM�����2 ���~����X��ŵB&49����T���%h�:���]a�de�v� e��(���&�9�xm lS��=��(Q�bD�O����Vo�u0�?K�EZ����}��W?'��u+ �k��L~2��4+��I��A�����;7>��Z�Z���TJiH������Tr��1L�k�[9�Ulf*�4���+�9�ˬ�����|��m��L�ed�����FL��"�;m���lѮPZ���{�ȁ8��n�Ɨ���z�I��dpr�F� �7y"xf����`��l��#�{�^�1�+�is5��П����A;�N�d`��g�1+ٽ{73v��<x������C ugϜ1gh�
0z���Qy/��
oХ��( 3�%:�=.��`V�^����bf��@���:����&k�7�&����/_6��<���f�}<.Z�̌٤��f8�| �gX�q�<p� ���)�}�	}|�?��A`WqN�0��Ο�1湎ۏ���YPN��)ϧ\����hd�Y>Wm f��n�!1U�M���\D���e���=��t�(�� �]�^Jy�$mv���3�Q��c<�o�֝O[0�ח�au��X������c�1�2�v�M`t؄�-3\�O8��0���>>M��>��i��N��o��w�Z�$j�2v9DئxC�i���j�(�R�	���:�m[��2�&e�L�f��cg�ǀ���W2��rl�+h8�{���o�6��A���V��T�s�p�Wퟤ,Ty���w1�|��+�hUa"�42�T�����j�Sq�)פ���|���!��b�G�m��O?����/� � ؿW${���K/E�FQ�`4�'�	p���sd4�#����l�_ ��!�R?��JIK%����fí[�P�/� ̴ ����~�g��������-���?7��W�: /��7�7��CD�b��df���~�����$p��>\�c	��Hz��4�s�`��pi�u������ϝ;�c0�����H�&h�Y>Zm*Yg�D��w�e����ڟn1 �d��tM1��ˤ[<�Ng�k:�DˎF��p}h�N�cJ�����$e1 ��mf�z}m�1�Z���r����-FB�0���D�p�W�3��/I�~I:�ڑ#Gf~򓟌z���"e$�r��b��0�@��� &���\w�!v'%�u��3N�>�,!n4z;qԖ�xH�T��G���6y8����=;vq�^D��c�5��e��EzF��(��6Z#�b#�)�kc��������g��
���@��	��j��OI��������$�vc(�&�ܫnڸ�K	"�@�0ڥ�M�`��M ,��O��R�~�@�O?����@L����3�;f����_#@\) TH����@�	�c�~�D`2ᧈ���B�$���֫�-{��Mf�����p^`�m�f֬���_Eog�O�7��<�x��I�3H}D@O��>|���Z�"���k ����¹̅$��|W��l�G[�8��� ���X��W�����=(&r7�ms�y]' ::���38`ʱ�f���FJ��)$��8���'%�9�۠Қ*�������m�]�:FL���C��EU�G����6k�[d����M���uft��EI�|�@c��l��{��X�9�@�I�gR�c�ԇ	�M����_&�r���&�|�}�����NϬȲJk��U.�*4�p�Ò̷xȑ�d���u]:\����fÌ߃?6�דյyîuLbƴ�?]E3I�.����d��W9Sjζ�y�v�̮s���W�}�EO ���bE�DX�oX�&��33��+�
/��1�~n��B�4|��|�^�{�yK�����7����~ۼy�8�t�	~���7ko�� �W���_��/`ݼu�Y?�/��Ԍ��8W�  ��| d�rʡu1]�/�� ���޽{� ���% ����$�8F�x��'	@�'��D(	��uR�a����q ���n\��n֘��_�˫v�8�r��]�S̺����+\��y�
`B����1X��)u��tNm) SO�e2���D]ZX�x;��<�_7�>�L���U���^���&Y4@
�wӲâ��x���)~\]_��Ձ�a�s��;
@J��8/Hl�q�m3~�VdR�k��.Zn��������s6��$��+��r��O>A^�����k��&���(u�*�Uy���0Y�~Z�e�g�3[�B�} O2i�`�z��"�*����lc��t.�����V&*"}�N�
l������B1�J�{��^(��pn�0�x�0\��{�.���0~��2<��Cg��n�,��4ۤ�׳<nq<}|����1P��V����D+��Z�Ҟ��g�� �YZ��2*Ϊ��p J17�:` ���ӧ͇'N�y��{�ۑ�����8
\j��(L���Q����f(��30��a��� �|+BN��k� ��^�#��M&�:�<r�o`����1�E�N����N�X�ь~���`w<�QW*N�N�/}�><AU,�t� ��/����1��l����a�|6�R�1(W���D�@��B���
�伴.p��bP�DM�6R%'���`61jr��tJ���ݯ"�n�Y����m�?]�j��w��гS�~踦rK^�y�����i:6�G�����-Y���U�Hg�(����,?���@��%�E[?l��ʨw��N��@`�w��(;�T�����;NҺ/HW�[IҾ|�(L��T5(�:(��U~�Xs�Uj���6+ڔ><�Մ�U�!���q^|55�e�g�X�������/��Lf!�`
��\@f���0��",��?��׆�FJ�4����X��$h���ŋ9�>���p�l�9��	HB�J0f���m�A��$�K��������\<t(kG����P��({�  ������$"0���RT�ٳ��,� .�<��30�5L	�@�L�0G���{||���~�i�#�w\qF�?��	�3S��UV�+��ADO�����Q�05jL��
V���dI~��Hyn�}�m�) �ǧG:��`�
`.]���r)&�a����̒���qU�Gw��ի��lذ��C����W�?�����ٳ�jhF�Im�D��~� �I� 0C��E1E�o�L�v��tW��q5�L'��SmX�6�����`���1kƯ�$l�t|���߀%\�g�p�.�@:�>|���������_��_}�_�OXZLzl��C�J�z�� 1��1�Q`��l21�VXH�]��3�x����#�R	�H�(7�:�?R�Q��"�~�
(ss!	��0�K_����t�a *�1zڃP��ea���#V����� �Ah���I?���E)��#��f����P��q�:�@��3i�XRѪ?����s�|'f�ҏ�Jd����}�m�6_ ����ޚ�������rFe�a�O�ݸy�#�/���pP|:K���q,,��iP0�fn ���rD�#��j��7�4/ ���S�g���$����M�X��ȱ�����l���0�-��zv�ﭑ[t��w��H�����
`�6F�ǻ��T�x�t�l���h�X�����>Zm�&T�=�M;�i#��ԣIo� f�!������'_s���d{�~p]X����_U=��{]_�����X�昣��NLL^=x���?���% a~���;1>��;fjWV�Zu����g�󵲩Kv��㘈\�6� �����y�x&sB��F��l'�ա�����t��� P���0���D��a��N�N���+��wf4��f�M�4G�hB�ku��������J���e�*����ܴ�|%�[ `��)�*8���ٍ�L�,��[���������t�O�.�|<��;�J��*yT|蓼,�r�ܒ2��ELHج��_�]��o�h�ȓ;Sg&'&͚�5��#b�$����)�~�b*i.7��8@)|=��յ�a��h�?�!�ǚ�Np��~�!��#W&XP��%z�Y<��[��K��Pߛ�+F.  �87D�cA�|?�[:�}���g�ƍ��:`����(��-����D���F>P�H ��A]ȫ���E��I?[�JQ�[}�"agM8_�}_:�����]q0��c����8cҼm��˱� �#2^Ǻ�k=XNA��vJST���)�.Фn����=>z��b��c����=z���cOS�+	|<�<N��N��2-�в�v�
�U@�8Q���:�#3.�#fn����C��M�M���,�e�����z���T��oA[`��q\M�w��^���J���1{���e��f�)�ȅ�+FT;)�&`˄�E��3+�y�,>P��qy���z�|0%*��+�O�_)��'��^��ӊD�k 
���6��&�I飜_h�U�c����R*�Fv&?��҃ns�G��k��2$М�(�ԾV���h��6�Hs#�k��˵��u�8�c����7�^�u�q�_���]��N?$,&@%���XN�<Ɍ�H�鼟�ݐ?/;�T���L&jl�u�%'%��}�N0���׾^�s���M��6������ce�6r`@l�o�@���Q]l/�bܷ��! �0�|�(�iBJ"D�#b�n|!����);��ٷ���8c<y̐���y��	�lz*$�[Sh�\O�����!��eݶ:��'�_�쾖`����K�A�8!���od	�� fv��#Q�W���T�<��H�.~�����R� ����d�u���M�X�y�&��)x��*�~I��-��y�#�#h���V�o��O�����0}�b}Ś0fy�����J�1��Q�E������g�d�\�们߉%`Uc�-׍���u��a�\K�4��5urzz������֭�y�ĉ+ sLi0y�'<�{�8�*?��i?��dH$8c��9�\�ڰ\.���RRj�lm6��b�G�ۼ������e@��x��#p��x\8�7��hz�9�j�J��R��I�w�榬qE��_�&�7�]��9y$9��ߏY��$�� ������{� Ϩ~�%D4χ|�̮!��a�}���zHɋ���0)�!e,z��5��4�`?��(m�L6 r%�� N��6AQe�R�c�Z���hr #ρ 3���;82�@��b]_ :m�I�QF��>p萹H��XB���!+��	���X9���	�lSr^>Ǫ7yý���6�&n>u���q�N=���� M�`� ��)e��f�8���\}R��֭�$6�p�&�(U6;��D�����W��]�C���e��	��u��N��S �=���.�&0���s*��p��hAT�����va݀(A��% ���u����ϵ�W�����X(���� �g;��ӫ�۱�^z����G���O�0+2��� 1��h����ȋ���c�Q�s��c`�MTx+g0+ł&@(\a�/�^���ȶ3�{��Grپ��H���m&�#����Mdxc�}%e6M�Ol�B�fs0UP�ڼ6�xv�HO֙\���L�����˚�a�t9�*��f��-�f/�AS`����d�؏�`�-�@� �nظ�sa��ƫ�Y�*�Є�`�p�9:֚�t#�Nm��IX��LLNpP��վ>��d$.�E*��!�;:��.����k(U)���< C9>XC�_m+�0^`/ĄtG��G�<�KYO9�M���_��|�L<[�<`�,�t��4WB�/9�Q��B���k�x2 Ϫ�u ��%�4���l�y���Js#Ǎ�->[� ب�9izr�#��뚾��Kic�+zkkE�zv�'�Uҏ7-�{У� ���S.��\�J &�-�/*�y��n�$��k���[q�n��ی��ܡk���v>�[0���������;�j	ہ�C���(���,� <�&k����6@���\��&���u�w�uWѷ��S����1��?��������o��Y�1eQQ�.[C� �b&���mg�8o�fS���M�T�iV�A�)�X�f�����$"2����2�x�w'��!UX?�g5ƙA���80�q��4>ݖ 3*���UR�^"��׮]��s>�u뢩T�R��ܡ�fH�= �(Ae�9��U�e����c�`@
`V��w	D��b+!3�%��L�z�?'�QA{��)^&<�\�b\0n8�D���B�:�!Q�3v5�sĸ��D�"�ADH����iA�<����3��O?���i���@u2��Ă�@(���J��q.�_��������d�L�3���z�~&t"���'���.G�<��+��&�#[hX������dĴ�T��"NNS>e��fr�W8�VMֶ�]��q@����������Z0�tn�� ?���e'�;�'���|pA0[���q�5�_qЄh�VF�7��hi�=,�ڗ�����;��]�?����;�Z3q�ԑ����"��� 3�BG`�����S��_�Yg�ZQt^I��M4�=�v����)Ѻ��*�AK<-: x�id_�ѩ�Ǩz䮊�R�T^2����%;�v��On�Ih��_t�%��-�`��63��rJ��b=�vͻ�_<�WU ��� �I�W���Y(7�
���	�ph��;69��`�L�1��O��c��<M�x���uA8 X`�S�c	�YA�iPo�	��_
��b��1ͯ�������Ă>�`�>!�� ��~�x����	�"*��u�K����ĂR�`+Q���+W�CjG��Q)�6n�`������xG� �'���R���m��:"h��cvf��!�/G�~���!�ha�=�ܹ�=�����Ä�F�kܝ�e���C?������N�\_.<��U%:$�G�V>G��u��?(9��Y��G�e���`�.�[tNP,P �~��i�]��@ߟ�O��3��aBd:Dƥ�5,�$w��v[�h[w�QRN��zi��O��d�ݮ{�m�����N}�ck����vO���Ms�����֣-�����[�1`E�}%��W&��HzG��BB*}��`�_	S5� ��2G�&�@4�]�������vA";�|�zM�\���b ��VlZ�>D"VuZ����8f���|R��Fz��� ��geF��L�׀m�o��7�w\#��yI]��Ш�y�`�P�:�Ĉ4�
>��f�n��9z� L���+}a:G�I>Tz���)Ct5�U>��#N�TLa��R��C���`r� h!�k���=�9��^kN*�I}>e�0�#�B�cw��%�A �r�a"f_�������7�1~�R{kiBp'��� $�_z������ᇜ���D� �q��!�[�J��h�^���16�o!�F�6���f<?�������k)>�ggOß��Su��o7�O���~pΦ&�?yP���F|7A�
�D�8y�q"���%�a�z��p���oU�ʡ	��G�-�	�y��0�_��Q��)Z���_��?C�|4���勵Q��sDOg�f�mzv5��-`���zt��4!l:7l��Κ�f��C����z�|��隍�0)�	��u��fn���n�̇���{�l|m�\�f���ٝ;���v{�=����N]�y�W+Q�#&8x�������NQ�*UJ���˷��80�
���Qr_
x�L0� ƫ��^dEH�����(�H
%�<G�S�_��9�I���S(�N�H�z�>�w�s�S%�w��A��b��D�3�}�0����0%j�?ܨժ�ь5�]���.f�AG���BJ+�X�C$�����A��-[�2H����0��r=�-��f�0Y���IE�?�T��-���͎��즘��, ���X*X�{Py���A�/������R#u��;~� �'N�`������ѣt74�aj	`�36 )���	�������IL\>�1��/�?�ƀ $�[W�q X�O�<��U�P� �Ak��Rt�K�bf=3���lb�&30���ҏn������ ��5ݓu*@ ��ڕ����&�4�i�u�@0 �&�~���/p�J�2M��cg��TU0�W����5t	`��r!"x;c����Q04+@!_��u����_H,>Ec�������Dr�u�`=�5wV�ʍT%��؀:�QgRhb�ۂ�&�S�0�S3�u�o9ֻ���w���3�֬ro���sv��c�X;�9��3?w�Wto��QϬ2��L۹k'֮7f�ḱ��8��i�r��s�nx��#��&)e�i;2y1�ăoe6쒹�+�������ʛ����a��X�m�d^g0:����^�包M�q;e����G'E3� G@5βnN�(�*0���{�-��M߆���S�&XbRL�e!(x9?��c2u�/A����*[,�!o�0���;W���FV���A�Ɖ�
�ь�rL��b|���Q �D�㞘��Q�[��*��N��V b�ޤ�R
�d��q�������R˰;U$�����_���"@��o�i�;f�޽{Q���3|"��>���;��:��s���&�rvD1M��1^׮\a�8"Ñ�	�� � ��N�D�!\�\�l�D(��\�`!T?�D�"��Gnw��9��Yf��Ҫ�� �g�9��Lc���2�4�)���_�/��ͽ�0J.a|<'�V�̨��y{��y����0{��5���׿#�×�4]x�x��Y��sA�,�A��ʪ��~K�䋓y����ϻt���%MD1K�D�U�K%�s;���A㓿Ç��,&G'j�(ߛ��6 R��l��8�6e_ �"��>��ؖ!=3i�lZE�Tw�ZK�d~�ף�����{��={f_����&�9�묚7]��]��u�R����sv
7�%׿���/������3�TZ����AƩ��.>�}ӵ65Kx�#�~)J:ۮߋ�I5m��%�Kb&3EE3s�(,�Ԯ_E�M��8��M|2��idr��Q��F^��׽�K������D�(��q�<�����6rSRI	���	���GQ��>>D '��|>���4d�F�Ϙ���C��nx��=`���c ��$� �oP40��Ŝg&�o>��3������3`��,ݺ`����=;���!|����?C@v���{|�ǰ���+r�O�2�L@��~�����[o��ɟpya��c�h�3�4V����5��`������`Cu�҂=�8K���?�O�Iy�1~�i�j�̜���<1z�)��9�H�8��k�>
�N�`��f/�r| `0�L�XL��=7��[X���Wa��	�c���`b�`�<��% H�������k�f��M��L
��p~k��:�R�>ȧ��C�\�'����&����M������s_�nZV���s�˟����?�A��D�w0%H(1��z�	hB���Q�3�I�I�~��N���ի��cr�N���ىk���>=��뻩��3;Iqp��f��^���f�3ۡ��<���j�fr��m�{��߼b6��_� �F�Cӡ��������s�l=k��)�����[���ub����%s�	k(�N�8��rI1 ��"rc/�E�g��i��W[3��� S�q���y_-�v
*����l�hH�1ѝ��J؛� Bx�m�x��,Hq��L�I���q�%��;��4�����N����#3�\ꋼؼ��\���T�R�d���F҃��R���ߠ�gV^��M\;0J�'$�e��_�����cja�i@���/�4���*���J�	`t��i���X3
�%WZ��,V�9��G	J���`$�g��?����o~�&i �z��-�����xu�(/|������s�q������oݺ��~''�ǵ�M@��?MO���۷ٍ ��ᖠ��Eu��)0��'�
�;2�Ϛh��j?2���c�	���0�l)�ĕ'�d�x�eE|��<�/�ⓔ�\��oݩI0�9��D����y�ܧhn��,`���fa����He*%��	�"'�R�|�ڵk��~�����A���f�<��h|�os}��e=���>��9�~G9�X�R����Rg�n2�7�6T�q��;��ȥ�n��L�s�_u������M�:�k��L�s�u/�DoMw���۹g��8@�����tC�|�G/�K�"9g̚}�w��f����{�v��s���O��>a�wX�����ͮ4@)Kmۮ��Ra�*	�U0x3
��m��F�R�l' �d0�5�I[Oܮ�3��T�5)�E/����Vl������2U8J��.A��8�J(�R�	.��`6uRb�,x1��)��Ǳ��Kt�H��G�Q�� '�����y�gY����	?H$Yxs,����1`+H]�ܚX~��l
�' @ݳ�>k�������8�u*����6P��5�(�/DXk��5�܏�AKe��F�� {��䈄�"��W�G�\�~�=G} �<��9>9��״�$�'�٣G�2+� )\�����=f�v=��8x�}��UH5�*��D�w c �O>����XL�@)��Y�f�Y�O� z`)��c���:%��MM�4��2ϲ�� r�Kxj Ѕɯ0��Sf����f�)�	+X���9F��v� ��mr��(�EINH���Uv���|W��"��%@N:��lٲ���u�}0�O�|>99��~�h|YK0���hZ�	e*��F��I�y�\�vJЩ���h�A�-%YL$D���W�E��x8��3�ٲ�ƪɽ����M�����Ě7�z ���<�`��-��&�n��~d�,�j�~�6f�)�����&]�?s��/�>=q������O=����g������ j�I@��U�<�B�f�0<���|}8���2)GYP4�~A�At�ed 3��;��Ԡ0)�^����a��8��d��F�����dJ�8���9vB�d	�=i���y��L��S��~<��M�$�/Č���V��� �~`M�ť��ULf᧙�Sy	��Ͱ��\gLF_U��^�Ƚ%~W�O@��x��Y����W0hS�D�*̴��~�%��K{�]�F��_x���O���J"� ��SC0���8Ƈ� ]�b��q�C�P����3ZW�fb0�X �qLT�i#lm~ƈ�FM\�|���}8r�<G�;ȕ�n����8�����}��3�x�����:JU޸�K�w\��� ǵ�}��^|Ѭ���BH}�%-M���3�\�|���*�	�rf�i��s�E
\�$�M/Do�i���1�d�o�hUܖ�&Qp{༪S�<�\��#"��ٹY����?:�����7�=�d�={)H�P~9w{U�,���wV�ܹS���Ȑ�D��/��!ߦ���￹	�������j)�iS������$=7Ռq�41��W��>p����O��C3f��T͝�_7N?��vb����Ո �j�(翤� ���k��uZ&s�Z�Xgm�͉���Y���?����~���}��y�����}{��5�qiGC�����я %���� 'úS��N#!>n�h��LS�z5��ͫ�\;�/3�j")�8s-���`͊
��U�c_�1ߎ_�G�{�jy{���x߿�w�wi�&"Q���. �(����
���h��N�.�F�	0u;���r�Wy�hNlXL�}�j��L�"d�U{%�3��@&L�`3� ��"�ݻ{��)L���h��޼iS�"��]���pl��k�)���P.�jE����`B�K0� �H��"��	� /W�M N��Mm���G����{�Y^��`��0�c����������h;\��_|�S<K�-+���ň�:�R|�.I�AM S������eNy	����&���@8�w�ܾ�4kک������][$k1:�	`ց�`z}�2W�JͬW�I4��JC��|H��k�w��X��>��A�����&���V�o$���>��`�M�G��"<��N��D��u:������Nu~QY���˫N�;��;�����7泿3w_��O�5;ߧӣ����s�`;薂��c"ma޺�|��&���_K���g�=�-��s��+�ts���v��%�@�B6Q�c1c�`��'�^��0x�^�%z��l�̳���qX�fHO��m!���E�%u�};�O�������uvթs�8�T}OU�ڵ�j�o�]̩m�v��� �QڧZN�6��r���C]d�<�x�ɭv�e(mZ����]G[�U�܉Nټp#�V�t��P�`ۂ��v�6��s/��>�5n=5���?�e�V|�5��?t;���8wHP�1��hK�1Gʓ�$� �|}j.r��w;���1=��c�-2i���������4"���Bl>'C�D�%y�3��`",w
����p@�D L>�R�S�/Yp����na{��n� \E�{v���l;J�ur�ġ
�m�(�Zz	�&�n ��(2��p? �ؤ�4�`_E��,����벞;NR��`���m1_��.x�Tⳣ� �w�w:ڇ"�C��jl��J<��Q�4������a�&xƄG/��ZR�j".&�U�XN���A)��K��4~;��0֨zm��R��e���+�)�)�;���"b��!�a��vą��D���3���P�P$"�C�c�r�I�QDpY�x<����-�!ay�~�l�x&�/�x���1�)��td5��"J�-�x�}�|��v�77��q��s�:q�F��YZ�l��HY ��� U�+Q�#�'O�u�N��l������^H��~S�O�+���Q�����8�g(վ�l�i�.��cְB��D�z['��?�P�G!�]��n��ˣq;�ҩ3j��[	M����*)����y�fƢ�}_f�џ��;Q#/3i� &�9,ب���;���� Z�2��Kh�n^!�5.��|���ؙ1��O0��Oc��OJl��-�&��9�ud�#� &/�-|������*�����c�����G� ^� �b y9��2��Aei�o`֭\����݌<"@�蘰�k@o���z"S�9��/]��Qe�6�eώA��?���p�� ��#`D�1�V��رc�a:�+�/�5����	��葍+� K�a�� �!��_!=� �5/D���?���<�}WS���#����^Peϗ���l-2�h���Ȁ����v>�l��A�C�cm�6�_�a��ͣMԗ6��<�y���z f���$��{1��+!#�u5]�KΕ9<�R"��&Db���ܼ� suu�k�*�#w,�4��$��	�٦ ;bB=)����Ϙ��;ucl^�s�y����y>
w�1�b������a5�2����`�*j���C#�!�����-���m7�z���و�B]޺�ر-�=��z�6�pG��6�L����dTV��-q���*�u��A[I�����a썫�јV��Բ�̲����6槈:r!��gGo���1��SPƗ��|��i}��v5.x3}6/�(㪳��b� 3����ٞ�HJ'�;R`]��U5B5�`�Л��!u +;��=�`0�>R:~_w�# �!�F@y~>�ԗ+�V�� ��ac�8�Ѡ&�W����_�c�����icLH���@2n�e{uD݋�W<;�dJ&?L�fr�����j�5�G�0��[GGI������,�����J:�!��*�<�h�XbZ�X�>u�LMNz��Ed>��`C��|f?W��P<� �e���>�{1I���}��~�+��\,���hn�τ��1,Q�'z�#PE����}�2�l���k�,��g\�.UV����60E_)&��k����څ���;�D3��S�z��z\ࠓe}����p�#?���;��,�ەk�Ԥ1 |�r����ε��S�0&}Vw(S9��z]�T� �5
��l�Ч��-Nû�U����<�%*���a�F��Rw� 7�Pf#�X�fjs�[>�2=l�x{abg�B社��N��/�%��O�h���>1ih������
Y|d)_�L���QwlSc��C�[a��m���X��0��A՞�aؙ2��yG~.�eG���^p��uN��@^&�*�DV�~��z�3��Ϧ>�*mߋ�`�r�I�EZӮ�u�j:��8�6J�g�qϘpy2?��b���>�i��2q�NL`P*r+X�:{��H �cO	q��ӧ�Xޒ4x���^~�����\\���6�sf���P�J�����DC=��Y�D�G?lBe���*m$h��4�!VyLV3��*M|��N��Lz6���}g��8���㉆�#���L�<�蘃f  �6��C&�0�����c�]#�:�����k�S�x��5&�m��(��36'���RQ!�r�����^{Fq*��td/�������"lӅ���>Rd��)�7�d��B3a������ݯ��8)��IՑ�
�an�	��)��"J��}j�X����i
���18������N.���nݍRw���l��c�@I��n�*�S�>E�ۡ�Ǝ���j5k��G�W%�s��s�e8��֊ �ce/�o��{�+������L:N���m	%�D�s���81/Ǔf~�bL*�=����k��A�������?x�S��率;]Y`�����$����P�^��z�UY��(A�>�t��k���Ag.u;J� $f²9��"@�k�iW�.��U�����r���	fҖ�/*�Mg�F���c&��yB�Mi0~��y�2)5|>t����*���Q7%�
�����2��	�A撅N6P��9O�,��P��:��6"���LD������Z�&�ݴ��C�BO�[-up`��E���`l�!T�u�E�x��-��Ԥ��������,1^d%���@��}�}�o��Q�m�섅�`H&�DG�c_�*sn�,"1H����.��W�5�u��������DL1av��ޭ0d��k`��A�HJ���MJ$��E��umL�rj��p􉂤�َn5�)���#!⛠���u�p �n*ؑ��1�Tږ������q�nqt3|;\�W�
�_|�N���\�G�q.|�|̦2)I���4���'�DH�@�t���r�N;j���y�.����������7�O����t���B����v��w�.������$�]J2c�@�=��nV�dL7�]������/���Dl��r�c7�mf�*rd��m�r$�G�� �[��s;EH�:*�Cz�����a]t�{�k2���E���$u��o,�н��E�*z�:�`d��Yd�LE�V���g�NV�M�|��a}�sT�
{+ *hI� ����*�x�׋����-�)�?�L� ̼��]%Y��i%�_αT����gv���z��%�ET+�m*�v���t�������A�	U��++|2���(��H s��_��Ϳ�l��D��Mp'�^�a$�� ꛭ���y�U9�s��`^M�?b2���kv�dޑ\Ӵ<�S�n��F����4�dJ S�{�*��`����0[�WS��r�(��5��ۛ����Oz`sl2����=pIJԻ��$$r=��({ݨj��z����ϹI���kVܨY�ŕ��F!���\a�]f�L���|��ӵ���/��P�	��&��T,���ۉK��;JH�>x[ㄤ�V�Qh,ەb���J�ד�����R�$�U��/���:x�Ho@O�U&��CI�߿i[�0�����+�4pDf;�� e�����e`�2&.�6�.���w�R:����4F�R��[���XK�ֱ�{�y�H��l(�&��U�"�w����I��h'Ǉ����� 
r�JB�3��y᫶�(��QS.x(��i�֣� xv��~`=ǥ:q?����:pcDS5��&1�Lp� t��X��(��b��>ǝ��c���� )O
���r�&�X�܂��A+�پ�P��_]60Ó]ה�����o���R�r�)�҉��V�@v-X�ՙL���|�k���
��W�`3�״��UU���|>�����V`���1�&l�໣�|s��D�)P_�o٬���&�o��q�Z�Sԅ������JJ�����N��g��[H�!��0��[��͉%�h�5����g��v��op⢐t����%x�5R���2��msN�x��n���m�b�$���Ye�N?C���}�o3/~f�|�6w*�}��;?b�D�f0U]g*�TwBXr"�Hp�,�$zK*���W'�;\�JF0F�@�$/%(:fw�p�<9��8D^�ڝ�0����@3�S��P�/�Ʉ
�˓I� EL�QWq �<�!��`~8�S���ōy����V�G2;R`C���`�a�x5Y8��᳛f�v�9Ÿ~	�͙d?A�K�`�7�F�z`��z�s�"�q�Q�qR��lq�51q��y���<&���/]�!��Pbx$s5�o>�
����y�rU`@'	��	����c��'jJ0z���4��)�\�<��tY�RnwT؜��Q�nҁ�A ,�L����o�g�L1�d^a�B�Y8�1�a�� Y�[��a�T�~����S�0��%��y���@���C��P��z��m�#�(M���htQea'�Nݢ�w����P��۽�N�o'�̭z�<ꔫ
��Qhg��ɮ�xW�3�:�x�/>��#�G���nu*�T�g���0G�I��R��R���L�،�(}C�R��u�m����rB͗_M���v��`c�����-�Y�#7��a�HG��)��x�zG0tN0�̠ E�#��n���kk��F3�x
ՇpꩫBꝜ_Q�m6�pG�w�IH0O���E�.o�`
 ,��:�P=�N",o,,��ll���u�g��|�L���+.3Z�M�%�W��UW�o6|� K!�	�O�AQ|0�d6�\�H6�!C��|�"m$��x�N�J,v�8	�w��F�xW5l����9��Ž��p���L	C&���G�ΐ4l��N�<����ѡ���V�&���j�ﷱ_[�m�PI��:;�;��Q$��^cS�d��ex�DQ/,�ۿ���@q#�K��3��j�g&^��m�3wu T��m;�����x���>�kT�#�(JEq�������<��dL[�sb��;����--�L��#��٭V&;�
���p�R�:�ؐ���~���O>���y	�^s��{�2{���t �P5R��Vy�i���1%�=Es�J��v��r�U�jk�)F�6�$�g�Hu�8�_�t��_��\���U& '�LR��{a�����W��N �$���FU��"w|�0���0��8�W�q�zd�T��VF<8g;��T\���r���v���Y� ��L��M ��n�"�Ն�~ ���]���z�yW�'�x�J��P_��N棕������t>ꘗOX��
� <ȹ}�`eĻ���M ��^xv�#�&KzΈ��I�jr=0��{�R����m�B&A!�IJz�삡���m Y+t���an��|��e�y/�`��:��`���I9���k�"Ll�0�ۧս�HW���{��a�|���1^��W�G���$�As�pq[r���=�@�<ھ㺩A�t���� �UZ�ײj�{� ��T�Ap�pf���eT�5�ϳ�ޖMJs�<�H\^�d29�S�� c�L�~\�o4m����[Z�>�Ė��9j&�m��*��P�b�R'3C��_�-��.TX\+�k�t���'���@텥X�X��7�tw%I2	���)���l���씎B{'E��ع�J&�? _��r7]I��:�{�Z3��X�3+�+c����1sDq�]�.�8f��hAl�a�\�ڿfO��t��{�u��*�\ZZr��ƨ�8h+�*E�ϟ]۾m�ۡ��y�P�rl�oI���5�.�֗�� S0Ri]'�F�1̊��\�����4'޾���9�����B��������A4�BP��y�I}Y<��'�n{�D�Tl0��\y�X~���<QX�%���%�C.�L6�m�q�ȉ�	�n\����?	�~!�ά��m���SC���Q�d*5��Ꚇ	VY�}0����d�����A��v����3�p��G�aWB���O$]9����B�*L" &� ��K���+��t,�
=Q��EG��� h" �c�v�f�0NA{EFn�����6�I[l�����F؊�Y��øxY!�>�+/�O��)�;�C*���rho_덶u�8�)/�&��9�T.ﱋe��Q�R�)�O�'���oΐS�lz��kg3�QyIN�ǽ���L��b��a�<]`���
;���NZ(��{{R�L����w*]�ֽ��\a����|������\`vww�J����L���P����ɹ`MW=�u��	m&i]�,��p��Ȫ���a8O�:��-*u���� R"���z\i����%�!�����;(O\���)qo`�OhiA\U[a \?'�0y`m���M��<4�4�Z�O���u"�T��9�λ��3����#��]/���J\&>�`�=���V3��;">k�?�x\>�[����땍��w����>_�s�)0=�TB�q��$�Q�+ښh���_��x�T����G0��h=�~O�C�(N�Z�k}~0�mޫ���*V*�\ݶ}<���e���r�����UT}��!P��B;�S�n��ne���sI�R�50��J  _�IDAT$��o��D8!B���ǨR3���wD��OK��ɔ���^�-�_d��K<�kB�o�}�P���p����1� �<��j�r�y}n�8���<L4���#�Ć���N�3 u(�Z�/"QȚ@�\,;���bdd䅮������w��u++&Uu�&
�0���Ć	�9F���%��Y��dƜ`�R��J�)+��~�Ԥ2<�u��Y��l��r[�3�̗�.fu�E���F�q�G̪q(��l#s�B�!�n�R;�`R������{1{��Ү��M+�FeU��e�L��B�d&�6 �e���4U���������U��P>[��Rn7<O"���*�2�+K`%QT).��!��U��O�ӆ�m�@l8\���t*�:�-�1#(�6L8��˨:���%T��2�"�����4U_�Uk�Q}>�x^�pEL<���<�
TW��T��w���<J�8�"\�̖ኮ'��g���ײ�Q0Ŗ�y��M��״�U°t�z�D<Ld0q�x�����Ҡ*�s�q2�=��K��<42�2Mo�vD��ڊ�����}PU��K=Ħ�Ԋ�����;�n;�����T��ɓ��\Y��Nyh*l�
�T�W2%��l/Z  �8��.�}�7;n'l%ǡ+)g�Є���`0���\��W���wC�9�y	:�I�#c�A:r=	�ф���u_q������s���'�#P���}.�6����d29��g;w�|�����z�i�n1�/W��+��i��i����ٵ��1f�{~���6ݴv��"�fT�a�f*q>��5c�bl*{9;շ�/Gq��	� a&��o�H�m3f��:�I�8U��ɘm�t��^�h�6Cl�U���־�ȟ-$�f�r��������5�L�
0S��R(�\��G��]��x">�Qe�V���7`KG���J~��{�Æj_��I%SĆW�A.+vuu�Z��)�� ����l&ƥ�(�r�(Բ.��\���:s1]��̹�a�0�)rlgܴOV����g J�Jt��}�E�;�\�CU�Y �g���&��w��P��z�O�0�[��p��e�]��E�u���p�E���LD�낔��5��zj��roT�½�Hi|����.�P�����`Av���l��P��-R�L�l�}����Z�d!���!���3��k'MԳ��&�6��YQ�۽_�tkaR���DU�{��!C##<H:Kǵ�����\��%�K\�g~c{�:�+���cab~�T���l���uU.�O�|	A���6���]�)�_XS!�6\�A�=�dWb~ǁS���/~�lnn�&���n��t�Z����|ZE��1���$\Jy��wb�"��҆���We���P&�F�/��̕�')H��OA��p�g���r�<w�ȑ����IG�;1dN(D{Y�~���n�߷�o�8��|�2<q�&������}��]������o��E�Քd�`,W���Պ�*��E�U�ZaTUԵ��YCoMJ�kӳ;���YZt��8۶N�R�s���/��g!���z|�"��%/~��9�X�/gT��e?1�7�dF'F���)���I��{��|�^� �wj���r�kH�O�5�U&4J�3����=�i"�=�}��� �AoH \,��DV�/�ĘWp��0I�kvBe�籂(��c]���W�c��"T
�՘�P4��9����Bz@�tT�a(�^n��X�d j�iMU�����E�6�- e�"ۘ�M�K02V�~hJQ�KT�0�9)�nc��9�6 <X��d4���t�'	'6^5�j3�0u��$]P�A���B]�2<� ³p����&������]��!�,�J��� SS|G#��RM]�]W�t����¯@L�=�)Vi� �%>{��l`��C�����!Hߟ7���7G�7�tw��z�먟� YL\�g����C�����3:�--.�:��'^�k�oݺ����djz��ͅ�L3��a*�Cm*����M?�*�ɏ�l!$S,�ef�Q[*^��z�-�ÇW`�T��j2�����SR��Ɖ��>^MF�	y��{���L��P�'�a@+�6W��A]�4h�y@Oj��Q�N�:u*[�;�~�V�Tf����!fm3�����c8~g�8Gmd5��"AM_�R
}�t��Ғ���(�裏�{�L�X�ѣ;r���f�)Zbj��X��5;�<�LϚ�J��X"q`��wk~ii��-�5�S�lfv'Ա.%�b���t��~!�YL&�vn�����l�+��6=�3㘹�ױ�,1ӧ�m�=�e�� ��]V�;��E3��E��=��s�H��$�L��,h�i��^��v��ٝLn/���4�1d&��ʳ��_R6�@��c%�vCG0���eZ� 
O0�>	5c�\��L�vm�!�npbPs���E؞��s�QV�Ng;s�\���(�k@�yñN�<m�jK��N����g��!����}	��3���.�t3�{�
���<:U�;m��iǢ�tU}1�iJͲ���S�C�^B-x�R��~�A�J��k:�
�����+.ޱ�{��P�	��,&�."��C 3l�b$R�Q���U�J�;Iy�щR��:�� ����$ɪ#=��Q~	���c�vAv4s)߆��U�e��4�ae[Cy=6��Z�jl�����ܹ{7g&ggf��7��]�w�>��_�E��;�$	�d!�|@乳gy=�������F�W�����c+�4��)����x�*A-�� &	�5��1�IC;j@ϙ�'V�� �t"��YD�璂�7�}C�tǿ#�oP*�k˨g�Mɕ��ꜹ��&|�i��	�f?�U�,���0	ɜ<y�.�A�L�6G�� �^	�'�r����(|�!�;[`�3ާ�:N4�]�v ��q�ܹ+ 񑑑�w���>��#����稓��:�����_�J��h2i�C��R��� ؖ�������P���Q�x�9��<C6���mT�]V��Z��.��Kb6az�(�2�ȡ�x>O�b���ĭ�ڵd�z��#�N���X�r#�*�<z�(�j�< �v:���~��~��(�Ǧ��,�k�m�P0��@}O��/����1_m+4UQ�x,��������Y�=	Ǐ��vZ�0��tMۡ�fnovz�g��<iR�b�MmԆ�F��S�R��=� �NB~qiniʖ���jR�t�o ��1��������y(�
<^j�,tHH@ �E5�a�ִe�K �.���c3����wQG�%�7��/0�<U�I�D_@k h�
 �@��U�ζ������U���L�`V��H����w��[�"�np�h;H�`�%9M�c�jŦwhq��]f�	��;r}� �%���|E�c���|�+y�@���#G��	P?~�9��s������m۸}&_� %���2����z�dȬG��o[�6���m�&t8����H%��R��:�.���ޢ�o	�� !P�7�����S�N~
ܳ'N�X��o(�FĽ��o������2ls��w�_Ԉ���(�NB[O�j�- �\����}��Ed,Q�:��Ld/���]�ۿ�ۙ|����r�Ȝ�_�<VTӔ�̦�37�K�W�ī�V��b[]S��sT��}�;��'�{�����4+˱���P�G�f�����%�g
��$@�9�V��M����q���K�����W�,f�5���?�����|هz���}�<��Z6˴jTM�Vੌ�:�3%�T�����W`_�h��N&��D2��I�R9��b/�-�R)��vT˵����^e�cx#'K��,\�`���aP�8t�%�'� ���c]v(�r�|v��V,:�/A�>Uaj�d�3@}�Fu�����##itՁ�����
�=����*��K[��V�T��0����R��'��30L�P��氌�j�+a������x�F&3&�p��\�t�&Q�N8��z�Q�BדUE�ZmA%@��YN9��C��Ȼ�})���4�LA�}�]��{��l0=�J��ì���{�fr��m7��ȋ��xTRP9y�2� F�?�`� � 9�98�U������\�|��0}WWoh��	����}�a����j{qy]�9�l��������� m�U�&
�m#c���qNo��ް6$TJyt&��ʀ6d�̌����}�ʔ��ɎG�_�Oؘ��^L�30V,��e8p��y�i������4�ȍ,e��]��^�qm
�z s�����V4m�	j��too�^*�FaKB��	�w�����1�/���^z���������[z\+�y}�y����r���J��_�f���g9#�m�vJbN�8���U]����N���V6�%t�9�f�o��U]�vj˃��u���w���T����,u�T�
��Π���m��:}�8kN~�G=����d�0��_�j���y��N֘$QM�̙s��g�͈to?p`��s'Q��L%/'R)����x|˖�_�җx'��O|b�����:E)BJ*%L��)��ު (���l,�B���� +e��z�ݳg��K���̘}}}3�7�@Vql�{��5gT]?�ڜ(��w�=�����ej;�$`��������{�(T�Ub� fF���"��a�uZ1,� ��C�����r4�9V�BT�@#J&�:\���,Oh A�a<��$fa01�
42w�Ȑ��j��q�D��D0�%��i=S�mFL%��`z	�i�$'�����
����?q��[�A����G>�J���:� K122��O�i8��SOq�M\r�����:���>P��v�``z�D��>�
�7"I}�`�y��:*�Wi)l�zb�p�U� �G��3a�}D^� �ƚ�5Q�a��m��@2j�Q�o4�<O���X��
ԄM�-&`�9](:�������������5\	hƔ<���.�7��~� ��1h�{*��V[� .g��A����uǎ���˻�����S,w��}
7S1��{l�{�)���r�8�����C��͇H.�L��c׬{R����}�lCD�jozF����|�[_�4�I����G����H��ҷ���=e�&���ՙ>���P�2�ȭ펙�w�I�*��Q���������$�x���O8�>��z�\�
�(�����_�5�\6V�+1�>��S����w�q��0h,��0����,|�_� �����_���*��1Te���T�KϜz&�#�M����趝����|>�/�WV� ��H8.�ʖ�dC����p9��O*��?^=��wOv_�\u��{��y�fY�?����y������"Z[Ѻ5x&�x`����
���+�>�]�Y�YvɎޞ�TL�����P����m��{kfXv�B5�V���0e�ە�"#[F���0g�d;4!�G{$�]��
&������~���p��e�}܃kb����aF�F���n�w�6S+��m.H"��: 1$2�"��v��єCx�{��9TCp�K��7�ƕ�6��;���|��6��帛�(�Y��><�������*tO1L��I<�)�8�!'�lf~�L��lLKWٗ���)�L|~��ڵ6����9��U���-iHr�帣8���-Tc���/�IG^N�x+�6�[f���s��ã w-��c5SfP���ׇ��~�W`���q��* S&��_��_*<����~����ٮ��U�'��IU�Uˀ9�i�2����E��67F��E����ӽ��z�n���Ώ�9�sƷ�%�S����"��%㽚��e[�W�F�N3�t(ޣ3��CQk ��$��K�;��w�j��p�b������B�a��u~�qj �( �ȩ9�B���?��,$�bY�W��o�_��W���_�5��W�����>y�$�9Q~��ǳ��B�qUӘ��R�XN.8><��ߟVi�djC!����&d���g`v�q,�^x��?;��7�_����##Z
j�����\�2~�[�Zy�{�{z�y.&ɭ�d*�B�����-�*n$|0�N�ƎXt�a�$�� ��3��Z��ɍ��8���� !�Nޚ9�4� �PϹ�RQ랻T�"���*r�@�z�@QZ8����'�sEd���sBy�t����.���-�J�����j:Y},�ㅫB�垽{��%�Q��r����{�M&�C�rd:����9{�Y\X����7&O�;pۅ�tc�L�\�����0}��:��VU8�l^�Ίv����<����kPD�F�����Kb
�h��4�����V������ܜ��c;�߲�îe��k�M�{j^���-������exӓ0�LPǙ*)�|�+_x��u�t^G6,X�qL��A1y�KP�����P��/�@��#�0v��YXX����=��~���i�W��2q���hK�����~��R!��
���r��b�ƽ�BP��X�=����_}�9��t&]9t����#S�C���~u$ٝ4W�ء5oY�H�	�h�@��J��_dv��bɥD�^����z�LW����S'��S��������8�l��8�~3GɆ��70%�̵L�ή���Ǐ�6��eb����[v(�l�~��N�l]ƣG��.�nK���q��o~�	���x]*�������y ���`A��,���5V~���i	0�}q6(a*B
m��S5_�'h�& &��X<�� �t�(�%b��5�.y�W5��b�����$ggg��W8~\��S/:zz#x�p����wNA����#���U���n%���6�B���Gʙg:��G�������ˆ����9�iz!K�Ⱥ�L^`�V{��-�^w�L��]���65��޼�,�ږy�}����Wþ��|�6��n��N́	����D��!�����9����C#���3MժjL]�h�DH&��t��|Q٩��"n�2��2K<D�
;��Y�pJ��K��,<������y���/��/9�~�~��>���m�W����g�Lm����}E���������� B{a;I�᷊1�����]l���2��ù���ͧ��[�rl��z��Z����Fz��(��L�����2�=J�nJ#Y�{�o↻ť��{�O�W���نm;+̪,�hqı��
x�.0j���g��\�����l��wu��!�8��:ރ3�>uMڷ�	�f̎�l�WU>s�6==�fk���'�� t�e��p{t<�KW5.T��=d�8>�3j�&�R�a#�����޸�)�,�|�3M�kl���FB�&�1j`DR�7�zPoY�iz]� Xƿ�-K �P� 
�h���e�Zd�[�9�x"�#b�8ٹs'��א׼������F����_,���!.���Lt���[ȡ�o&�zի8�DP��ɓ��Yt�M���y�(��FK��T6:\߻�HS��ـ�Z^!Z�&���pb:�V�J/3øan8����<Z&��{w\ь�J\t �8~Z��_+r	Go�b4��jEx��x,~��D\�WX,f"�iÃ�I�Z�|2�� &\�U2Iz�F�Rebb��X�����ߕz��)�f}��_���G?��P����*�:����B���!B�����o{c�%\���������|�c��i-ݸi8o����F���P(�h��D̩�4�_�?�=r�m�Gn�ӂ���s�@�@���J�A �����$Ѡ��hYr����x/o'j��T�.S����.x���)�}�w�! 1)�u��;���#�����W�Zu�Ζ��4Np)���T��G��iNM�ȟ���A�5st�j
*�*)K�ه/�'��X�ӽv# ��6��Z
�iz����0&��Kv�,��N�.��q�J�D��88|���*>��>&XCx{�������r��;8c>77G�HuVV��w�a���3	 S�.�O�Ls���z_C��t�Mh��'6醗�8�%%W�R1�4q� f?��4q�n�ڡ�Z/�Km�`y��jT'kF�ԕgR���D"�&G2�P�{n߮�,��h
����+�*�_G�?���ٗ����|��ar��۷W�sP=�w�I�6.�
uJ{��ȃ>x�S��T���5�7_�^����vժ:����z6�W���f0+_r4?�'�8��):֛�G7�ɔE�X�Y�քe�->�8��Y�0�\�G�!�&;NTur��l� �H7�L�;�cP�)�	�v}c#e� �k$�x�)cT`�ĕ��0`�p;���/���h�h����G�o�7c\MY.�I"�>]�${D9�g; ����y�ؚJ�S�}i��f�9x�&T� B�.������3��Y��Ȳ��U-�aG���D�Њq]�$��4& 1n[��QElL�� R�z�v��j���z����1���̥�\�qի���~Pó�R6����9�����gϞ->|�֛�U�������)��J�/>�0�_!J
e�*�5a��;�u�8�zE��i�d`�n��38��مT*a$2=��g@�u�������iS�K/�������$�8������#č��[7��y�̙3꧅L���K�M�n���M6���7�|L�Ǩ�)o����Z�����y�5���
ef���e%��2r_�Y~�1gjD��ԁ�Dg�H
 f�x��+-�(XTSYB3tjC���$�����W�}�l�s� �k$��h0�R�m+L��NA�En8ძJ�"rq��q���N@l!�LW-zeWY��g-:����,�N�բ9�'��W��c��o$�g�X�[|O�@�iQ�~�m�qvu ˅���W��ô��9���z$� �4�(��@�`���͜ە]ʮ��+C�*��pM��Qޤ�bA�O��}Y���N?�CН<yrÙ��v�#�?~�<v���C=�f!&\���Vy4�)
=�g���d2I���o|����~l'm1��������bU��@+{̲�ǫ�>R�1;�#J2�%����o|��yd�*0��˳�vO8���)-yx̡J��L�ًĶ�ĲkJ�9��+���2'%x��01r��2�˚����'^�'��n����ʴ�=�����y����נ��ܑR�Ou ��H� �!,���؃RW�y�F���j)�О-S����NV׻�q=bè�J�B��*W����<�V��yf���� P�=�5���s�����~ݟiv���َ79�gk��^״�q`����g������޽�lۊ��s|+
��ǽDed*	� W�B'�'N����o�F��~M��rIu�,�cm.��,:�e[Ds��^}�8-f�GQrP�k�(��$�b�6]���Ϻ��g�q��GV��ل�hĺ#�Z��q ��=���g���ݭ���ϭ01�}z�߄6���.]���V��|p��ѣmu�y8����;f؎F�1à��zumG�T�ees���'��
����
�I�\u�G��e�	4�aZt�c���EX��CQ�v�����p2KhM�񙽑{��t-l�9v@( Q;�L��+��?P��XU�k$��h��Ts�)y�����c7
��F�%�ό��^��2���V9��cI���&u�t������ b��U���
1�:z���XWz���r�X����u/d~od@���8�ĥk1p���\���+MQ�w��K{|^�)����H� 0m�A�P�A�_���9.�1Iq�Z������YX$Q�8��8R���q�HG�"w�y�������XA�G:������ZM�����ѝ�f���py�������	���_f�������	��SZ�VߢY��x���.V�OJ���D�e��N�7ǲ�\&�������s=�7%��-TI�K�d��w��L�R[g�q��T�Z�T�a���u�CA_B�)R �h5��E��%V#$���1��Ls�%H 'u4�S�v:�0����g�ǳ�`:��5�����/��o%M���fS[�FWR)?���y?&Ww��8 ���L�$�cE����ykP��O���s����3���rc-�b+��u7�A�QU����==$ �>PjR�tn3���Nc���:�ո���ۯC����Z`5F6�*�l0qs=�U�Td�J�\*r�dzz��7::��	���0l��O4�y��7�LX�i�}��-o)�*L���ّ��U���/:hw�s�N�`��.]�~��m�������3I��V�����'����)��ۤ+�?ti��r����&��n۰Y�Q��-�&�"���d���Ѽ��'���dD�L|��:��Rvud�&FvC��ԩ�4�r/��*s捌 �iYW*+����ڀQ+�
�kw2NsrU���� �k-|I.��B��*�eX�W8������"�v��i�e��^��}+d�'[�l��tuw����v�r����ο��>D�X�&&#�<Y^^�l&.�ೝ:��<O<uo��/J�~����3\V?�� p^�Ѝ�����#}�9�Q�(z�����#A�o���΄Q�Ѯ�"�P��0=::j�Ǚ�#���L�>8 @��H$`��G`l����WVVv �<u|
 ���-���+�����������T�;A�TR�)�=1��K��>�Pd�wijo�bmI�ُ?x���?��J�k,�O!x�r��b�@/ѻ�bqmqʇl3�C�r	𛲊=.S����r�ڎ���PE�Fhb@���)w�1���GE���f����!���D�K`�Ѐ%U�P'�B$�.�������f6�Q.�r���܃�4LX���R q�3��d
���%���dK6��lʶ��O�4�؇�[�V�NLP�$�[|��ȭ۶�C�a\c��G'�s�A�>1��bb<L���E��K/�c�>����R��6�X*'T��b�~���Vc0�XL�iݹ C	�w�, ̋����)��/�4�EF��P���%%JZa�C�s̱'`�^:~��շ�HGڐ�G�:2��H��s���П��4��X,n x3��L������_������]����gT�8F,f�]�w�jꨕ/�Q-��,Ӷ�Y������?Mȕg2��r��=,Aߐa�?��X�E��K��5-E-���_�T��=0��C�zUb{�G釾,��hnTa,��x���f�N>ItHq,��^�R�k��������!�&]�pq0�(��!�ဏ ������E�3�YS_�P^��G�J��f(��=����Z��j��,i�L�3ȺE_�| ��g���BDP`�(��;�h�U�� w�%&1&^759IΟ?і��E��67<�
�����NkQ�`:�ی�Ur-�s�����8=PH��4 �B��-�6'z13vz�;+�����k��ɓ';6����s�Y��G?zrttt�,���FFF����}0Qe�.]B��VVV�3���3�����j+z�U����c_%��f:��n������Ϝ���]3�������ͧ^|w���L��=4��M�$�
 �M�VT�O2�xIcΔ��n���f�1\e�ޚ���L��H�(���
n0i�X�?����5�dΒ�԰��΅ӆ�v�Tʨ�5nZ&g��"�u�� �T���pS4�Ky���,�|�JJ/ҬZ�6X�� ��0#ڊ�\O\���*2�h�P���D�B._��ˀ-.s�pe�NBp=�6�뮻�/�}7ٶm�Wh�`-Ó�0���Jxb��MN�vG��+�p�����k ���UP�H��mrʖ`�j9d-j:�-,K9(-�{_ܻc���������#���s�~@d-�ۃ���4M3	�7-..2��Z0!���?��8Y��6�����?��Z4�J2n����Ӵ�J&�G���*����i%��C���~"M�����G���l��{z��J���Y5����`�v��I�$G�fb�}���m�0������0�2�(��*��������$8�FS�_ĭ�cr��J%��TZ��>l�����7�u��U�Wi;*}��t�|R��Q]~O��`����;�\��e��,�p�|+���4st�*k�`��]Ў��cP~�6w/h4c��	�;�X������g��x��Lybj+^n~�yC"�5�'��0%v��0�[e��+�mT������$d��ե�;[w#@'	��֑#G*�<�����v�#�H���6���G .�r���r�7B��b�\��kە���F;E��x��+�O�x�3��-4[7~����F6��P(*v:��I0[�v����\���a����gd��m<�؃v.=_�w�z3�w;������$�� �k&�#��,b0mt�UwQ��&v��A�����7��h�T/�l1,�m��k���F��s�k�7�I��v��j�n��7K���
�nX�w��*��ޤC���48�b��21���O��_"��ggg9h���4��M�K��|�`� �x���� �ޛ����S�HG:r��W�򕅯}�k�}�;߱0�Y*�z[>��W�ս�t�<==�hY�<L�2�v��u��s��?>ce��k6��]��2T��Z�ƬLήQ�؎�M�3�v|���y�*J�������0���\c,O83#�Q�7-�L;������|aھ�h�63,���p�L������1���M��� Q,V�	��5��@�
���U�V��ÿ���N��>���o#�ڂU�L�j��M�� �1~ %�42j5R*�:������U4��H���&>�-��ͮ�5�;ґ�W������?��?z�R���Q \��\.o�t��Nhϻ��ƶ��=����?����w���2��=�l�V�tJTK��y@Uw�VV��sy�,gG!�Nm{���P͙̍H`^#�+�H��:$D��D��E��}���ab y\�j;l�@+���Ր���,���l��Vc��\K����6���0&���9�2�M��wD�	'j�$�IJ,L�Mi�rl��k�Cޑ�t��|�3����׾��7���h�{����e2��Z�6���۷�������;���<�_�I���f/~�cO�̄U�٬̜�z	���>V�2s9è���&��S�[��K��p���P����H�܁�x=�\��8ĸI�9����i�nr"A�o^)��A̈"��� X0,Q n@�|�[zN�Q��Q
����z�W�2�Q ���Q�g���g���<j��Oݪë��}d���u�������T�6$���o5�יv�����$�T�
���P�h�v���HG�S��?8���x2������ӧ+++{fggo_�~���rd���/|!�L�iW4zS��گ���˻�|VqVrTQ���Xᡇ�ʲ�WB:}\G��Ȁr�02����|ۅ$���0���{�̭���e����M>h����;��'#��yG:ґւ�����޽{_��b��
���l�
 Ө�j4����Їj_��WQ���A������+vE�"&%�;��q�:�c,���=�������w�ü���NwM=g	��r��H[;���K�ˊH̤S�w��[ 3�w����Ii¾E~h$�9E����v hCLM��B�=V���v���	[����R�si��kR�Vi���J�~Iv�jt2��U+���%M� M޹���[8,�Rίn�*xh7|�2�΂{�q�q��7�
 ���};ґ�U����[�lyt~~>�L&���ӳ�T*횝��.�1�w�\.�v��=y���u�|�Or��X�1U��X���^]�Q�[�U�f��N3E�mE��?��.�����_x4s�c�n�sޕ�Nב�#>n�V+��aB=�g]d���v�>��$A�e\Efey�d�Y�r��_�IJ+[0�)�e��������+<]y;ƎD�r,�@"p:�X�N����Ahb��L�η�HG�w��?��������s�=�K��a�E�߷f2�]�7d,˺���5y�-�̯`�������G�	MRی�5E�ޢ;��$s�م�c�-�6%#j2uQ�763�ո�<��4}�k׳�9J`^CA%�	�.o��J��vd�k"c ��M�ؒ����k�gD�-����5
��>99I�;FΜ9��&_{]���~s�0q�ěo����U�"�==��H#�S�ҊElum���m#���7��y�D�;'��nk�'��q0Y����7����7A��+^�8��HGڐ���}�O~�����D�P`���o5Ms~oUUu,�Hl�s i~#����<��_<�3��t��wk����n3�M�����t���L*T;S��9�z��9����� ̎\	�H�o藯���Fk8��L��WV��ٳ|Ml��e����p(����.,,�< �!H�K �?p�AeۑT�z]��HG��g?�م?��?}vii� �Sw�@@s��}===���������H?����z�C?����G�J?���O�rB����;��� ���m�����Ƙ7{������ʽ��������P4�[��J�ߦ�L;l$m��.���2���r/^���H�22Nd�š=��L��.i�DC�Lx.7ɫ�-$H\���X<N�v�$�|�+��ݻ	�t�e�Q-0f#z'>w�8^�}KxC_!	��lG���^v�
{�7�J�����S��6�®��{����Ħ��HE�롰��Q���J4��"!�IG:ґ�]���o���߿888����+�ݙLf>��@�^ƾ���WX��}�{��g�/�p�?��۲�����Q�܅���m�+�!�*���9ڶ�,��);vl��yg�\�����:�jdy�������p���Ȝx���"[O$���W{�v��\�m�i��Kg×�y��eG:ґ�td}��OT^��םQ凅B!�L&�Wy�\�p�Z �N,+�����<��%�qG��O����?]�j:I%t�i��Rq��}�j�dT��1�iU9?Ir�~�a�W�#��@f`^�k"��H�4
��G1s�k���餵�ii#Rk�������G�KN>�o39k�4�-�����99�6�/�s�y����)*�Oنo56A%�\���^ &�<,����y!�׼�:�|<��X�0������i�{�xw4���4�7�x�"m#s����N�U�c�3�����?�%A��@z7PDԣt�#�����7��'N�?�J��T<��8��v�T�蜇�'}���)o�u�������9�m�8K�Y��rӳS��MB*�21gfm�Z��圲��/���Ǯ+uy`^"�k-m��CC.�E�ޫ[϶��wns�UU�MT��$�{{+��w+I��^��<�����!���!�p�,��̤�dzz����so��nBћ\�u�r�냯L����r�-����7Q��\�4φ�`��T�Nq�c���$�HGna�z׻��'rܲ���8�i��o�9������ݩT��w�1�Q�����w�?�S�st���Y%[�f���^z� �[�8PJ�PV��İ8������j�h���sv������\��t �u#�x47$�F��ЀG[���t�CQ�w�=���'s�P�sX��q/�&�7��QX�s;��d��`����A!�!B;�`vu�A�ںmw����p�a.�^;�o� ˇ��/����244ĝ��<�Kf;ot�w��,BJ��qiەԏ7�����8Ϣ��HLQ��d�58�5�FZ�$|�=�(ev�@��HG�G��?��������B!��G�x���$�Uegww��X,6I�djr!G?�]��'b5VdC����F6[�U���S��R�|P�V������1���J�p����n���jE�_Hl�O�{�Yw��H`^��6iU2�5�[\�<T�WJ��!T�����P��C�|��}��ɛ���%����z�_�ŏ�)�;�8y�PG6\_31�%2�h/x_�U���!�ܿ?_'=�O��z����s�"++i���@����]�v�-���)�d�u�|#��	�l.Kʕ�4����NT,���/�5$��	_#�K���Ν�n=c��Σ�s���׵�p�
ԍ4�,7/i�fj�v���t��O��������o>W.��`R�㡯�^��B;���r�w�}w���Gu��A����n���Q;�w͔��/S�jE+���7�j[����j>�e�J�B1���j�֛lk�>S��;�y��9Fȩ;	1�U�����~��$�FnBZ��u9�\A��g�" 4-�vM\���۸��^`�j�J�X�>s�X�M�����)���Jl��;���TW���i255Efgg9 U<�P�rp2� ��|��ťE�˼U|�E�Y:4��͒Ix�b�t�c57{t]�"��d�Q�*o�M��U���I�E4*Ơ�P��d3�v.�p�=	�Β����w�#ٸ����e˖˩T�"��= 0{ `S 0'��[�@�Ĝ����9J�Y���~HV��J͠�\�-I��R���������L�3��7EJ���#��G��I����:Mһ�qHQ�(M
8�{\{\���ii�j���)�� -���\Iܺ饭zI,���-���c�ܝ���D�e��-Z�?g�����P�����'�ig:#���Ę��oU��DǗ��dO>1K�����A�(�ۉ��W!��~�W�&ͷ3�:_�li+8]�Xi>,�Pڄ���l4`�X�b�:_;�¬����t�͗+�ܼ\n��r�$-߿R���&d-�< dm��8��3 7`iN�ggI2�&.��
�i�+�T�G��8�RI	GHZ���j6{�#����bQ̄ۋ �lp�lNW����,�ޟ�����밸Q'��:7^�1yWq[��_ҝN'I,3��k�@�j�Jߗ��7n�N��fYV�0Ud�g���ii�������C�T��qNI����;�&D�C&���n�[#��p$��ȡC������﷦��fx����� ����l��㋁��_:<oW)I��}3�ȁ�&��%J,A��a"�$n��L,J�m��x��r��[�ȿ�Z����3��*���*�d���� sԵ��7��{��_X�O���%ˮX<��[���jQ�a
�����f~)=��P
���T������b)�%_�C+�G
�7�h�D\7��Jn�2��G�ٿ�ҟm��i�K�:ѻ5u(3jv�]6�Gt?XW0KN��y�����4,��SB&�R�B��[������|k�ȏL�e�l�ùg�r��	�����,<����'.]�����G�F�ԩS����y=�n��[����%��1v���w�\���rKſH6=��?��>+�և4w�c��&û�?aK�.�u|�hC#$�v��-��55�G��½vZ�[B���t�/�q���Vo/'o�E�~N<�o��9S�'
�6"~����B3]�>�:ڶ�0ͪ�޺%ֿY.G2Kn�ei�JϹb\c%�̲G��-��Y��qIV2J~*gqg�"�eF W]�8�f�ۈ�1�d�ȒlJ/̀#n�tM]���A��d2Q/!�9�?�!&�^�G���VI��Q��A?���v�sÌܙ�I�_NK�8����34b�ɬX�1]�.��粺d�B�m�M+�r�$Sb��� ���{%�Pl����^�+9�PR����ϟ�4�3޷�ږ��8'y���)��g�J~����2�2aSp�ix�	�LdsVA��;�#~��ѹ������"+���d["��P<��a�������m��d6�˓�O?����5灃>��w@1���{��o����y"/��zF��v��(-�嚕]�).˗j"���Bz���4��ѤJ�m{���O�<�t�uD��F8����؎�2�����xqYNX�1:	/:@97c�&qC��^�[>HP���BYQ�Q�q�La��|� ð� ����"R*���+u��\ڬVS4�В:q�/fQ���B!�D�����Ab���_5[7��_�й�2�,��xol���fw���̕��߁�9K"r�J1�{���r�Ukb�N�xa:|�Sp�Yx��J')c��#��#U�A��#�F���?2y>�톿s�\.�����
kv��9���ËW3��Ft>�xd�������7��=��xJ���H�]�DO���7��6����٥d+K���j�6$�a��1%�p�S��.�nԸvg���ɓ���h�z<���89�?���B�ש��(�ۄ�KH<���M��)N�#q�M�W�ZՏl���^g�-�b�"�)Z��������1�_"T�1���0h���e/U(�
'CLI۸xTL\nF�������3��7�L�5�X��DF�50#�%\��)!�U�DZ"�'^��f��a%�*��ru3
e�B�{�Y6���/�2�l�|�
�K��߶�2fnK*z�f�*��X,!X���~̃ ;��`ss�oA.�p��n��b��[TU����������dD�lJi�#H-�s��#�I�"�6j0�{<����(+�����S�����|].�v�l���7r�vk2]�SvF�<����LÔ�����z@���7�����Z�?yV)\�4�g=��J
?ka���MȲ�%���МD��fs��ƅT�M�j��~j�ǖ��E_�A�0���K���1	�Q��R��XF̈��\"��żY�+e�:�k�^G�+Ǳ��:u��Ϡ�Y�?�����\'��go�r��bI�?^D,+2�A����ٳ�cǆ�].WWCCCW0�K&�Mp/�}��i>�kҊA�ߙ;��!���:|�Q��uX���RHJē9��'j|���]�t�Ԍ�S�CU5�K2�i5K���M��I"b�R&�Q���⶚�ˑ|߮�JH�Xe��O��:g�h�C��&�~Հ�Y�+*)JT�(i��8D��)�������b��5m˛��-a~5�S^8C~�g��ԐR5"Lc���� !+�.��?�9s��e�\��ѣP�r���5u,<^�6G��IȪ��Nݎ�X�+���/hk��O�ڳ���>%�!��\�p!�v��===6��3�N$�JyE�w:�m��,��E!(��V��C$w��G���b@a���#e$Sc�f�����Qo�g���=� �Ĵ���k9�2"岠�R�t�b���0�%3'785�3B��8���>����%��d1�
�6a���7`ގqY�Z��q���0WņwT"BIB1�V�:l���e�R��M��lQ *-��K���&�(��HٙjU�j�We���Ax��W���+�����d{]]]��iUU�p�������@  �O�S�����q�����6ջj�.Q�%ɒ�9Jd�
Y���i.[C�T/Y,����kM�3�LײT3/M�(�pq�*�Uz���b
=0LY�͢`n���ZKooНˍ)�w�l�2Ƽ�`� ��Z�,R@7~�t�$mK>#��c9ֹ��W���L�|ը��v�H#� ����#G�,���aY�;�^���l�5J�T���t���r� |���������g��%��?��,-��x6��v^[kS\N7a��˖=�U9�$|���4g4��\�d3ϋhQK���I��}��cj�F��>�Bz���N����O3f�_�I��ϷX��/�haM�������2��\>z�r �Y�/���A���ק�<yr�f��q׮]� ��aA4k��h�������l�ԧ>5q��������C��щw�������*K4�L3��wF��y9�q�c�܅ҌLrin�YN4�"��3��,�� ��13�3
�6�r��Y�]04m����d����-�d��q�墺2s�ߘ-:i!��HB3��'�Ѹ,{5�r� ���?~<����_�pA
��֚��F�:UU}�����+���:u*�裏����t��FI1/g,p��K6�%x.;E8s�*�:/�5n��[�n�IXR���Rݳj���I�Y�嘈*q��'��*|s���wI�6�s���q��+��ܬ����pJ}t���Ց���C�ڷ�8���$Z����E�<�!��Y���n~�*7�AA���zH=w���8 IR&
���Yo2�잛�;�p8�KKK����ӏ=�X�TM}�%����3��CY����?NHoo�@aY da~%��M��P��m;"G^WWW��M�p�Yj�9֟��J���Z�ܰ�&�zE��k
s�X�S:*���n�������Y� � ;�_���9��p�\�ew$q�`v�����T�n7�d'O��8~�xU���3}���mh�*���R��������9���k,Lmm6q�F)�g�Y/Q��
�����_vuP���*[)�<�㪃J��ʊ�%M����?��?�l����!�^"� ;���>�;���H(�o���{��a���go:�& ��@ ����H���v�D(�U�aI�0�L'�`��5����1sn/���$	�9�:�C��53;;{�r�!� �6|���cǎ�FU�Z����v��R�Z���D"�(�u�\G���`"ל���Tl~~F�(Ä�NNx#919w��O\�Z�S��5]�A=婈V�Yݟres9�)J�\bU0�烕�9�K"�L�U�	�5�Yx.�r� ��d�^�{��A"G:;;/H�T733ә�dj[`GCCC�޽{'�H��CA��Ξ=�wuu�]��l�2��P�B$�]l&�����s��9�E"y:���%BAv6tzz:{�m�M�\�����%�Z�����p7���Pf�ĉ��X���o�M-��YELMMi�H\�9���,�̥EJ󭯒�5�ƲQޥ���r���'��6KB�����$�?�Qa�<�l�0>De�n�/�KAdg����SG��M�v���yH����EH������pJ�����cd���Y]pUU��c3�:@�jĀ�V
)VJ,��V�5�lb��*�N���A˂�U��D�1�� ����AAJп��oG�|�ɡ���߉�}��t/�ef���l��t���:�S>��={VdV�1A�����&/v_�6�d ���&ç�x�mm�b�JR�^��r��+/[�>u�3�O�6bZX3�Azc��s�I����oi�M�� � U���:u������r9e~~��l�{��+�x<���%a�X�h���d���Ye�!g�Ý�áP�"!5@ר�kDL��w��e���x�)0���K��@��)�&�'��v\�AٌG}4�9�:~���v��եi�͆a�d:gffn���,�s�ݓ �(Ov
(�U��s������E��,&��	XZ��l�pDθl�-�UIi�$?�:�Q���'���{��Ο}KP0A��R���>���="�.�򌍍u����������S�U��؋0�!�`V)B2a��s�mĪ�*�F@"r3�DN�Ƭ��]�`�L%��dX���%NG5��Q[�f�BA�"SSS�[o�����j���^���133c	����SUu6��ľ��/��^z)Jv (�Ս1��{��~��g�����>��K�oG%.pE�@nB�N��a���f	\�w1LΠ\"� hX��'?��IY��wvv�Z�=p߬��b-�\n���b������#�\:}�t���`V?��w�]looO�
�V)'�&4�2�ױ���y� � ��g�y&��O477{t]�G�ѻZ[[;@.oJ�R<�NˉD�]�t��z뭣�ϟ��#�(�7�p�~�)� � �:�zj��;;55�u:��������0���J�� w�\2,��d�:u*!�p�LAA�����;����S�٬�J�>�iZ�o������ւs���^�cn�H&
&� � �u�?�A�g?��o��_�h������r�z�=�d���x�<��3����7Rp�~#E3Q0AA�3_�җB���7��� {<�s�� ���T�{nn��B!�D��aM�?��#��O�>}C̊��� � �|���]���p�6�M�7�b���hTLmQ�!��N�����޽{��_��򗿜"U�ѣGeLAA�m��_�|��_}'(v�]��_�elwg2����.��Y��1%IҐ��?��O�?��SK�
av�^��� � �����?��G?:��o2��j�<�r�Zc��M�H�yzz:�9����o�X,v��G~��O�y���� ��/�N�>-�N_�Y�(���f���~�����YS`���NLAA�m�+_�J������i���Nkjj�;��_���D�=��Ի�nWMMO�R�+��RBM��Z.��|���C�"}}}���goo�D��)�yZ�>���S��ޥ(���AA�
x�駃'N�8���$��c�u���H$r3]}(��%X\����'\[[����$���� w�?�|���i/��"���i�L��(�x�����'p>���`n�u���b$��we�Z�s�=gi��r8� �.!�$�HX��&I�z@xw�`"� �T	}}}�O�� n� u����;�N�}�X���tڞ�d��|:��M�/	۪,�1UU�@F��A �333����x<�F0E��K�.�p8ln���Bl6hkk����9�/���p1	ʹ�x,���ݰ��X*�<P�륔���&LAA�*B�ɄU�ĉ�C�5���q��ͭV��A�v���<77w��r*�� �3�$��2�(JR�4џ���v
�	c+�3ŬA"b)rp
\.��C�kjj���p1����@ E���P�JI��l�u\�d�&����yY��:XŹ@�1M� � H����%A���Ν����d����t:����I�?9#�A�DT�eEu�2�u]}#E4R$h_N�.d�3ES 2)���~1���i�u#ȣ�J���i�p~!��P�#�iN9�9��Ρ��Һ�:AA�J��ǹ��ǿI&�R(��F�5 q�I�t�����`����Ox�)�p��S6�\8g�;��I���~.�2�ce��[��h:"�?!p�f��kF<᱐�����B�����&+����|(�� � ���?����߀���8;;;���6'��G`[�����,M�P���I1 G*,��)'�H
ɴX,	d�H�/���m��r��nπ@�A@����������f@vE3;6�#� �T;�H�� ,�8:44d=s�L`aa!!Fo�$ZA����X��9ʋ�+�#�Q�e�)dR�?ae���2<�:I�����'"����"�p���p�EQ�^�w	�r�s���}��{>�������_�(�� � 7B5!�@�ĉA(C }u��ݖ��*�����V��M�z��^X�`���`���& �����<x�8t营���Q��FME���D?�����W���;99)�Ù��¾��>�9���(�� � 7(}}}��8�"��\���/�_���] �s�9��"�����i�̲b-"�b` "�.����z�R}}=�*a; ���?��P(R������7�\ӿS��� � r�ShB/�,b�x�,��^R1b����L�.}6�٬H�N����-��B��Ns������+�t��wG�~�m!�dppp���`"� ��\�$/������fr�=��s�FFF�k��F�y�s�ltt��P�i1���s��� � ����	�#y��g�e#Ξ=k.)(�� � HEA�DAA*

&� � RQP0AA����� � �TLAA���`"� � AA�((�� � HEA�DAA*

&� � RQP0AA����}-V�jm    IEND�B`�PK
     �8�Z�J��T  �T  /   images/91777b75-38f2-4118-94bc-a70a6868aa47.jpg���� JFIF  ` `  �� C 


�� C		��  ��" ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? ��	��2Z|�)���U�E񿊢72�1%�l���y��Qd=���(���=�`�����|`��|����6��K���&)�O�X{0�{+|Cn��ܘ�(��i�ڥ�ŭ��Z�F�M�$Fee<A ��5�c�f~ΰ�̟�-߆�wF𯈭έ���KYG��C�xVV �+����������7���ڣF�4�^v����I��;�=��$W���j��62��#��Nx~tczL��X���&�h��� /�G�I��_ƀΏΏΏ΀ΏΏΏ΀ΏΏΏ΀ΏΏΏ΀ΏΏΓ4 ���� �G?������F}� �h�J��� ��0�k_�_S�D���6�FOM�A�&���S� =h�޺��?�4�a��[���m'�*O�� �L|H?��5����,r��Ύɮ����һ�:� yld#�Yzׁ|g�:=C[���il�P��u�8��'�qT��[?�����4�� �`��{���8��+bE���9���U�Y��N��*2*?�M�_�m�W<�"�eQ&���WI��9�5�� 	���7�G�&�/����/�a� ��~���g��ϡ��Mt_I����~�7�j���㈡7���2J�[���,�9ojA�\�kC�u���k�zm���u֫o�}��b8�kf�J՘'�z@��L���)��)?�$�1��� |7�W�W�Q�^h� ����Y|���i6�f�y4��Pe�9��2� ҫ�|b���xoL�V��)x_P��a��;_E+���ナ�?�$��Y��=އ_�W�M����M'����Կ�i�Q� l��+�+L���Y��X�d�Z�a�Aq�h��Q�U݌�zW�j��R��o���v������m(�v:�����U�='.��=�N�M3�{;�5��&��n?S��޾�� ��izz���:���׼1��aj�F��W\�,����U�@��麽ZZjmnsJ<��f�F�Z�%�r���=�4Sn!{�;�xpf�3/����~��#� g��5_�#ӌ����]y�V+>D� ���\�x��@^:�ſ�J��p���o_y"����'H�7X���{������\��˛sׇ��� [�~;� �J?gko�� 4�xM���_�,Y����Dt	�c���ؒ��0?౟t-^�������6�MR��0I����c�''��/sX��Vܮ��^g�� ��W� ���h�e��� ������U�W��鿲��Q��#��]��|�����c�=�> HU��x ��#����k�?��/o���k?N�i~!�m�#�A`A�Rk�ᵿ�<Q�C���k]�:��յ�~�L�#j�<	⽻����t��GV�5m?N|5ՐC�qr�{[�		3F�eB ���e4�r�i?��gm9MF�\����U�
�^�ᯃ�g�<Yp�D:��L�'���FU$�6�'?�R5ėWW7���z��/慄�k�2N���<��L�H��bӠ�����ǹ�Vh�`H��\.[��0�U�N�� Zg�"� ��G�"� ��^��� ʏʙ������������Z8��}�/��{E�u�<~�u����tk7�0��,i6���k�S����@|q�᷍� �,� �E��x�����?�K?� Y�Xw+�]�?Ώη?� ���_���"��@|q����� �M?� O�C�r˱���FG�n¿���o� ���"��W�9� �m�?��� �Q�!�9%�����#޷?�_������� �K?� I� �?�x�� �� �{HwIv1?:+z?��:��'�_3z�&����.����]?P����s���u<��j�%-�����z�g��GPT��i*�D����@��e�]��W�� ����|� �x���>�M!�Ƌn�jQAG���	�q�0�n�@:��?*���'����0|w��wDԼC�?�b��z]�O.�[vfؠ� �=���(ʜT��7��='�?��V~і�'o��;�� ���]�jv���${Kd����=kĤ� ��|wL~��`㶖��i���x��q���x���ī��.��v2i����U�3n���5��2��6b���é��w����QV��ǚ:}�� C�)�')[�� �������.?g{��B���𵴩X5���-0�l���g ��������O~�?���ă�\��>���N�X��q)e$���I ��������5�����'�o/���P�Bqg�e�č�3Ͻv�'Ï��u��?�(�ᔹ��O�X�n�Nd��C)8��Xzk�J�����K��NJ�����::�d�[���]7��uM?�zχ�����r�O�,s��Y�ҹ��XJT����>��x2�W�<g��x~�t�j��%��$�Zۿf/�?Z���.� ��3���F��c�����o
��7���&�eb,�H�|�#�#��� �^��Qxoƾ��}��@�E���J�𼺥�����Ⱦgr�^E_�V�$�^; ��+�5��&��@�ƫ/�?�x�X}=����N[�p���8����E���Ox�V��ǌ�|��`^���P[5��1�a�����V?����fD��_]�4~Eܒ�O �bY@탑�������c�b�u��r�Y�>b��GpD����4��]��pNM%���:֓�v���+�U���M�)����B����)S�����Z���>k� dYC���_A����K�� �~����5�.��,�v���p�_�ߴ��?��㿏>�'�/�6��-��b[pT��A��<�w��6� ����&����U4��f�-�͝�H����u�_��f8j��[��_�zt���u!��=#ÿ�P�x���Ě���[4p����R~9�̟jV����#������	nۙw�GZ�um��6I?�f�5��n�i��V���Z��=�ҵ��<hR���xeh�(�6�ې9��ҧ�R���v�� Ҽ´�y��u��  �?�W��I�V��>�$���mo��~F�Q�J�J�U��~�O�[�?����;S����g��ٛD����J��H��ۏ,�|��5���Qh�u�̥|�efv?y���<W({9-U� ���;��(�PH=��v:w�/�:���
�isg9���:<��pA�C��5�����s�0����D�t!�M#5	=��_��&��~%C�$2�M����n_ۓ�|��U�:������
a�+�V���x�x&� <�l���	W���ڿ(���~/���'��E=WF��W)�����n�|s��U�'1�k�l'lr���s�s^]|6.zr��%�����
����ޝ�Id��↉�ʺjgO�B�)�bFT�2z����U�/k�:������,�$yo�f%B��tP� p �-�Ӳt��Y�Evb��4�2=���._{vEJ�z}�� �O�|�SmW�as�˝�	�u��Y���!Y�*n#[�2z2���W՗��"�b��ĺ����M����d��Ր�"�	��W˻!1ȯ��o�	|H�<I��Oh��w��(��G�Tb�9�N1ҽ����������3O�Q��h�'�tɡKw��	�����"���v>�|�l%iVT�o����������7�~:񮱧kW:���G$�3lQp�+�`�nq�5��?�a@~תc��^y�2�d���;*����x�^�<���=�<ʵ|=uN�F���� !ьe�(�� �G|+� ��[���G�(�����j�p=?J0=?J�>��� ���?�����Tr��� �έ� |��� ���~uo��� �]N��F��G�1��_�������?�G�,� ��W����?B��W%̟�_�
Kx�Ig�i�}�O�Z�(��b������C�t� ������x��� I� ���X|e� �bq�KǵG�k� ;����=�?�:M7��>����1x�"�y�zW�w߷G��-SR����$we�����8f0I��yΣ�3�V�nu�MJ�k�2�kJQ��Fz����f� �H���7���������� ����� C�� �� �Y��z���J?�|� Cf�� ~R��V�g���#��?Ỿ8� �����O�n�?�?k_�k�� �Y������J?�|� C^�� ~R��V�g��rG����r��o�t�7ǚ��M�$IC���uO��5��o��ί��"˪_���p7d� �J���_x��!�u��[S���[�"��`A'��]�[Ϫ4QC�C(}��"�b��j�}���{�ε�؋�R곶��h.t��c4������b��~�?�x6�Ş(��^�]�3�23Fm ��Q��;x2�Iӭ����[M�q�} h�(�H'#1^I�b�h��?e��g���cR��X����a�iϘ
�rq�׵G0��p�����0�i6~`+����s�d>�����zm�l6�������O<���RE}]�"��x?�p�ů�W�� ��/c�d��k4̑�gV�|6u��$� �y��5����� ��� ��:� �wW�3�~��Z���r�����6�k�M����9x0h��p��1�",��%�-a�j/��9�i������	�� ͭ��)uK���M�kN��	!>V�䓎����|�?Z��MO��t�骕�C�0��{/��:� ���1n�"��� hiS8�O����Y��Ԟ����P�~�w����xCN[��3�z����݈�%Eʷ��Ǧ+�t9<7/�ZO��eu��B<�.jd�ҒU~�N=0M_��E��3��c�,h���{|��ˋ��kZ.Ui��k�J׿U�J7��+�	�K����eS�Gz����m�x�N�uIt}2�Q΢�b�OW9��M#�<���%l�1h�k��%2O�ģ�C�_�����־��-?��1���~��k�#��+�ƺLqE"kc3.Yx'����5���|B�
������/%�������́�3Ҽ����1�d��^; ��+���W��~x_�g�/�|S�K_Z[�4��]�l����k�+�� g��S� 	M���u�����ʺ)Ħ�?.�>�+��k���܉�,�"�7BInȒ�8�����ٳ:CV�TY��Z�{}�������������n?�����:��}}�O�A?����5�q��G���9z���;�Ϗ��l_�L��O�W�(�S�E登���~��q���w�`�����-��kw�im�[�$���6N��mds�8�#�_�� �Lw��½�7��1�������s�_!RP�K��v\���h�#u.d�#�Df�\��2�l���4��$������J���jzG��b�|%kj���4k0�Ό�Hq�y�M� ������ �#T�4|~D?R��g�����|<�-������l�!�&Rq�F�`�*�nN�K� neIʤZj�נ��n�I����s̖�R�+ ,���#=	�+�k������&}F�ȯ������� c?�Zw�]� B��I��Qmb�ʚ]��~�3]���w5��6��|���	�oZ��r��'>� ��[D�� ����>x�᭿��[u�>��3[[1�&��\X�r8�����������5�<i����({i5粵yЀC���c���K���%��B��>i���W�~������o�s$lYca�Ҿ��W�4�X���"��]��}4�����<����1�)N<4#��7-���]_}OB�;ǞoC��g�_�G�M�񧌵M>��H�ԭ��{I�'�#�p�J��ڟź��?�%��O��vռCqym:�w3;n�w��S��_M~���mg�_�<�=���%�ڎ�$����H����={6+���7�O�1a�����I�]�f3�1���i[g��_"*��wN��6Ŏ�R� !Mo���� *s���!Mo��C����E&�(���2*�q��ږi��c+���#�־����c}O�Q�#����V�c�M�C;��d'�'>��n��E|��cb�Fs��C83I��ٞ��1� �D���{|������?f.~"j�������|�q���_�݇�z���׊t�>���(?:Z3Fh �QI� /�7��?Jw���������>�n���������ϵ���� ����s5�p��	D��\3V�*+���f��o
W���4������M����A�]��@��s!�t�9ÎI��k�� k���ׂf�x������+�jV�0kw�Tn���m��ֶ���M�yz_��~�qKmcq�ml|�p0?
��S������6��O�������Ch�E������a���A�e��� ��R|��>�v�O����xC1�5(Tv�5��*�V�2����?�}��`���}7�5�Z�%���>+�1�U�t�=OX]n��O��a�#w"�}
�־e�i��"FSs9̊>��lEoT���	r;�R\x��l�?�W��`g�ty����ۜw�[m�� �;�#���~�}� �8����?�����G�ˤ?��¼� ����� �W��{X)�<�� �����_�����G�L�>������A�_�k�����K�-g�#�ղ��o}�L���sF� 29�NM|q���g�� �#]n��m��v2ȁO�U���]J�I� *�����Q(�ֲYZ�e����q�k_�z����/T��ċk0�販)v?�@ �U
���P���c���}�Y��͵�n�:z�io�?]Ns���<��u�[x���O1��'�4ڸ� r�zW�W�|^׾!|x�ϋ|S?���<Q�� $@�(UF �W� 
�_� �!� �k�e��M�JMy&��cӍjv����]7�+ϐ� ���4·�������X� f��̿��C��� �}�3^��3��C�/���s�!����p�v��6���� �[���|���_�F�'㟉�ψ.��	�����\L��6��n=�Q]|����I/4���*��v�*;�5��D�L2;:��r���U][�:o@�5ni��{�I{��ieo�3�������������>��}w�N]�_�O�yC�t����9����U� �+n4���i��b� hO���ϗ���󎕧m�C�w���-|/�_�S��ׄ|Eঔ����&Y�~�R�
�r�bxu!t�|^̼���v^��E|�H­��+{��~����U�.t���9�z��!'�DÞ�a_t� �A���i�����6�}�[I�T7	����Ȭ��|Z����c����k���$�S�.�J�rKh���AOK���ƣz[�o6L�*��q=7��y�`��>7q��e�f۟�5�����'�����OƟ���_���/����k�0��-�� ���!P�1��UUI=���R�K{ZJ ��O)�r�1�W����N�G�Q2����� �
Y�M_�>��ó-����m�"vl���7)��Mz�ۛ�~4�MgO�Ԟ��!��r��t�+��q���<�+��,�w�9M�|%1�OL8����?/��5���j�~F���FC�ug�^#�0��Τ�%�(��M�^��*2i+�}��_~ښO���x�ֵw�k�St� �U�f!� ��ÏZ����� ��I�`����|I{��/�׳��.#��CwD�OB����ߏ�򉟄c���� �sW],��[�ha��m�[mn�{YVnR>-��rO�)��[��9��?��?����o��U�ǚX��(��������o�?��n�ot�4+ǒ�%"gR�C*�{_Ϗ��M/ńeU3鶿���D~ ؿ��<����g�AO��� �"�s%�'�wbz��0��P� �'�o��X�k�?f�(ڇ�y={|_���^~q��� n�����OZ^)+�:D�i8��~Rm�mR�� '�Kǵ'� ���KE f�
N� �SF�ڼ��	���1� ��/GY]��c�$J��}x"�=�o�)���n�u1ub��fL˽�*s��5矴7������xö��j��B(%������Ğ�j1�{H�OF�eF��6�^9�qX���!��I�9�X��|ЬBH� z��3�+��ԣ���u_h�'g��k[����/aI8⤨4�K�'��2jz���
?*)x��A�QG�G�@��&h ���1�@�}��h�����Ѥ�ҍ �7����4|��o���d{Q��E�9� �������'�i8��� ~<я�~gڀ���n���@I�)wC� >�� ߵ� 
��J_�~���?����F���?����L�(�?Z�sI�b@���#PG�⳵�q�8�t��������g����<�	i;��[���eo����+�[����`�_j.��ͪ�i��?����_G�x5�����iQ�A���T���n������ ���g�1�L��u����|,��V�gͳ�����K¾��{��[�����_�^՛���J�(e� 0J�0���z��9�=)b��}m���{~��٪�x���7��Z����g_t8$��|AuX�sE*� <�s�88���:��%~��0GϪ�(�d���i�>�9լ/o,����ŷO�b%�J�d*�#��������o��$��T���'?�<��d
����˙�;�kk��X�sy�S����$�B�� u���S���� \��
k����_�b�(�������?�/�� �;�������� ���A���H����� �����������ʾw%��N�OC�� f�(���y={|���^'�0�>:��O���ԯҼ������_����R�IF}��:C�J?:8���Z (��&�΀ h�(���Ɨ4�Q� �-'�q@�jOz8��Ҁ£�R}"Hn��L���a�����Immu$1������=x���C�	��'���ۨ�A�Zyr	a����3�¼� ����~	x�����I�B%\��+��]�.z���{[~Ԟ;�ᶳ��d���oKW��r�`H���Ñ�C^s�J~О2��_h:�����wQ�_շ}��o3��pNZ��bq��"����,���[I�Y�˷h�0�Gl���-Gcn��EX�Y�Z����B�p����z-�⛑�@��sM�=M����ԜQ@�FO�z�dz��&���E .i8�����(�( ��Q��K��p� "�h�����/�P�5����i��� fZ�� �֐��*��r��KAQ�u�S����,*�� �Jl��F�������Ɲ�;�͖�(������k�o�(ׂ���?�'�	x|��� �-)B�o?�+㢨�^��g�'�k��g�t�^x�X�EMK�W��=��+b@æz��� lQ�)F���RM��{i����hJ�潒�~M�p���]Gu%��ж�����s��?�}��� ?�韄����� C�����*�-|��6ӵ�#��</z|�: �{�z�����O�2,��Io��� On���`EtR�hfn�j-��i�Ӷ��J�jG���b��?����o��T����$�B��u���W�qb�(�������?�/�� �;�������� ���A���H��/��� ������������ �k�2_������=��]\x�V?���ν��+������� ^M�ν��)�5�f� �o��� ���cޗ�h�c�N(���(�� �h�h�h �h���Ҏ}(�֏ƀ}(�ҏƗ�Z n}�}h� ^*��k%�q�~t��l���*�n�^����a�����"�>��G�sY���t�9�/�v��X�KI�%W�� ��t�y'���~+��|e�i��?j76ʉ�X�,��~�[h^��
�o��� ��5oJ��须`�#�o$כ~ҿ�W�_�� ���a�K]z/i�	,漻/m���8�Mz�x���,�{��s	��z#�+��f�
� ��*j������/$A��I_py��s�G�3�E4m4 ���ϥ� �R�4m���Eq�@R�P���R�gڀʏʖ���J^}h��J(�֊ _��q�M�0�.��֏��g�>��� ]������Y�[x�O�K�_|׵�|�'U��i���Uw�e>˸��?�?t��ˡk�t�;lg���J���S��ڿ;�q�/�J��L� e�#޼��I�S�o���m�O񇇡`����ف�X��Tc�#���#)�b��`�h�֥�Z[^�k�z��B?�����ߵ��M?�
<S�+�yt،2i:\7C�,l����� �|������ �%>!�7�?�$ƾS����_/�u���\���e�D� 趨Gݎ0p��=�}m�@�&~w��?�9���K.q�Y)T��+m��^�β���7݋��'�����?ʜ�v���S[��� *�c�,QE��x� �#����� �'z�w�.q����� ���A���H�����'z�w�/�  �����_;�� ~�n'��� ����-h�f߭{��{���y_�n#�<C��������8�V@��+�ͥ͌���m�Ҙ���Q�4q^I�&ih�(�Ҁ(�=(�Ǝ(�Ҏ=( �(�Ҏ=( �"��J8��>�w��J( �QM%�2Bڂ����!}O� _/�Qͧ˪I�,�!p�wN }�������'�� Α�'���1y8�<��>m��s^k�M��J�  �N~!�� m���jRh2��	� 6|�}�8�G����3��Z=������ ��R�p����A�6���l��?> �����|O>�n�u<C0p�{n8�ҽ�=B�	:J�_d�S����%�E���������ڟL�S��m��V�jJ�C�
)q�F�c@���F}�q�� �4�Q�OÚ _4��!��'�M�D�7����8���m� ?0� �b�'�i*�Z� ��?�أ������(5w��#�9����A�z?/ʏʏ>�gڊ_(��)��pn�F�?�
1�V���~�'�s�>3��[GZ
�ď��b������6����5���c,�I U�I���	�b�Z��_I�I.��YѾĸ�e%O�}��׫~�W�z_���U�cn����m�Kt��o��FW=q���?�E��^4��K*�a�e�EPs��c����]:��a���\�V�{h�۩�S�:�W�c�����������>*�����3Y�g�O���fP0G��׮||��&~�[o�j����<'���5���|6�Sǭ�Q�Kr�a}��o#�|i��:K�8���O2lWvW�b1�C��NV��m?5�&�(�w�^����a� �I��5��}�?݋��'�����?ʾ���QE @�?��A� �~� � I޿��_#��wa�+�%�鱾
��H�V�o�̑��&$�9=���𽌚�VdJL���P�zrv��d������>��+��`�}B����P�
�|T�a�G�4�*�4�>���#��Q�c���EOmZu;��劈�qE'�\��EP��ǡ���h� {�����K� '�G�G�G�@	�u6�m .=�:
6������4v�Hѷ��2�����U�gբY��#v�zd�n��}�����:}����_]Kk��H�|�h�1�kʿk���1�,��R�>hZ.��0���D��ʹ*OBFG�k�K_�_5υ�9���ƽWK��ۺâăi@�S� �zW��ߴ/���l�^)���k��+\�vH:�p;W���⽤[�t����)ӵ�8+&/�Y�;��R[<��R�**�TQF}.z�Ԝ�T~TRn�P!*?*)7�(*JZJ \�QI�Fh��� �<!��2�O��gk�xE�̖��D9�pN�k�o����\Ϋ��
2 �_�9_~�����1�hz��G�Ȍ\��n�ֿB�e�˜�j'�N��_#�Ԝq	E����zu�_�e/��-� �� ����� "g�@� ��� ���� �\�'�� _�����.�_j���+��տ������������~��_�?�i~!�QIs���H;�ǌ�"�C�����~h�g�;�k���U�)�@�i�=+��0���9L�<2��������>�f����+�9���4����Aϭ/�R`�R� � �Y������?�%�?��y{��n?�%����+!���u�����
�=��U�]J�#�X>� ���z=��ď�I�Ku�� ��I�mB00|�H�H<�V��j����W�If-�|#7�.0>��� c�_<+g�;/���-ғlڭ�Vs��|�$ �=�9+���r�NiYEKF�-����J����J��w�k�?�ë�i�bx/���y�-X����e�� t��c�hæ���kk� ��_,|j�3�߁s/��!Ӆ�{K�9{ir�$\�n:g>��?���	5�%��?ߚ�i��P������}�D�9JN��ů�b��?����o��T����$�B��u���Wўyb�(��oO�I�:&��/	ܽ�����A+�r�gQ������A�w����I��u����Cє�h��f�cjg�:����K��**��煯��ɿ����,i�<�ov f�,D?��2T�z_�댽�]v;��k�n�m�c����})O^��= �>��;m@J_�����̃�h����T�^٣�ܳ2��#;�m=Mgx�ƾ�kqoi�},o�Ž�FgU�`�w>���R�\J�}�a$�G�%�Ռ�~x��¾4���ỗ�z���ؗ}���
)<G4��џj8�{��z8���cڀ4��b� f��=� � ��� �/�q�� A5����� ������ ���|,ks���~̿ܖ�i;���+�{Q��fy� T;��>� �a������1+�k_��� �!_����x�%��u����Ak�J�OeI����.M@�"Ӕ��+��⾻���|���9����7�����x��:n��`��>bbp	�񭯆����-�#������r(�����Pܫ n��Ey�ƨ��.�?3f|S� 	�������"ӈ��G�k����a��#gg���1�=k�ߴg���Z}��?c�?��He��mC�0pH��l�-,ڍyr����O�f��ʚ��> Mj�GTU�V~���5u�km$W����o��U��__|��o�X}�=^��|�0bKmVG��� 0=���b�;��X�"g=¹���i8٦�g]F_Iuq-�j�s��֔���O>l� �zt�V�̂A��u���.I�bq�^&a��P�ʝ9Yi۱�F�%��O�|��k�����+'ئ�����ϥ}?7���M,��,G�۰o�8� �u�w�q�Vc��I�����W�Z�\D��;��1QVG�?��?� ��� ����C� C���e���� �W�� ښ���5ڷ� ��Ն���I~�^7�����	~[�z���P\�#����2�5����T�E��9� ��w&�{ �\>�ڮ��뺎7B��e�2�8I�H�nŖ�6������j���rt:���hS��J��F?r�J��[9������J���P��4��W�r�?�� ��~��u�n��j\�7
�� �׿�i����	h*;���������C�͆�m��-3���Ehͅ�hز!�Qǵ}��� �:O���&�jk��	�h�(=�������� �)o�5�|t��/J��֗ᶼ��$Hc�-�FT��5�_� n���EMO�����Z�Ϯ�z���!�
̄�8���Ng��*���Ԧ�-��qvZ����=��+�v�ꟵG� �'����ۼ;%�����;����cV�q���c�|����� ��N����Q�z	e��T�l/�7J�/�u?�9�� �#��\���ч�H�m�bB 
�H�:V�����&~m�|�gǹy�^�K�����X�)ɸ��n�.���yFR�]�>.~/hS�
k}���No��)��5��}��O�EPc��� �_D|� �Cp?�(��W����� �_D� � �Cp�(��W����Tta� �w|U]wP���7s{�i����m�����-���Z�8<0+�L��9|q`W�IE88�d�Tۯ����y���j2Ŵ�⾊��:���v�� 矚��cֵ���"��G�2����~ןt�d:m����jϦ����|�+�>���le�ĻF����f���}�X�����������p^����I�ϯ=�&MQ��Y��<�w>q�(����/�|�T��x-�D�K�x�<��3�#���*�����*���u�z_�k�_���uIVKXT���!�FV��
�o�Jh�)c�6=9�h�K�Rg R�z� ?*?*2=E��ʓ����Q@H}sK�Y��K�$]�[ր+v����YO��'�Mx��>:=��/i~6��m<1n�-���*��Q�<g5�鿴'ËEf�ڄ�/��GҦI��5����f/���ӌy�_<Z�>ϷX�����>��B�P�m�JZ�ˌ#�Ǖ��8�(��3��B�y�t�Ѩ5(���;~G�%m�ӗ����M��;U�+ dd����u�S�#� ����%��{e��k�D$˕�#�?ޮ[�	������.k���_�����V���IU���RG�J����i�C��x/[�5�|E���voP$,yUWR&�*��Ez���7ë�H,���5	���c�[t`���U�(*�%iuK�z��ԯ������>���~�� �E�����]|�� ����w�_o�'�H�Mk��8����H��Y�q85�������X� �8���Զ?�w��"9��,�-ю�� ��������6UZU���-�Kϱ݈�K�%�`� �&u(ou���+�e��3PWt�$�'����_X� ǔ��~�q�?�5�>��|�� ���{�5�_���#��g��d��@�b�m����^��i�� fI��v�K�I���`��U�Y+t�N޿��Ե�L$� ��O��a��W!/�}Z���]�v� v����^��GUᡴ�O���jM��W�t�z6�Z9�s���O#����h擏j;}q@��� Y� �����WA����s�J�<���=�q�6B��@����=��z_ƀ����<�KZ�T5�s�)�uҏ�}h*;���*���;����Fc�=>q_i>���6�×Z��>w���8�J���>A�����/�K���� ��_j2!;��\���@#���7�tX��������[�V+j�i@Q��l�|޽}k�jg//Q�P��U�k�%efߙ�G�}�;$~�H��:��%�i��D������@=����� �&�� �[_�j�_�S�s���=j��6����B�K��V�%��D,`�A�pG|��'[��$��v������a]x\���.Wŵ(�gn�SZ�:>ŵ{����ؿ�!Mo��C����b� �I��5��}�<��Q@O����}�"�J�~������̩pya���_=.6��޽/�o���>�Ӿ.�[ƞ&���gsᛔ��* Fˏ���^^eNUp���Y������ �c�����OZxW^x�c���g""G�1��_~k���߱�l´���%� D~7��c�d~,�S�� (H� ���>�W��������%�:\�����&?y��5ac��f���;���?dn���*����� �(� ���#�3��� �(��/������Ώ�D�K�o���L��u���ۿ��ӿ�?do�&_�c� �� ���#�3��� ���S��Ç:>a�יg�:����t��s��o�N�L>&?�ih�i�=t� �?d�&�a� U��#~���� ��]��o����~zS��Ç:=o4���'�)~ե� �b��2� ���G� ��'��� ��� ���G� ��'��� ����P�G���K� �ſ�Gڴ��[�u�_���� �#|d� ���]���� �#|d� ���]/�����Ù���/��� �j�� �1o�י�{�#� Ѝ�� ��t�{�#� Ѝ�� ��t}N��� ��߶i_����=֔u Y�U1�������������6�� �����df� ��(� ���]?�Udy��n4��j�Y5��K{)Xn"E#lb���#8��<;�O���"��/����z�"���}�i�ygl�~�q�ג/�/�86����S�ܼK�q2P��#�G�߇z��K�cu�cH���x�W�[!���br{v���I(�jK����Z|}�9��].��(Ŵ�
�ǥVN7c�U��b�W�(�a���Z��4���j��� �_Y�¼'�ۻ�y�j{I^���e����?�0�C��95�U�ξrd���o��>���j?�2W]M`�&�ď��oO�����O𯂿���7}��ս��|s3�gW/��+�`V���xL֭����n�0��P��� �냃�^� l��i�	�rN�:����@��z��
��q��0�ѷ��OJ��S�hU����H�����g͐���<��� 
�=d{;m����~:|~��f?�	<Q�xx���j�~���;�E�_z��M7�,�}�U'���W��U�[�]?�`���ե���ӊ�2L\��V��m=�](�^��~�?���i�*�?�5O�O��$l�1m���
O=���F-��
}ȯ.s�B9��?������'��b��/�WĶ?5����n�a���Ӎ,D�� �yU$�Sd��n��y7�k	����_H�/��|m����o�<%=�~�%���\g~��O��?�|�z�����!�W5�� �r�'�?g�hzG��+��D7񒤗,�>�5ɜP��c^f����'�(|G�J����|W!��I<�P���s3k��Y�Ґ���]_�e�;�~�ZƳ�ڵ��֐$��)VE	����!��c6�v�}k����iBr��OqN��&����#ƿ�%k�	\[G��]�(��wy�d��p���k?��U65��o'�=0_S�ƿ�G�O�:n��h7Z��Z��ML�d`�@�_1~�^$���w��V�i}5�V��J���?:�0�J5��0�߹��J4Ժ�mƹ�8Zo:f��=k߼�|H����Z5բ��ݲ������#5�n�hC�z���ӟ�?���3���=����l���ⷸH�Yt��^e����Ҿ������g�^<�������3V�0x�G��q'"2�+��Lj�H�!޺�����(����b�.������Ўƹc޽��<��� 3��G'n�K��n��w����0z\�Rn�?�;4 ���)k��nT��kD���m�['�C$��6�bGs�3����'���W���-��$�G��� V��8���'��|tK�A�x:	> �?Te{�yQ���PL3���?�Z������?��U�}�/�g��t��/R�յ#�c �B���l�W��?��4Xd����|���2Eg��hx��_��^2�N��Ui~[��ѯ+i��º��%t}=�u~����w�i����5�h�t{9�I�Z2�6;�8I5��E��_�*�#���<ٯ7�?b�  ��27�+��� P�B���������5����-�'�� b_|�����K���O�\	b�P�3@K�>�ׁ�c�P���nRj�v��%��[�7'��|r�v/���S[��� *]ے"z��O�H�����}��(��E WU>S;���'�*��$6�� $�FIF<~��?a�ؖ���Ԯ<Q⩮t��l�l�k ����Qs#�f�'���֓�&��l��~�DEk�tky����RI'�xx��jrE\��]��v���|���O.2�����{Կn��\������?��?>3�fF�֑g��Ŗ�J4���;[yd8*�1��D��FpOJ�~���x?����Cg���-���[�*�+�,��F=��px��ݙ�J.�!�и����o��� �j��4��L�'�u��� SGۮ?����b�'�П���4��� |�u�	��?����u����y���Z ����oΏ�\y�:��Z9��	��q�����u����y���Z ����oΗ���?�Aϭ��� n����5�� v�3�Z?`��QIK�@%\��������6�7V���� "Ȅ���U:^v�� ��&���I�����~�ߴ���#�^����K� �V�aյ���
O����t�'��D��mo�?�� ����mH��tʨ=����x?Fv��y�`G�� ������?¼H��**z#�U��}�� ��y_��?�XM� �UK�'�?�$���ڏᦽ�� �]Sįp#� wq8����ѽn������h޷?��� 
�����2K��)ք�?J?dφ~������~1x�pkZb����d�ft��	$� ��.�#���do�i�O.N�f&���]"�U�y$C����i��l���+���9Jswl�5-Ћ��g�������
��ο��x�]�I�i��	$�c�<�g�|���R%�ơT�J���&<���n��~=|]O�� �O�Q鍢��	l4�Hf@�$��5���Y ' �5#6�,yjOֵ�8�GdL���}e�7� �B�����M����E��%���.�n��ݹ�W������~.���*M.#��,09Z�㸒5NsLf,ķ-\��Օh�Y���TH.�E��X�a���	� �w¯�~�|�5F_٭��#����##5�^�9��U
`/J�F�**5�T�:n�����O�Y��Wㅵ����͉�q��vFX��GX�z��JORy9�z����������j��h�����9Hde���r����	~�Z�;�����ѵ� ������ �#i� }��� �'�I��<W�;�_�u���7+mk4�B,ӆE*�V,`��Z��� �sA��1�����q��FH���W�,Τ#�8(�7c�8x�D�|=��a��B�����[O� ���������/�ԼM�x�B�W}��χ��-GV�����c����o��P�hVfU_���_' )��P�kT�4 ��w��6|���C�A*O�H�FjUf^Q��Q־�� ��x#�����H�-��
������N�-��<��1E n
��徘�W[���c��y����
\3�cw���O�^)����=����� �W3�)ѯ��d
���e}��r��oBsƗӹ����U�}J
�rZ���&n?����I�����ǳXCq>��]�kZ�h<��qXa����߅c��z�W�c�W��ӴkO�������4�.���i%t%��s�b�lF:�|��mo��
R����9m�Z^2�wP���
���pUYH���U�q���3��ri�;���X5�Cgu�H*�:���j�r���]��CW�o◎M_M��-��_[�o�D�� ��p��x5ф�!��%�ȩE�]��[�o��ߘ��>e���?y�d�������:�pi�A9� �/�+�ܳ���_|� ���y�?����M`\\���,Z���i31�2N����#v�_zn��_��"�ZI�=���k�'�
Ѣi�O�A���KHa�Լ<�x�ZvI%Tg�R��G�~�^^-���.��F� q�W�o�9��������?L�i�t��C��UV��Va�7Y�	��~WMκ��gY�,��s���T�����<�����h� '�G�K�1@	�Q�R�P~T~T�� ���.(� '�G�K�1@	�Q�R�P~Tb�b�����b�Oʀ�J8��b�Px���Jv(� 3�_ƗOʗ�oʀ��N� �{яzw>ߕ �{���N���h�֗b�^�����Kᷡ��� 伵�}�c�^7��S�m��P�x~e��$$F��(��i��Z�R��� �+���p��[��?n���-ݣ6і`���W�^(� ��| ����-�\�]�i!�O�:��2s��Z� ��A�r�]��xTׯ"Xn�	ĭ$�RNN  rOJć�
��u+����9<?_��GC	����sYv���R�Z3��}�G���]�?���^�|G�K�wW��������w|q�' ���]i��AC�m�L8��~X���
���٫��wQ����8?��^��
U�Cu��3���q�Ilv�s�d�������>_;~�ί=i�I�w��TI����&P���4/���3q!�޾=��>��|l��u�ڛ��|B����yon4�,4��Dp���y'q.ğҸ/o½�7N�O��y�V\�
�����xd��0=T٥
�2��tLp����]����� �`x/����|;�ĉ��o�WYK����	����L����J��� �E|l�E�g�>^��4w����w��RHXpAB1�Cz�Rպs���
�R=x;�0+����� ��,��~��(!M^=N���
7�[Ԫ�'�q��ҡ&k�G�
��Q���Fj��%��|'�cnѨw�*�t��rd/� }+|���b#n�U��]Ϝ��⊿���#�����]�.���PK
     �8�Z"9��T  �T  /   images/0b0a0ee7-c404-40e4-9217-cd21fece1ba1.jpg���� JFIF  ` `  �� � 


		��  ��" ���          	
   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz�������������������������������������������������������������������������       	
  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? ��	��3Z|�+���U��x��Q�n���T�l��ݨ��|rWي�p�x7�A�_L���3�+YӃDm-F�sLS@2�b��a^���!�VW�L~R�4�mR�{K�#������	�:H�0��x �A�k���������hK����o[�[I�����{��W��[waɯ��*_�-#��6��ir���]/�?T�.)�w�.{�Y3�H���SU�a��d�ϒ�������k�,w�G�I��3�s@����g������������������������:?:Nɣ��h:?m;��>j:�Ү�{��� �/Z��>��O"�d�́���qP@�iI���)��~uկ�߉�K�^)�8��d ~;i��#� �2�� �� ��>ޟq��y�?��/?��Y� 
s�aM��O�]��2����o��3�ޝ���\���}��^ںč� �W��8�Ua-�����|�_Ɛa�A�=��q��~�"��M�\�*�,��d��&�7�ߕa,E�TI�2�$��f�>��}c�m�zM�Q� 	���7��K�8���9'������ϡ���M4_I��Ķ��M��|gsӎ"��,j&�8I+�i�f
���(彨e��<�Z�|	�߯��]j��\G��ʡ��#�ƶn��Y�|E���O��ғ�='�x������S~�:?���@���V�	�h�M����M"4�`�C�� ��  t���>,�>�|S��ʞ�4=Tn����1J�rF�G88����~�|��w���U�l�� � ��J� ��� |5/�$zG�T�&� 
��>#�k�"��/�/�V��Ff�\�Z$�rUwc'�����v8�k�k�<x����#4�:4Q>�0u�=@�D3	Տ=.Y.��^�'i&���7���.N	��~��׽}Y� 0��8���^$�tOϮ�f+��:�� �wȮ�Xe��|�0g�����]jJmns�<��f�C8��K��#�{ h�������i�1"���{hf~�� �$� g%��5O��"ӌ����]y�V+>D� ���\�x��H^:����J�Qx��p_�烮N�2n�;��	f�S_i�縹Iח6��1���j�w� �����~4�>8�A���6�X&��-���mQ<�>�+�b�_�;�W��+�.��]x�v�^~��]ɪ_[�	6�{c,{d���Z��kB*[���+��_��j� ��� �o�� ��W� ���j��G��� Ǩ�(� ����}������<�i#�?eoڛ_���a>��Zc�ڡ�kZ���� $*�y<p{�����
1�#���V���~��$��A"��DG��������{ox�⇄4=Ķ�����m�j!����,F��bx�{���߲���j�~�'��j� �X��a=�����J��� ���6�u�S����3����v���iO�*��t�3P����'�<W:��E�6О��T�8ۜd�`�a��]]\��˩�׎d���f��$�;�7$�JD:jI��Ztu1�}��5
��	W����v�g=J�zt��S~���Z>���Z�I?*?*���E���E�	8� f�)�h��z-^�4]_�RO��-c��n��]��L � �M���Z�T����w�v�m�B?�?� G� 9� �k�?��� �V~���c����@<q� D�Ɵ�%�� ���t� �m�/�O� ���!�9%�����#޷� ���o���"��@<s� D��_�%�� ���C��%�����#޷� ���o���"��@<q� D���&�� ���C�rK����V�|u3O��4f�4� �M`�F�}Զ��K���v�cv�9�oA�5Q���qkp���&�huH<���(�g� l�C.:�?ʾ����-�������0�4o�$��m�mJ �!h�\�Wq�<n<W�|��VR�_T�$��/�&���蚗�5'��R}�K�i�ثn��@�g�y��S���FԷg����� j��.7��~�� ������;f��b=��~S����R�]�;�?u�@q�K?�r�?ey<g�9Y��<E�o�M�x�L{;4�F�f*����ۚ���s�b�ᇌ����w����8֒�G�:}�� C�)�')[�� ��������?g{��"�����X�����L!F na�Y�&�|*��~#�ӿ���-o��:v���-�ӭ�/%�JYF	,�E �H#�x��c�x�dmCട>$I�����#МY�YC�1#wL��]���������j�J<+��i.4{a��2[�d��v��N20EV��R�����K��NJ�����Z:�d�[���]7��uM?ǚχ����Gr�O�,s��Y�ҹ��XJT����>��x2�W�<i��x~�t�j��%��$�Zۿf/�?Z���.� ��3��FO�M�x�X��}s��־�1��I��X�8�0�#�8��=��3^��Pxoƾ��}��@�E���J�𼺥�����Ⱦgr�^E_�U�$�^;!(����GJ���]���x�U�ែ�k�>��qk{�-���RFӜs^+޿d�C�?�5h>x���z�V�n��Y��3f1�8��ԏ��Y�;���r��w$���nX�P;`�b��� %����X�x� \�VmϘ��Q�%�r��*��p�3��Im|�������G���l�co
}"�@���y� ������~"���mf�L����e�}	����7���#��"Ԥ�t�V;���� F��#��>*��_S��O��=����ľ?Si~�Y,�%�K)�Aڻ3�'|
�c�X~�3i����J�	�ڳh6� f��y�v��:����B�$p՗���'������Ӫ�Cu�zO�ࡿWK��ǈ�Kw��h�/���s_�^ ��[D�
&�ipoo<�7m̻��#�}�����,�?�4�bp�t�O�� b�u/���qѮF����B�x��ou���+F9GQ�6܁�<��<����et��������Ϟ{�/�%� /���O���p���m�� ��Sk}�5��V�U ���k���
��e/��������Z� �4ٛD����J��H��ۏ,�|��5���P�:u�̥|�efv?y�����t����� ��qU���=(�PH=��vZw�����<gsg9���:<��pA�C��5�����s�/�����\�t!�M#%NOdC����f�P���)̢i����W����8 n�� ���*� �������=片���Ͱ�(�	�
��~��}��O��������R��$S�ti��r�1�{��B���_Krs���v�*�I�85�W�a��-N�T�4g�ǟ�*��7z����'�&�*�ɝ>9
��Y�Pz���2:��g��W����z׊�Y�kx�X�徸��cA�B�� 
ȷKM?'M��Řa�Wf,?A##�� *���!���fu*��?��z�揲���� ����
��n}�s�� �>.�{�7��"hJ����L���C����U�?��إ��&�}��%�B+��6Y.�d>A��d �����Lr+�᤾�ď
��Ğ���Ƒv�Z���	M�y�EF ����+ܿl���?ڷ\�4�j:G�=$�.�,)n�W�>���0أ�Q��n�ޯ����*ʛm��}��5"�ty����O�^6�4�n�TH�Gm�.%b��v��;�]~�,(��L�+�?fY��eU� Cbz/�ۣǖ8�NeZ���J�J�k�Q�e�(�� �G|+� ��[���G�(� �����j�q�qF?�+���/�K�� #_gO�Q��W� ?:���� ֣�¿��տ���u8� 8��}s� ?�����?�G)� 
?�g�����������.d�q�� xV[��KL#L��}���G2�⤹eU���������>?���� ��)?�?�����X�R��Y�z�����ErG���gG���Ƿ�:��U�3J�������e�jVq�A�d��ᡌ��b���^��	7/���9�fjڍ΢|I�Y�x�Ymc�J#���Z=�^���,{~g� �����g�� � ��� ����� C�� ��� �Y��z���J?�|� Cf�� ~R������.H�9?�nώ�>k?����������� 5�� �,����S�����>� ��T� �)G�������r���_u+�]?M�޷%��l�@ſ:��O�_�k�b-[�:����Ȳ��in�?�ұ�+�����C��wڶ�g�ȷ�E���N���P��Th��$�P�1�ETq5��ͯ�����<�Z���4��;h^��A���3I*�xO+�NA�+�����ǃo<Y�Ae��%�s<s#4`��p�+��㷃,t�:�_��E���G��������r1�䟶/Ə���^�~��x� I�5+�u�>��&������'�{ts\�8h�[3	Q��g����g1��C�)*+ ���q���R�����<�Y���RE}_�#�Xx?�q�ş�V�� ��1c�� d���k4�x�Ճb_���k��y����_Kx!a?�J� y���'P%}�8���g��;*j)��#jV������~]���D~�S�0~�,I��g4�~џ�%�O|},y����5��N?�F�,�1K���zg��o+�Zt(I	�g$�t�������b\p�&�MT��q�g�}����4��x��o�	*gh�B2s��5sZo~п�(j�~;|`׮�#�-�����7�ɻ�J��o-�'�LW�hrxn_�&.��e���GR�y�\ ��[�$���z`���_�g?���Hѿ����-��lִ#�)���%kߪ�	%����ل֥�k�Z2��#�k�{K�׼E�i����>�s(��Qb1n����V&�� s�z��t�I5�?��'���Q���/��W}���_Z����~<x/����w�x_�q��I�(�Mb,bFe�/�<W�ע�uO�)�
�|,�W�������3o�2�J�ֿ=��VO���EW1B�ҽ_�{�q���)���O�-|ioh��yw��Hc'��(�z����
�)�?N����F�*����������+���r'�ċ��Ma$q�"J���֪j�?�f$t���J��L-ص���9o����Ͼ1U�_��	���5������Զ� �=�fk�F2��Z@��G �^���~y������ ß���U�iƊ5�QCy�n�s�ߥ{�x�����a���Z5��kw�im�ۙ$���6N��mds�8�#�_��dwi���%� �&:k}�=:y��}��jT�J_W�����G��s%���#����LdD)q�y0I�+����.���B���Ţ�J���,/�h�a�������^�� ��ep|��F?"��k�7��c6�|<�-������4�v �Iǥ<<�a+*�nN�K� neIʤZj�נ��v�I�~���q̖�R�+ ,���#=	�+�{����	��&}F�ȯ��������cO�Z�}�B��I��Qm^�ʚ]��~�3]���w5��>�Ӽ!���	�oZ�0S��'>� ��[D�� ��~�� >��ᵿ�<Yu�>��-3[[�1�&��\X�r8���!��������}n� bi�
��粵yЀC���c���K��<%��A�������W�~������o�s$lYca�Ҿ��g�t��\��!��wl��N)��5 b w�'5�x�t�JL4#��7-���]_}N�S�y��?+>5�t���^���<c�i��
E��m��O�?$�3�x8n:W�~��,�~!�/�x���6����i�R����t˼�R�Z�g���_��?
�_�e��I-��t�$>�2D|��>��ٱ_$|p�i����	����M���1�\q�H(ԧ+J�=.��V���3�G�ر��_�)��{�No��rO�)��[��}�����F� ��6�ʷ|�����V����d� ����l���S���F���.�o�:�ذ�3�M6By�s�����z�Wά�6!��a��=D1S�.ppvg�~��Q5��o^����� :�ً�����y={t?���_)��|��wa���sA�G5�!ϡ���P~t�Q@QI� /�7��?Jw�� /�E/�E�� ��(�}�G�G�@	���U]J�k8�	��T^�$f��TWQ�42��"��=O�h�[o�s�-�cuy��M����%��C>�d s����ח��������^.���Yh>!��W�ԭ�`�����1ۑϭmI�3����.��� ��]�I-��q��d��9���+�� iO���7���ߍ>6��<7o k��EHdPTg�s�W���m��� #I�t���KY�w�3SR��GhCY[���h�*�J��WܞX1H=�+�ٯ���=3�r�W���Z���Y�z��V��}�����pc�Wn��/sO�q2�#�1�dPq��r�h}b���.�w>���� �0V�l�)x�M�����:� u��8�Ҷ�H� �x3<K�%����� �q_"}�Ϝ���?������^{�W���� �W���h)�<��$�����_���A��O�L�>������A�O�s�����K�-g�"�Ͳ��o}�L���sF� 29�NM|q��=,��b_�k�Ѻ-�Qn�Y)�*��VR��V�?�]>b���J%:�K+S���=Mk�oT�мU��:Bx�mfU%.��$j�W�?��׬u�o��6y���ݱ�C���]�-�  ���|�;��s��x���O1��'�4ڸ� r�zW�}+�>.�� ~;���ž)��_W�(�k� Q*�� p+�� �s�ϗ�D_񯋫��%6�)5�_}�N5���G1�WO� 
�_� �!� W�h� �s�� ϐ� ���5��v7�|�� �W�����9����_�O��Ox�Q��~��O�kCzu�r-�p>h��+�� �s�� ϐ� ���5�<u�+�{�޳�;���^[�K��8�� ��g��+���r�$��K��L��i�H�#�5��D�L2;:��r���U]W�:o@�5ny��{�I{��ieo�3�������������.��}w�N]�_�O?�}C�t����9����U�+�4���i��b� hO���ϗ���󎕧k�C�y���.|0�a�O��ׄ�Cඔ�t�2I�g�߱��B��\��+�ئD\�Ə�/;?�ݗ���_-QB���+{��~������.t��tI�Z��!$yw0�W�� �P]~;��?@�������i��t��ĂA#9�_��~�r+/�.?�r24�~�[|8�����~3��Uc�[D|�b
xha�X�oK|6��Ȕ�R<�'��÷�/��GF�3L�<��s�f��� �O�3�W� CZ�J���9���>%�<�]�w�#��Դ�!P�1��UUI=���S�H,�9i({y<���?8��^��*N�G�Q3������
U�][����ó-����q�"vl���7)��Mz�/ۗ�~4�Mf��Rx_��>����Pm��H]�##��ȯ!� �����o�IM�|'1�OL8����?/��5���j�~F���FC�ug�^�F2��u$�(�iE��h��7U�FM%tϱ?k��SH�/�o�	��Z��5Ƨ�Ox��3aF� T��aǭi||�c� �M|$�0�͏r�f�$�����k����ۡ���r'� ��U�����D��1� Mm�9���_C-�40�]�ޭ��l^�U�����C� \��
k}���No��rO�)��[��}9��E���H�W�� �C���U��dЯH[����H#��A�E>��It��ʪg�mC?��@� �� ���_���� �/��+�_�~�n'��_����z��ՏƼ?�a� ���ד׸C��~5Ü�� ۫�4����֗�mx�H~4��R�G�E&� 6��-P~T�{RqK@	��ԴP�E��@�4i�����`�n����Tu��o<�D�wׂ(�f� ��� ЄZUݮ�.�PZ��əw���Ny������~�`�%�xv�RM_T�E���S�6X�����t�F?i	���l�(�!�F��r+�?n+�� dOI?�4��"��I�T��Fs�zz�}�=Ϋ�$��?"m�k{Kx[�)#�S��L�'��2jj���
w�M�~T ~T�w�G�@�~T~T� (�y��{P�o��M'���� ��&~�n��!~o���h�����Ѥ�ڎ=���� =��|�����K� �ך1�����V�`V�I�s $��n��}c� �k��=)
q��� �h� ��� ��� �h� ��� �3>�g���Wc�H�{��a�>����{�1�����]��{>n����KR8��O�sᕿ��ڟළn���M��m}����6��T?�`�k�/�_��|7����<b-*;H#�{�ʂҾ�m�<�������� ?i��^.���/��J،��~`�s�ic�W��9�s��5�X��'���y�xҦ�t����9<u��!���JX��_[on{+�߁���j���1�m~�� ��K����	.4]~"�6���U y�pq^���n?���
g��#��d�W���?�Ϳ��:��{yg7�~-�~�.�U�!Wixݜ�wϥx�ǋ#�	5�� ��$�����\�V�Q��s?g}�m~W��no;j|`�v/���S_��� *{��� �!L�� C�����,QE��y� �#���� �N���xc�A-��� �5��y� �#���� �N���x_�AL?�_�_7���;q=c���������� ��x�� ��Tc�Y>+�!� R�J��?�� ����a�߅/�_¼S�8��8����&�΀ h�(����ii8�� ?:ZN(�>Ԟ�qG� �G6��D��G����Ã�I�L����Hc���,;�2z�(�5�'���kG�n�`u-i��D%�v��?
�� �?�z��'����<I&��is���2�v���z���Q��O���/ٗ�ڝ�1,q_�e��"��G=y��+�A��Ɵ|E�ꟳ� �<��DMV��{A�|����8kݡ�ƺ����_�a(��� ��e��֖���$�>��=���T�[���V0E��֟_`y�N����ǽ ��qL�=h� �-7p�4n���7RqI@��2}h�֛�z��G�i(�n��Ғ� (��p���`{R���P��jmǥ;�( =����4���� �-i���gkH^}GV�P?怒q�u�SK/��x
W�9������h8ӼGu�����q>�?�}�� �^��G���'�/����%�(Y-�g��|tU �k�>��|�.�����H��x�� g���%cH�t�Z�՜Q�(Ɯ��RM��{i����hJ�潒�~N�]/P���K�ɡm�7/���:���� ��o�/�u�� ����b����� ��iڇ�u��k��>g�\��=x ������'Ǚo�$��FC�'�_�I0"�if437J��m4�i�f��R�ڑ�s}ؽ�O�)��[��9��_��?����o��U�'�OEP����H��� _� �;�����?��� ���=���H��� _� �;����_�?��� ���d��N�OC�?e�Ǎuc� NM���!� R�J����_�������� R�C\����E�� ���~4��G�BqG�G�G�@4sG�G�@4sG4�� '4sG4~4 sG4~4���s�K�G4� �*��k%�q�~t��l���*�n�^����a�����"�>��G�r���f��XY��ö�ƒZM�*�D(Xv#�+�lo�>�_��-L�����Q��TM:��e�����B��3�Ts~�_�� ��W�-�Du�R{���4�2���^m�J~�_~�Ͼ'�-��G��$����a��;�h�i5��������-�&�Y菀���u��*�
���8�i��f����y"��i���/<Rs�K�I@�jJ\0h*9��? 9�ӿ6�s�?*J)x����p� ��-'�@�G�KI�P�6��6��6��6�z� ��7\r�h�:��G����z�5����G�w��8�ҿ���:�O��ල���i:��[H��6߲���)�]��l���
����B�][+���c�?U�ejP�H�:����� PH����)S|O������{ׁ|5��>)�-��z���0��,�#\�08�
�v�zb�:���1qX����ԶkKkѭ}O^�hG�u6�C������a�/��(�o.��M'K��h}Q���� ?w�נ���~8[o�$��t8��"~=I�|��k�?��.j:�uw�.m�d�Ӣ�[T#��8A��澶�� �� ��I����� ���Y,��Ud�R�����Iz:ʫ�d|X�v/���S[��� *s}��!Mo��C����(��(�������?� �� �w����[���C��|@� �~� � I޿��*O��5�y/�?S���� �g��q��oֽ��������r�G�x�QQ��ϐ� wfq^��*:W��K�%�/���1ԜQ�4q^I�%��P�Q�P���Q� Q�Q� R�RqG gޏ⣊J _�QM%�2Bڂ����!}O� _/�Qͧ˪I�,�!p�wN }����oo���� ��H��j����|�fd6�g���5������^'?����	HU�)4K^�� >r>�W���y|��-�U�z_�D�\m)d�8PV�� ך�ҿ�W¯�� |M��j>'�]��	j���!��8c��p�^��!U��%k��a)��\��"�����cfz��O�Y����6��+�4��S�
)ߍ�4 ���3�N���@	�K�i��4 �N�i� ��~t�$HS|����c��������(}��Q}���~!� ��l�� ���@�L���$sG#z#R� ~4g��Q�Q�Pgڌ�RS�
 8�����@	�5C\�Ѹ��B�{��j��'�s�>3��[GZ�r�RE��ſ�Vm��j7^kkkx�Y�@�?:����B�=-_�?����D�$�E���b\p����>�}k�?h�=/���.���Qq�׶ҥ�Pʷ��#+����}k쏄GE��^4���K*�a�m�I@�;1�b�1�c�t�~�5��k�������:p��5~�? ?i� ��W���1s�����S0��Vpo���Ne d}�q��z����$��O��m� ��_`~�����|F�_�����x���<�n^,/����w���6��[�@a� /�c��M����F9�b4����ͧ�dU�n����վ�?��?����o��T��b� �I��5����<��Q@�'ǟ�"?�_�� �w��sD����̟��J���:l��>W�8����#PLI�r{���5h�tȔ�5��L����~߹ۉ�}Q�WF:�8��,����U���מ��>���iZT#bi�}�׾GΣ��5����ڴ�wgT#�h�Oʹ�ƒ�(:8�4~?�� ���h��������Siv��ޓ��mZ J��H����#F�b���3�
�*��3��,�c�l=2i7ep>��������υ�����3%̑6�Nіb$ו�׿	�xc�Y񞥢|:д]N+Pa����mɕrT������̶��;��q��o�Z��e�u�E�ҁ��� ����� h_��;��ҼS�T�t�V��.
�u �v�����{H�R�[��s�S�k�p6l_M�bw3B��y'֤�QUB�ڊ0��)s־����Ѽ�@�����o�P�*mP�
m/�% z����������� Y��^ds%��v�:� ��o젗3��7��g�� �W�߱w��|m�Li��$��#16�'���л��o����7ډĄ|ӯ�W���'BQm+.��{�W�(��K��������e<ȗ�P?뼿�r���<	� ?�����#~˾�ڇ�8� 
�}�o�{:l|��t|3�'�_��z��� ��_�F�R\�l����ı�8���P��@��o_��������@��i��c�E��0�A<`J�8(��}�S)O�'wvy��0ϵ%;?_ʛ^��/�IN�I�@	ϭ;�)0})���|��G�w�֙���f�����7��8��!���}⸒���=��,U�]J�#�X^� ��I�cm�#÷x���m��#�y�P�8げ>��� X������Y�m_	M��K��x������OĿ
�����6�v�t��6���>�;Oc�GJ���r�N	iYEKF�-����J����J��o�i�?�ë�i�bx/���y�-X����e�� t��c�h�$��3� Mm�9�反?|{�.q��� D:p��/iyg"�m.A�D��-�L�ھ�����&�wĶ����Wu:8J�����ܺ���*S���n|Z� v/x��
k}���J�v/���R7�o��U�=Q@h��_��|rMK�>�{OC z�W��BΣ�y;�>��� ���Q������۽���)�ћ������|u�y��ԗ�;�TU�#�_C|�����X�Vy��@�xX�g�d�n����{j��wSN���8�,�sCL�R��{�z�}|v������I�����d� u� *`;�hϰ�噕V9؅i�k;�~5��[�{Ok�c0�-�3:������?ʗ��W���	$�<Q(o��d��t񧇼ܾ��~Ļ���QI��9�_Ə8��>�qF=�ǵ %:�m- �)}� ���� � �]댟�	������ ���q�� A52�X��h����/9-��w��bW�֣�����w���=� &����?�bWζ���g� \�~�K�_��ȕi���(�?M��+]jV�{*M�n@�rj����_�����k��߱獾.���ſĭj��_���u&�&8��p���O?�m|5����j����t� �D�֚��X�p&?R+̞9F��u����3��Ht�g7��(��Ï��y����ńx�'�I��^.7t���Z����������?c�?��He��mC�0pH��l�-,ލyr����O�e�*j����5�9QV�Y�V�2��]���_�_�G�~~�6_<9{�K�e��a���{;��F��U-�Y � �����͚�V7s,���D�{�rw�Ū�q�MN���Iup��j�s��֔�x�O>l� �zt�V�̂A��u���.I�bq�^.a��P�ʝ9Yi۱�F�%��+��~|S���~]jh��SHQT��rA�Ҿ���
��i��O�Q�#�m�7��:��;��+1�֤���?����^�"\�����#��z�� ���t��E!� ������ 
2�� �� �+�o�MC�~��R� �~��ԣ�?i/�'�ߴ���<!/<=W�y��.d��PFߙ@���m�b��#��� �뺓R��p���G�����:�P�%9Y|��Nw�8k��e�--Ǉ���#|��Z��r�܁]�q<����Es��ܧҾ�+�V��j��d�3��8�.T;�h�M���v�?�� ��Y��։����s��+@��k7^� Y��n?�%�q���υ���� �5�Qye�x5�H���MD>�*8���<!��J��%�jk��	�h�(=�������?�^$�<������=*�kz_�� �!�@|�S�#�ץ|<����5��
�E�|�Y=���|�I c�oq_�f8J��O�Jir�.ge��� OCޣ(�'g����S�*�u��/�V��m�����v����#��a[9�C`͎��G���� �Io�� x]�Ǡ�\~�G������x7S�/ÝS�9��>"�la�0|������1����� ��I���x_>���^lק��+a�V<�rn1{�[�K�leZQ��{-ϋ_����B��u���S����
!Mo��C���c�'��(�� Tݯ�> � � ��o�+�c��� �_D��� �Hn�E�
��o�7ꎌ?����?��otM5��~2M��� �Y⥳�BܫZ'��|Q�!�/�,
� �	#H�l�ʛu�㝼O;���FX���W�Sx�Uݶ]n����Wu,zֳ�dW����U?ր>So��⮒L�M�����Y��c���zg�?��Z-��5��h�!�V���\ o���=]��c q^Һ����Y�6xI#V��dɢ�7K<���C���=� p�%�����t�ڍ�G%�ռJ�S�����dT��TUr�:�޽/�寄~�������*Gck��#+��y�슥4�1��������3�)x� ~T~Tq�(��P�RR��(��P�\��Vt���	z*���
ݲF�_����S��I���^#៎�c�O_��m���xbݤ[51 U� �*2x�k��hO�����	�^󴏥L�i�kr������/�K�N1�-|�i�  �>ߺZ�Mc���x{���u]C᾽)k�.0d��7W����Xb�8�cE
��ҿF�ԣ�t��D��{�=:7��)%���w��@ g��]&g�� 	/����� 常{e��K�D$˕�#�?ޮ_�	�����>.k���]�����V�{)%W00O�I�+o�H��u���I�o�ޭ��Z�ٽA,yUWR&�*��Ez��ԟ�� ���.�����8��F��_5^r��BQv�T����]J� ��Io�_�'�@����K��\}������P��'��|u��� �~3��ֺL��ml$���p0�w�^�?i� ��#������Kc�V�>�#�m?b��uc��6�2G~-��2���V�j*m�t���v�1�EFvIy�_�I�F�C�Q��y�dS&a

�d�����=��/��pO�n2����?ok�~�|>��u������3FE�H� y1
� ���M|1id4��$� j��H%�$���k�0Ju+N���k�o_����&�է���0�}+���>�O�Y����^m��/E�#�����]��ߵ&��+�:o���9�PG'����>�m�q�Go�(��?�M?���� R�J�u������~#�W�_G�����<F�)}i(��8C�zw�Sx��~4 ��fx��f�;��� BZ�=���{�O����@�>�� �������/��;����>��� ͳC��ֶ�� nN9%�ҿA?m��6� �j��>��{-6	5��"��U�:'�D?��éSF�L�,��1�[E��b��f��f�G���־Y���5
|�^���VVm���p��ߓ�G�U�ke�Kn�m�Q:���cn�j��� ?�Iτ���� C�������"����Z��6����B�K�_��-�!c�C�;�=8���:�� �%���PG� |�0��6i�P�+��ڔw��~��P�bڽ���ž�_��?��o��C��[��� \��
F���?ʾ��	袊 �՟�k�o��V���h�Mv�G��&eK��?:��q����|C�GJ��Ɵ�s��3�6��&k;�]$pGP6\|��z��*r��p�tmE���� nxg'�+7��5�xn�º���=�{9<���H���\x��>�~,����� ��G�o��9A�����9�2����K�|���������-�G��`L~�3j¦��+6���޾�� ���#u� �i�T� �F�9K� S�F� �i�W� P� ��>�W�� �d|�'�_�}�/�g��]����ۿ��ӿ�� d�&�c� �� ���#�3��� ���S��Ç2>`��יg�:����t��s��o�N�L>&?�ih�i�=u�� d��&�?�a� U��#~�7��� ��]��o����~zT��Ç:=o4���'�)~ե� �b��2� ���H� ����� ��� ���H� ����� ����^�̏M�V�� A�Ώ�i_����̿�=��� �G��� �h?��?�=��� �G��� �h?��_S��Ç2=7�ZW�-� :>ե�b��2� ���G� ��'��� ��� ���G� ��'��� ����_��9��mҿ�1oW4{�(� 6�n�co��y7�'�G�	�m� Mo���1� G�A� qh?��>�T9��>	�Ҧ���d�#��,M�a��I���� �⾹��>/^|k�OԾx^�������ѧ�坲��89��^F�d������N�r�/���}Co���?>�~]/���}'_ޠM�^9l�C����ڴ�
�I(�jK����b��}�)��].��(Ŵ�
�ǥUN7c�U��b�W�(�a���Z��4���j�N�������87v��cϫS�J��|���?�P����95�U�ξrd����>q���j?�2W]M`�&�ď�o?������¾:���-n�����݃:�}�9^ ��t�m�c@�5�}C�è[��0��"@���?����׆� �Z�o�k�d���������:^�'¿2\jG:L?4m�����Ҿ'jhU����H�����gͱ���q"�¼�Y��h����o�kٓ�O��=q�m[Oӣp@'q���_tI��������� � 
���
�k}k��,�\����\�Cazq^fI��cQ*ֵ��.�h/t�bO���4�4��gE�4#I�{��f-� >��I��4l#���]΋���}�� �l�|w�l]��� 
���洔� �����5�XJq���#�_�.���l�m���&�ma9R=���� �/��8x7M񇄧���ڄ��[����!��򯙯B�����q��~���?�I����������J�+��żd�%�0ϱ�sg)�?Xי���/'�(|G�J����|W!��I<�P���s3k��Y�Ґ���]_�e�;�~�ZƳ�ڵ��֐$��)VE	����!��c6�v�}k����iBr��OqN��&����#ƿ�'k�	\[G��]�(��wy�d��p���k?��U65��o'�=0_S�ƿ�G�O�:n��h7Z��Z��ML�d`�@�_1~�^%���w��V�i}5�V��J���?:�0�J5��0�߹��J4Ժ�mƹ�8Zo:f��=k߼�|H����Z5բ��ݲ������#5�n�hC�z���ӟ�?���3���=����l���ⷸH�Yt��^e����Ҿ������g�^<�������3V�0x�G��q'"2�+��Lj�H�!޺�����(����b�.������Ўƹc޽��<��� 3��G'n�S�:M��g��u蘆�/�I�c�Ө�CXR�:0ܨ��ց5CX���l���[�$�=�4�п����iO��0��{�S���k�Zk0��POO��ʾ��m��.�9���$���Q��b��G�K%A0�3���X=k�ڟ�?� j�S�*��5�@�K�?�5+-[R1��0*�0Kϥx֕�#xWE�O�?گ��BHs$vz�Ƈ��)5�����ƭ:��U��n��F�����
꛴�������J���ޱ��}o{�]F��G��4�E�!�c�3�ԓ^9���[� �&~���E�����6k͵���N�27�%��P�.��u{���� ��Mw� �w���؛�<+�]'Ǿ#��c7��X�T.�����v`r��T!�&۔��ݻtIl)�����7݋��'�����?ʗv䈞�5S� R7����_fyd�S�Ѷ�+��)���U��X���������"�Ǐ����9���ֺ�Ǌ<U5Ε��N��md�_ܪ.cBA�cp,�������W�d� �:-����¿���bS.�o#�s�c�I$���NH��q��+��Z�[�-��Sˌ�q�;�/ۮ: �f�a�i/�''�����5���?�]��>� C����Y
��h��21�� �ҿ |C�j��N��Y� g��A�6���ʼ��K'���pA��>8�wfgR���?�.?�3G��?����r.��	��q�� ���ۏ�����F� ��B���hO����TP�o�����~�q����.h�%�u�������o΢�h_�\y�:>�q����.h�%�u����}�����9�� ���� x�f���Y����sG�@=���)ۨ\���4_x3V1��i��7W8D$����H`�)4��Ɲ�����'�V��M�]�|u�����6%l�[YA m�۰�� ��J�?do�[����!��mH��tʨ=����xCGv��y�`G���� ����?¼(�q����:�X^��� �����|� ����UQԿb�x��mk���k�y?�T�+�� ��N+�� �Cto[����'�!�7����?pX���i^�u�-���7ᯆ?c�⮻�ό>�֘��i�j�$���$Ip ��}2Gk�#xd�L�yru�15Vi6�	Qg���w��ZL��,rq���a�JR���0�5-Ћ��g�������
��ο4� M�{�vM&y�[�$P�y�\�z�~�WץH��S�=+���&<��Bn��~=|]O�� �O�Q鍢��	l4�Hf@�$��5���Y ' �5#6�,yjN��� ��B;"e''s�/ٿ�
�~�?
l�?�o��,�^�uwUVf���Ҽ7������v���iRhiq�X�Aa�y����F�)��i�Ř�嫚��:���4u��ݨ��xK1��o�?�� N�U��¾�����5��dr Y�pddf�+��5"�J�@l�U��S�EF��
�GM���i� 7�w��p��`_\�ٱ=a�85���3��/Vs�)I�O'9�X���#�������x��-WA���X� x�)����� U�Q�ҺZ!/�KS��l:� h[�tj��F������ hOڋ�>;x��Zw����T�ҮV��i�Y��U��X��0�V�_��<�%�;��k������q��FH���W�,Ҥ#�8(�7c�8x�D�|=��c������ڶ����׼����3�ڗ��� b/Y�ZjＹ������4y z��o���e/��feU� �Z��p�+��UʵH�B	�'q:��g�QJ�1y�H�E�i�3���Y��b��u��� ��𿁾9xV?xn�¶���!��Ӵ�u���3�Q@����j�s�+��V��5;X�Gb�h�g���++�^�S?�л��� Ʈg�S�O1����������.�E��Ǎ3�s;c�櫉�-,#��m�cl��`� L�?�+�Wֿl/�a��'��b��jѠ�7�a�#F�~e�x���_���_�oNѭ>xn�;(DB�T�຺�դ�Жby���q�i��	���T)Jj�g�����Q�&V�
�橜VV8?ʿm�2~���/xRM xGN���s,�������M��O�y�V��~9�\�Q�|���|8�C�&����_��Ⱦ�t����A���k�	�C.KY�Ԣஎi�i��{�6��{�6��z���� �9�~��ɞѼ�8�>�t#�O]"	ȏ��|�\��؟�{ �_%� �7����~��w��y��omb<�[�u��W�2��IZDd,FG�Tg ��|�W�Uժ�y��]��E~D�Y�M?I���ii7���ݯ+N�$����B�2{(���I$lʆB!A �a��D��n>!j���ƫ�H����A� ��qsm;&�����<�*�w���k�-��w�Ϋ�Y����i*N��Թ��<�����sFh?*?*\њ Oʏʗ4f���������sFh?*?*\њ Oʏʗ4f��m.h��i8��f�����@�q�K�FE '�q�K�FE 7�_ƌ��*\�?* ?M���@ǽ����*\�q�I��O�&�@�G4���+�a���h�6�1�����O<�o�*?�����~���-e�F���2C�Eb����l�k�jRW4��+�g�ê�o�t|@�h/���3m`N�a��}���(�����m����kHa���<���/����O�P״����[����o��;��dج��+8#a_�a\~��]����T7�v���_/����pС���Wd�T�B�Yѩ���B�Q���x��{�ׅ4����]��$�����*�n��"�9�Zh��P�yAs�>���+�?oO}�+�٣���#-�r�=06�ք�Q;{�i����!ve�,�6w�9\���u�C,��|=9r���#:�U��&�;/�*�u���3(a���������_�*>��_�7�~&����W���Ks�F�~����q�~�� e�@��ϐH?�ׇg�½L�<�t���y�Y�!)��]2���HY�Ё�K��1�ݦ��i����Y��� ��_��1�+xv� G�Q��j���/q����x��_]����� ���߇|�X�i~�� j���:���-����<����U��~���W縥j�W=�;�W=��W�)�Y[��&�PB��z�ş�ox�#�'�U`O���_�y>��� Q��>��OH��V���og9��̏qm+���h�����3�7��@ϥm�Ǜv&��Y�����7C� |U��� g��4h��?�����y7?��PK
     �8�Z�|��b� b� /   images/ed998360-ed4f-472d-a3e6-52adfa722a6d.png�PNG

   IHDR  y  �   4�2   	pHYs  t  t�fx   �eXIfII*    	      R	               (              2    z       �       �   i�    �       2020:08:13 11:56:58 t     t       �    0221�      �    0100�       �    R	  �          X7  ��IDATx��}�&Uy�)��r���]`)RP�HU)DDR\@�F�KbLb�5�$� (*&�h��ш�X����E����}ߩ�|O��;�!��=��2�gΜ�93����<�ǳ�
��
O8888888888888lo8��������������Ḗ���������������Z��k988888888888l8��������������Ḗ���������������Z��k988888888888l8��������������Ḗ���������������Z��k988888888888l8��������������Ḗ���������������Z� �Z)�#Y��֚���y�,	������b��Z����f:��8CX0����e�������e�)l��j��g��y ������ô�j��<�SaqN�[�8���(�i��9Q�Ci���Y��O���h�e\RLe>ÍEł�b��O�?L��=�����0ʋw,|��S,��0X��Ǌ4q?�g܌y ���_���-���lJV$ʖ4����Y�����O阖������ãǵ��Gm(�̚8�o���o}�[=�вe�`:@-�` �f̠ �C��C^����(I
"I�&i�&�0�"M`.�}�嫿�'��6�JbW��B���TH��1�r=x@jܫ������u������1�u|Æ�:�9�y�>��뮻���|l�TK:���������(�q-���!�4<?ܸq�5k��%K� � ��n��,��xB&$�	�+�B̑�+�!vy1�a���]C�cx Lr�,��� x+ �ܘ�Qǘ�9�ZB�ɿ�wT:�*�_��1�~rr���@�8�����~�����زe���8,����x�H]ࠃ�����ãǵ1�T�<�ͽw�g��"�J^+LQ<e��BIA�����(�2V�!�%��y�#>S9��!��Qv��
��8�x�~�g��3"`J��R�P0+mbr�����F�4Kʤ/���D��� Gp.��
���P���/E:�~<�j�������p\z(<�eP(�O����Q��u��u���>h������&r���8���(�N�B���o���걱��`���'''{�^폪�W�G*��1+b��E�Ӊ�T�R�k���y��$I�;�aA�fX��.����z�
�s��RE�0<Ξ�����Y9��@c�-�c�~[� +
vd�3���� �Pc�у�k��OG}4;�|]>��rppppppx�Ḗ��"�,bP��� V�e||��<��t�o ��5$�55���yS��4&9mX't�X��V�,I�>&�M�Ih	l~�&`�m�݆f@r�+P>h���AK��0d�T�Ș�XGhƴ�F8rc=��^&e����I]�hI[L!�1�L�yo�f9����`���^��|\�`H�G�k98,J��¶7�tИ������� �~�:S���f�gR�'l�r��N�Z�vmS��;dNž,X�_��n��,"p�'e�`4 �c�f���=�ԬiZ(X��X�]�A:�q�HQ�nh�Z ʒ�T�Sjdd�ޯ��u�֝v�iK�,����98888888<�p\��a`�h7�ˋ�Vg�3d��DE�b\_a[jH�O(�PNhe��Z��*��1ݘ�xG��j� GH�X��2"*�ԙ0��(����,�g|r2�A���@ �j�;��C�[�-��5�ƨ���?���������R{0Ì2�K@ �85(_G4��284]HtRi���9{�
�)�ae�"����e^��	�۴a#�a��é��q�a-�(]4=�J888�p\��aQ��P��˗|��?���,Y����
T���k&D������Jkv�u�$I`������ �_����Yꝕ	��M�6AX��@{����� O����7�m�O��[�O	���4Tt����Bc�B�����%�;�h��n�:�V��S�0ݫ6D�H���XVW�1�Je~Æw�y�o�[8�M4"0k8���������h�q-�E�f�aι�]�������̤H�
�b▶
�í��;���5V2�@�)<��:(2��<K�<-�Aڛ�'���I�Hc-�
m<U�.J\Ll��{�e˖	L!K7o�+�MYh�`T06X@�-�I�|t��{q<,鎢�	
�NG�	����<���,��
ʶR%-)r��`�z�ra̡��A?��ȅ�O��lڜ춲����ﳸ�����#���2sz�������ถ���@��o�Ng����m���4ݸq#|ð��hV(F�U��(8���l���+����27�_��p�W(F!u�r�X��jxxx||�wlj��������0�6�YH�tz��rR�C��Dr���*Ma%��tY�5�*V�8U*.J8���x�6��lذaӦM@��V�|-v��g�9�v4�[9888<�p\��a`. ��W�i��:�ȣ:���~{����F�%��iO0��RLi�uX)�&h�OMM)�QaMgd�p��*�ǤkƖ.]�reE�/�~���	`A��Z��^{�Z�qÃ>����'�=��F�6@���#CCC���3����R�lQh!|�(p���q?N'��y�w"W4(TYC��h��@�p�D*_����Á�+!X{�.˗)�]�I��YZ;fx���S���\�b[}J�^\����{)G%�z�
�~f�=�5�rpXdh���~�Lf��կ{��� 5���f8�4ج���Ӵ���7n�X���q�n�;],F\U��m�7��t��sϵkײ� t�u�V�]˗/�c�=�5���q�-����q�)dx,�ݧ������`v�M1��bb	�SV�B�E<%o���e1-J�kg>����GI�s�1*��Z;.
x���pO'�Eǵ�����d6��@��g��=�n���GM
��[Uf��Z�?�	�(���[H��Egd��
BXȭ	;��X'��L�22V[�	�*789���׉�`ӦM������t䭷�z�����n@��l�`�VS���Q$ގ�O�T�(+�Sр�i�?3��0z��F� �{8�ɠ���6Jd�4����6�߰����4�#�N4�֢��������&}�z��rpX�p\��a`�_�2��|8En��{��?��?�1���b����)���#?'n¢XZ�b-A�%�7`'ʾ�'�*=������@�V�Xq�!�LNN�j��CCC��U�bq�
	b�>�X��#�(����/�0�V�7� ��)�?��[�xT��e��0c()\d�����b����ǵlE*�X#��Y�	���+��)IW�/"�A���ަr�KJ�P.4D'M���qe�H*��	�1I��	24k��0��=������]w_y��o������������=�@��ޔ�1L1j�9��-k|�"���qQ0k���"����l`VyJ��Pj�+���C����ȭ����g�E��Iz���xdV4�M
���=�����r����H��󟐿0�||î��{~�s�"�K�h�İUK6�j��o"s�VNB�L��#"&�J�l@�#�Pz ԼPX3@�,+2�����,2ߡ$�aAn�����g�(��0X]@�Q@RU�H`/��Л���WÚ��t�z٨P"�s�8�c��P�E�,^�LỊ��
�_c� �!R�)is���X�@X��&|�G�tR�"��U��$�7����
���8M��p�ȼ���Kh+�\O��5}�M
w��h�H;���.<�z	^L_e�ݪ}�.=�����c��60g�k��3�F������Y `���xh���a�ĔY�D���/��_p�v,ڞ�N�g��0J�B�p�簈�:�%{Q��
�撱	9�1#5Idh>>|��J��t98,8���80��*�%[?
����;|��I��	Uլ��"Z�"��p�.L�B���ܖ����y��s�*`�!5 n�K�,�ϡ���z跿��{�q�G�r�-���E(�|�.��i)���Z�@Ӝ�U礉��"Z�Ue��\yYP\"m%y� J�~?kS3�S��h�T�$��p&����7̑��x�s�+�i�_*r:-�ޠ�nI�7�
���jg6m@@4���2���$g�.� b$��a��J��тM����r�L����$0l=t��W��XL��x����8"'�(�"��7���*�X��$y�
+���L�;���"j$Ȝŝ���V�����â��9v�=<�H�(pHAMn5�/�+��f
A%�S�e��(�����c�3=0���SW^�����1��2�'�^����Up����g�����|��0A��nG�U�c6����o~�����Y�f��'�����L�p�;��myaD�%a��?<O�>[��)�Ew�B^�t���o���w��C�������N����)dA<��Ϻ���a�� fio8���Xถ�âS���*��mܔ� �X7�җf2f�Ŕ��q�D�܌�NӟV3&Hl�}�Df�X�^�W/�������,�e�7�������yZ$�e`�Uk�U�B�Av���(|��+��QW�X-�X\����$ˤӷ�|�<Z)m��j�	m� ˁ1�a]�}��p���
��b
H��aǛ���>�<�y��`�z>���5�@�t��Ԥ�v���pAR��-ˀ�ŉ�w�P�D�C���3��E�c����-#���ɱZ5� |' ��jeD������� �Rz�A�-�o����6������L��=�r�]���X���L�d/� h	?)�{�'����d���[4�:�h���Fߙ���oaҡ[U ����p(0n���^+H|/ �����5>[�a>�|P�{:Ǫ��%�Q�u�����o���g}���V2�x�<+���5#Q5�⫝̸vG���C-|D��?��G/Ma&x-�PSYă�{�������R��ǽA�*OY�2>>՝}[�������H�;�`��>ve��(<��8�"t�Q�-=�����"�{�;8,V 7H�$j�K���t�ͷ�vۊ�+���`0��k��`��(3JjŴ����{�R�V�����d��qIbh����gÆ�n�#Y�~=p-V���\u�o['��rJ�:�&I�mYr9vU�Ծ,��=�]v�!��H2Q�O��$����0t�q��ѥK�0�]x-�=���!l�h��h������x��O�s�e�����Y�<��|�#6Dl�N��� ����u�x�;~�5�v�&����7���/yɋ��)�I���[��w���W��
8�Za2^?M/���7_��ݾ���W����^U�m�UO��t�_��o}��Χ�<�|M���/P�x�߼�k�������w�-���DZ���^y�g�����8��C����F֛�r�7>�s��c{իΆ�0��dѠ&A��;�y�^0�#��rt�`e`�������:隫���?��N8�9������É��˟��������Oطr�ZQ���>�0��C��������?��*�*��������������}�-�u�~*�8������9�Bd��)U~�1����f?��?�O��������C	���{?:������t�I�s(?��(���z�K_�d��AO�^Z��)��B�}�{��o����<I
��4�l��*�@�@i"�[1K`V!�rpXp\��a��8΃ �'����0|��
�����!�p�0���������R�z�>X�!Ԕ@u�4�b��U{��$+�d{��diӦMe�a	|�������1��;���$Y�{iwI�]��6��[���N��C�eZ��C`*�� �
�F�G`�����t�1c4�{�X|�e����Q���E��|��,B��!8u��^�	Y���|�+ߺ�+����>�HOa��Vٟ\���p��Du�~.��n��Y�|�g�tʧ���V���_��3���/���z�k�J��m�n��W}F����x����ҥب�$[���{`��r\�htI�Z��e2�<[3+d!|�
t�f�`�&kyb����aF�41p�������o~�3�.0�,�")���;�ǂ���Jʽ�i��	��	�m8T%zB�,O��tBL5���8������z^���XEA<�i|�����W���_��׎{��0�Zu��@���Rf�Ga�`��x{�H���e��U�E-?Ic�`��³E�a��p��y�{/z�k����G�jx�:]�s��>f���#��Z����F�?���������G�_u��.L/��1O?��.��k^s�wo����8�a��Xa8=�meu��F^�+�(�D�Gn��.�i�$1�FK��Z�����~Q�-��e�
��>ܣ��a��Y���� r�~���` ���U^��ze�)k��D9�a����yV��Z-L��b��֐`O�z����Ӓ%K`v��^{m޼���@���	����-�JU�Z�/���7�I�"�nu*�i�������8:��tb�%87đ,����F���[��|pa寣K-�|>b'@�qW�B��\~�+_��(��@
`H�xÛW���Ї>t�3�87�%oxÕW�۾���ַ���3.hu���_s�5o}������3�<�_�*�+V�U^�f�D?i�P�2K�{n����n:����N�"��RQF����~;���vpb��4���k/:&�YbZP�,�*{D��^v�e�s�A�L`B\����Yg�u�7~��7����H1
U�md5%�	Ҩ����@�\���u��^p��R)�^��&,gy&�=[�\q�g��L�W|Fz��w���ėN?��_��cll��H�}���px4����8�C��(H�ַ����PP�zQŔ�'�c�aAN{~$��iy�2�4<��X��"���Oա�0���a���i�z��.X��+ƹ�_���I���[c|�V|�ԭs��yx��<����Fxf�YO�aT�f�������I��9��rpX�`�c=/�"�Do�ou��055��W���E%kB��PkέcW��ڱ��9���s�$)�MPP�1hV�e˖��vvH�6�
c �U{llH�������ۃ1�Z�Q-Q�$`qF
��T��|/(+fa��R�BR�W�EL��m��Ї�j�a�ƸG@!2�ʈ�v�X9�/�I�yE�3oI�[�#%u�7�@�#o���o�w��x�X�5k�~�s�Y�ߡ���O��$�̥�z�3~��S�?���_��O���~q�=��ӟ��}�ǿ��q��9:?�����U���������}[�<�2֦?��/}H̾�����#�cRm�e,�fL/ �>�ə���%���f�<��Z�=���}�S'�����@���p�gL}A���V�uE��n��"��<	�e��
�AnS�Y(��%Pt�-NZ��i�Y6}O��7�O�Ԡ�0h66:r�e�l��O~��������:�����i�e�;J��4�K���_4���L�%9T!��U"5I!�J�Yu�'y������om�g�P�b���^�D��e6�7�c��`�kea"����W��z�E��Q��3�dm�� �Ћ�GK����E�g������Ã���MJ�T���r�rQ��s������p����b
Iw�|�J\�58���hд�9�/�D�|���~��_�Kahhh�ҥ�n����������|���*0#���Ac���^#C�E˒t�y\̸2Jo`K����A8�4�O&Z�D�kC�6�����5 `Y�i]��B{�tp�p���b����u��%�F�S�rd9���.�������]X���_N"��T��&v2pzL �-`�BDx��T<�O��ӷdY�>���5���K�hy�9$R��zIv�Wv��_��.>�S/{��>�ϟ^�f�1��S�׿�u�%���gONN~��߻��[8� ���1w�}��Ǿxl���S<$J&�'ԗ��o�oYf��/���0&�`膾�Z����I�RgJ���"�sR9h�I�g����H�B�I���z�UaW�#<+����\�L�@����,����UW]u뭷�pr���6)�g�a��p��&�ՙ�u����3\5��x�i's�1"'_e�G�~��_~�9>��iC�`Kݡ������v<����]|����ߟ{�g�}�Uy���S�r(0"Cw�O�׫^����#m�^C�~E7|��Ozғx���tLm�}e%U ���~0Cʙe�j�����Pn^98,8���0K�N|�S�7�v+��yht��g��ɯU;X����������$-̛�`&B�9�I���<�Y$��Q�U�D;X����0�J� غuk-��^�J2��5�B��(lg�z���� @qB�Tu{Ƴ�.�����������S�ll-��ljr��7X9����kE��n5Yw����2!
����Z�[�����iݪ��R^���������GOZ�֠n?F0�t�|�{?������^<	l��Z�aq���(+�:MN���ڟ|��#+v}Ƴ����C�~��/:���؟��7�ݟ��{��ĳ�6^.[��KU�WV{2�lR�?Bc�/�g�u0Y0+�Pm�3_��[�w�VC���5=�N��c m��U-��KK����(�	���2�V�e��(D��-l�ږ0�P��xXvL��	'��{"}��O\��7M�K�g8����m$)�ԡ�FW��j�T�T�\Q��*��x?�QlO)�� I>��O���Ru|��TȲBaQ�� �
�8�GL��>z�=����w���^{�%�=��[���uڟy�S���|�߽�o�Z�BNe268��>W�ce ��y�P�2��� ��!ߘ�z
�
� ����Tr�	�Eǵf���� .q�m�m޼Y��9��?����.�K	T+�O��"g~�n�dZ�/-r�Zh��R3PT�LK؅Uڦ�wbB�^&ۨ8�9cu
����G�;`S�q��nioxx8tQdh�2�3���3YN��P͐��������>�̘"RҀ�y�b�ԋc/&�M4��������g�'?��_��w���t"���[�:�X�>e�V%��9x���Z�ꦛn�c�}�9�'\s�5�y�_��'?��ƍ�8��p�}�}�S�z���$�y��_����'���^�����\t�^I���
���{'>�X�/�x��_����E�ǚXY�V�z�)g<��Ob�p��	]}���:�TA��\��X��(^s�E�\rI��a�Չ��Zߺ��w�q����
uJ��s~�kt��_�w�V�bWdX6�eX&k��Jw���@SJ�_��������^(�>|=댳���o|�o<�����qzG���9���t)?Ks�X��1� �K���\���k׮E����S���`���o�g���rQD�>��ϟz꩞�A����A�����.� ��=��>���a���Z� i��-q��7}�k_r��{��p��̬9�(ٚ��q���S��ؕ��X7�c�!�bB&Qu a���
Pd�����Mj�
^ �K6ٓ"�8�8�~��p�6mڤx���D��+���4���N+� �''���,[:15�T�u����QXϪee�:�����<�t�Y�ל������`M�Z�D��.o}���db���*O1$|��`�i��V�Gb��y~���TwE���g����\�l��3_��?��Ί'������v�ԧ>���V�X�������AA��c���2��'-����u�L��,����A����i�)�����V��袋��u�V&�ڒS�R���A,�6���ʋ@�lˊ�`���"���®�4Nt�.��'�7O��T$�/z�V!����G���͠q�	:�H=_+��Fǉ�2Ȥ5C#�\�֣���R�3{"��8��8���������K�x���//z�KB�m��<�ZE�V��Ak^�u,�X*KѤ���ܢ75@����`��W��������<�y�|�˟}��ސ%�x�u��=_���MMx�K��Vȸ`���v'`rrv�'g�%��/���a1b�2,v���?�̥&;��ҥK��A�%D@(K�RBc#,sT9��)'7��+ ׮�@��'*�fG��.�n�D�^3�̰��&9�{���x�<iE�S^>����������@Dn��!eE���zX�̐�E6��wL�$�p|��	l����+�����BǪ�:��nz��^/n�#�!��^P��m� w�y�>��/����o6\w�u�vԷ���Vz�A�|�K^���~��{��կ~u���r���:��.����B =�J��h&��)+L�]�qb>��O���V�>t���f�tO?��K.�H��idU��Y�������0����8&���G?
�2'�g�}��`��P�2�9C�1��ǀ�[��������w�o��6{��T��p�C��&�����2
����Ȋ���G�x��^��g�t���c��i9�����y[@��d�i?�r�n�v�������5=��#O8�o�qӦMccc��L=�,�N�۟`<�IR���Y���F��$�.vD8���`U����[�mEw�掉��K��lݺy���bꢴ��ޤz\��/}���Fi(�G"㪪f�2��DU��o�Z�L�7~����|�fk<*A��l�������d�(bY`c�ga|�~=ml�����tH�+�����{�%q����}�����������#�|�a��C=�>�C�NTGr'��H;���~䓫W��X�XJ�� Ι���Fzh�}����p��n����%zJ_����D��z����/�?�x?�H%r����rɚ����{�|h�e���R=)c��5���_�ҋ^��^�N9�Dbb����
+Z�I�Q�(�M��w�#Uad��W��Iz6kI������g\�7�ս�����8d�ލn�L�L��&����Y���>�>l�?�Ḁ�
�%�oM.N�,�Zm��<�B����#+/OM�~p��r���<iiG2�EW	�R�h�HL��N�t� 4���QJ&�Jf�U�'���=�����×��'���?���=�Ǌ�>�T�(
��9\g�riy��_����=�����E?��כn����p�+a�6/�~;
�A���Q�2X�/�v�AB�TC�<X.(9<�=T�DD~�C3�6�	/�k�p\��aq`�;@�Z��9�GHK���܈ �x��W�,��C�V�%�8���Qu0a������T�}D�BSσ�xfMܡ�j<s����C�W��� �D�B�T8*[�J7Z�����@
Θ8A�˖3�6n܈�`�+(W���� '�0��Mc�<��l�^����
��Mo��_�w�%���_2a�0������w?�Ӹ��'=������wV�2��8����'��p�W��Gz�m�]u�Up�w�uW�f#�"r]��|P ������P�ʁ4U�����Ʉ�7#n��ݟ�K���_�ӏ8����yM��4-�{f[�Vd��J�ߍ�����v�p�YV���$�T@��\��<'�Ki�� >����z��_�r Y���P��#}�Z9�cG+�.-�h�M_x�W^y�>��SO=�)��@��)\kYHʰ2T�+��,M�V�+�����z�O��3�=�ܳ�� B�s��޿n��ի9���$I�݁�ۚ�����{�~���	m�r�ʩ
:8�p\��a�`>ǋ��8OE���vR�q���1�J�YL�p졸����u�Q�e.�.`s0s��-i!�vE��EM����\!�:,�X�~QG�a�J�f����e���Mi�S�����j+s�#��e#{��Y�
��΂�d��!�l���?_�b��<66�nA}�;�����;�"�0���$��m�A���߾����g|�3_<��C�������3=Ԗ���k_�����������³l�SI������?}������~����0����`�u��^��ˮ�v�'}��{�r�s	vՖ���4�0 �X%�S�-2��V �Oy!t�y~>5������^gM�����O}�/?����k���*��T��/� u/2i��%9d����Ҟ��#�:S�o��6"m���r���gŐ��d��Z�K�-�����z׻>���Xu���~���HF(y�3�5Dh��ʈ�Qi;�=AJ����S�B!�d���H��=�Q�jվ�}�_���o}�����>w9�ϰ̓��?��s��_h����J�Y�f�.��.�����~��~�+�~��S3#��?�؋���/�^�]��@��t}��c]A�щ�P��{��0ǸV���5wv0s��k98,�iE���E��Sv"�z=`�1����b�j��u{�z��a'wȌ�+E�W!8�O6�r2�kU	Q�5z�0/��KDQ-N�?aW�E�p��$=0�+���1)�$1�(�$�4-�t�-���E�iVfyI,G+I�~dt��*���[�rQ/1]�f���;0�=((��\'�KaI+�y�(e���?�#\����3��k�{z�6�
��>����������biԓȟ��g���uϽ�s����1px�z�S���?�G�8���Y&�:�DQ^��/���\R��P��(�Y�����]vم�����0H*��ӏ?�U���_����o����+)+��0���=�B�<��&Ĩ��\��׾���}��_��7�A�DŊL+�Z�T���r�-Ccm��j}������o�iE"���n�]v�@O����t��IUi���a{a��#��&Si8
� �|
����{�;�����+�^�B��},CL.V| fIҊZF`���%�uV�;��n`P�u�����P���+�<�E/�;I��a�L%�|vڭ~ �yګ�SSSc���{.����~���#�q-�E�f<^�d(�D��?9Z�"0"��P�S\���V2�g�]|A�.$�#�U���𭜭�V���˪is-M�^< K�^L�*~�,mS��L�9o��vLA�N��	:��3K1���C�ZzE^p�E�$f�`WN=�aXcUPN��x ��v��e`$��8�o�j�{���F����|�ҳc?U��W�"�{�Ʈ��G��#�<*��G�د���]񌓟�����7��\_��9�O��gg��2A
&3��e)\�ptծ�_l����;��d��w��?:m�n{n޼���?+l	��Q�����E�+�D'F}l`;C(���4K�"�)�J�N�3��&7#p�Î~�G>��k�������N8��g�}�	�&l%~��㬈��cE!S4�[��(��I��T��Tg�O�5�)����k�Ɠٔ�Q�̣Ѓ�ߪ�8㌿x������+��$z�+�w�y�v.R���e�*l�#�-}q�lg}~�$�C��﹍�������^�}�Y><b�Z���$���H�~7�Ŏ�E���q����]}���Zo~Y�:�o7��QKܻ�7�,�k`L�<k(��h�~F98�p7���"�mj��i����n����<�I��e-ч/]�uӃ����Z���A�mQ~�2�\��@UG6KZ5}G��w�ZF��Dڪ��$�]�Y�9�܃8fv���]�{�D���d�Vr1eT˨�-R�^ ���m��9°���&`
sA�_���{,��8��4�ԇةp�'�Yd��)s�N�B�#�;��gQ�LÁ)(�	%���u��Y@yP:��>�@_��kA�C�����+u�}k��%`�f�F(e��8�$`8��ڡ�Q4{sL�3Xy�f*fu�q�ҭ=1�&-0�UIM<<cYN��i�#�6=������	'�@ӳ��x/�^B��z��Y���g���_y.To�YS�r���.̼.^#JD�_�?�¬�MNv� )�0��J�"�{�^8:�Y�V��uMg͇zZ��݄qpؑถ�âS_���ܺis���H���r@�}SnƁ+��{�ka�4����h�b=M����yM�ӆj���Y��I�ةE3�^���,i�9`%=S��h���d�EU*W�&����j��F�EI���X���FTf��lH��.��������e��MI5A�d`�Uo�������p��p��2��R���H�|��L��ϳ��T(
`;�Hn2�`;�V��1*P�-e�M����� �Q�m�yZ�N<�rۊ6��q�i�F�
|t\hU
KJ�Ub��T��0O�{W6��L��Hѳ�٬�kKnO.���y�L��ʹGL�4`HmQ̬I���Be[/Ǭ~0�:0���je'�2YxQ��<��?\e��.I�4�J��E�ݔ�a��c\;�rpXhVl�c��d�099�|�	Y|/��R�Q0���N���y�D#/�T`��&�(��tya��W�	Z���9���rv�!\3(C�p�j�BP��`�����{`��1Ųe� �H���[�SH���^/Mch	{��i�&8]I����`�B���h턵�EEw�T0�l��y��2L���$A���`w��kUJ��GGVat�E�u�Pa�
�[Uf+lN�>�TB,E�и�&|�`C��%�P�ZC�$�q���`H���TAYg�n*��=��S6����j�'$Is�����,)�`(�h>��pQͥ�i@;��1�G��U�'�i��] �WzO�o�b�*�]b��c�Ӗ�bq�D��M�;�a��Q#��8.}SV����cϛo�9B� ƫ��Q�*|��+�F0qJJ�L�J���-[�}ڙ���b�U�^W����������b����J
L�X��T�c��)Ξ�1#��B�����^�*T�^��r��)/]�ա�J�GCK�X(�zú��V�ߏ���>� ްn��1%q;!���Q��W$X�&̊��DTc1,�]I�
ry�qҋE�,��ߖ$�Z�����H��.�0ȋ�r�ƭ�[әG1	6w9gϒ{�*\�ì���+�l:��0�u�Q�����D��(�cH�G�T��T#n.�b7,��q�):��<���t�h�v��3�����@[��2�bHe��|la�˱m�����*��,V/&��U�����2�凾�~�O�������Z��b`j7�e�o��FFF�@d�?-�����8AB"=>y�r�~�R���#~u|`���z��Jo�g��/5s{4��t����,*_/�`�AFI�p-w�~9SIk���b��/��LI;5�}��Jaq&͒�`(�Y�FH��h����|��V��u�VDЛ�V�"b�_P8?!�Z����(�d��d8����(���$�W)��O�>^���B�O��ABD++2-H�Px��U��,�Dʘ�f���H�\N�uGq�|��%%a�q�S���LS��9g�����7X
�ݭ�?��a��"{(0[Mfv��Y�HΊ�aKG�vL�D���)�	�o�:"ūW�^i=x���W�wH��S���:����ag��Z��|S�� |�E�����C1���D/�r�E���C�� {�E��1N�bI���ک%�l��e�U���gF�!aئ(�c͠G�Ֆ�{�X�,�AY֠�!������T���<�j�ǎ�[��Y\��e�Q�Ê4K�� |��V;�{��4ټy#����������a���Xƴ*i*v��˪��X�p!��B
���t�N���M�2Tˈt@�0J�\�	[@�s&"\����AǘR:Ș�D���� �L�'��L��ڏRa۶O.P�X*̢,�:��L33�c�X��R]X����ڭ{�y(+a�]Szh����G��lkO-(��@��rMU���#ѐ����Su��q$��F�?Ϭ�]Ξ��C	ǵfZ����>,�E{��]��Yɚ�4�JY��O\��t@y��X1�H���T���E^�+��dMݾI��n̡�ӹ[�a�@�Z�U��$��*M�0��䙕�6'O�˪�V����l�̺�MNNNLLp��`hh� ��7�ld�`�<>]C��L��ڟIQ��#�D��Rp)V:QRK�TL��?�U(�i��0�ɛ�嘣h:W�-s��;��1�rmX� `�lt��{�k�]�Rm��vM`ADP����m�2]Q�gC��<�u��y�vD�k��E��d0)@���g��=Lu���O�Yoy����%�Eǵ�:[��t:�A���#�\�z�߾罛7o^�d���ʪY�%����C	�L\��i� �s�Y��6�2+V�����J�)��J�i�W3���}�*�vD]\�ژ������8~QF�� ���� LYj�cr)�Q�;c�����C&��6A��޴a}�yJ&Y�[��íN������⨣�b�F�L����Qj�O Sͅ���	�d�^��T�9�jL�3��_��ۑ��eJRnd,T�]�
_
p��-RY�g�7�Wy��`��=aS����ԛ_T5 Q��p� 3�FN�|`o��i{�Fsfy�4�iVT���v��O<b̵�����;_ZU϶�&L
�ic,%�������g�s�p?�w���_98�(p\��a;`!n{����hQ��#Za{����s�=�A1i�Ӣ��X]�#O�bm�$I��Y	W���˪�BfA���)*/Y� Se�!��0��ظ��.�n17k��*��A>F˪R����L��Uh�4�9!��j��<lٲ�B"��g��]9zGƣn�7%UxÈ�C��*y�%�qHEq�Eux������D�m(��S�1�G�n}䘻��������.��J�N [MT����Z�sm�G)X���R�M642$
s�a����7\r�%Si����j#/�䃊B�i�ՠߟ�e�\�b�T%�^EM���oz��e	�_���	�La(�@GfY����
Y�̍ZQ��k�O��+ֵ����M#EAAhT�Frq�Z9���*�Z�^�26�T?dE><<g v�d� ]�^{��
`%;.�^�������|rʼ�ٿ�J�.5�XS�Qk�]b�i�)f�!^��\���׍������� �tk�#i�0�9G�ȏڈ鋮h�f��o���y�ռvpHE��g[h�R
����ط�?r%.~H	ǵ��<c�s�����`�zEс����~����O��}Tņ�Z �'q��h1w�Tu�SM��уM�U�����z�L�x��^�� �Ù`�9�� fnb�ٮ�jT���d�s_�#I3� ��8��l�244t��A��]w�끉���1u�G���KV��٣)�.��A�AF��N���'�}
I7����#�C�����q-�m�����̫� ����nS�!{���⼳?�����ʨZT��������z���)��E{�r�l�kU1�i��\���������1J�vʘ��=�]������(�מ�kA�@�w̼�Fa+2d� �0Ȣ��,Xs��	xH������/7��o�����4�#�=���[��v��%Ij�[�����/��7�r��8"Ԏ�z�;�����t�}��דsRq�U�-��e��R,�^^|ZC��'sI��xM�q�D�@o���u.�N��d����M�u�!lXuƐ��O��}�yT3��<��J��nKi��q��_<���;aޘ�E�Y�LkV�V�����kǞ�xx�`����ŻvT8�������� q��0��X��{�l�2X39�١DՇ��a"[���u)�q����4�+�&�^I��*��F�5;%؟Ǝ&�n�%�+7��lU��IM��*�L4���c�cL,��8��M F
���lܸ1��0Y�������+�����L�z���eP�"�� \/��X�͔~Z�ؿ3V��AH1�������ªqs�PJ�v���;�~���a�+g��rNK�>���a���Zی�q�������ϼFX影��J�Q��T��s��G�/�0�%�<�2�=ߏ�DyjhhHج�|�re�ִ��F�}Y��X`�V
�O�٪PCV�F�K�҃���6+r��)�)MŌ�l���Wz�h/��ג��jZUWLf��>o�8!�	`Y>Vl�SS�</�0�<�rfhhDJ=19�p��4��Xtx�6�� v:��ʜ�O��DN�U$�n4ORlCbPbW���P��AB�4A�B�by��:!��0>�����$�����@��挶l�𜍼jUF؜�0�W�Ӹ>���y��\�^�//�d�7�3�zm.7��kΨE���ŕ(C^W,'1k�3
�>�*�S��W�u������ZۀZ�a�Z�km�m��m4�HL���^Ne�/X�r�%�\r�e�}�?̲lbb�^:�m��Z����"�w�j�ƍ,D,+�f��,W��i`��{]�k�$T���E��ĵ
k8^�(��
#,��#�"R,"���(Oq<�r��a�u��m��:Bc0�j]��,���`_�k��F�w܁���73m{��^�ӟ���#�����j����Zh^�]_��m���{|Q��[*.�l�RT��C~�O�W��]^�G}_�{_�7~͌^X��r�5�N�۸I�����40E]鎵�If.�V�T�g5�^ܦ���!��l��΄�_8888�dp\��aP�},EC�g�b�2Azd*�r���V76���N�=3l ӈܣ̖2�e��TUm�I�������ҋZ��0�N��I<كa�:p�+V�[�a��W:NSY	l`�j�:Țz�f*�A`��Z�&X�X�B�Y��J��N�~��Ģ
��I��m��$ڃ���C�<6͒BK���
[�¼w��{�0�[03�C�B��h��$)�n��MMᵈڊj�%E�kُ���0JZz�V�Sޖ����q���T&�<ye8ᄫ6͗������i]�L�x�X�������\O�0��bU��[��Zc���<e�%�}�m�/����-���R�V҂*D{$j!Z�ޭA�vOѼ�L�B�63ЄH&�)���S�G�Uc��bs�ì7i������[լ�H\U[y��<��6s���D���m���5����z�Z����S�,��4��f�����+��=\�5�P�o�n��"��G�U�z%�lP�i�Yg8���<��:�K�i��kXê3Q�MǑ�욮K&p)�Lz�����y#w�d�RF҅R4U�s��V6��4�BFb@�H� ��>��a���b[`T�M�y$&Pc4��EHi�������O�WXػ.�*o��o�6a���~tppxl�q-�m@e��Gn��@��
��UH~,��4r�����о�Υ�����fy���� _�.]
�ԑGy�u�&M��>�Ö,Y2��k֬AW!�d'�,5��^�:��N�b���S1XmUKn01U&U��Z`��m���1~E��?[c	D��,�B��eo[��۰aý�܃Ś���,�7o�<��NMM-Y��W�\94���q�tmi�?���3����As�gn����)�qn�l�b�I�y�،j�;�Yk�&j.����1�g�G��m=�M�q����G9c�vN�a���{8���-�e����Bk�ox f����;���.�,Z3K�Fk�U+����w.F�9� �͙��,�JLS���7a�,py=.m�A��s�����pش���������懇��ߌ�cAѿ�����0kO6����������`��0��k98lT�$*�E�^�2��J�acx�}�zk�5�YV�e��%3����RT���)�V�e�er`�8�D��KƂa?{-�o�Hm%(Ȑ;lV��(D�4S��07��I����R�n��x� Ɵu)-6�(�
ǖ�u8��ə��u'`2	�	_'�Ǳ�s�	ipը�,7�M��,<��ɤi�\���@C-Q��F���Þ}�p0��^ӗo�C2�B�Wn�����vϞ�u����ε��#�3�J�*�y���E����Ƣz_�K���s�x�����@�:��5U#���������`���par�;�=L�����O���s�3����y1���Q;��<q*ϗ|��9�������Ͱ��u�mݺu��{���{��/��j�O����Z�a�U��r/Y~�7/�B�!�u�����n�����XT>g���-iua�,F��N*|!��"�%�D%��Ӽp����W������J+��p-\Њn�B*����u_��ghH4g�Q��w�F���O5�rz�f)����|fC;cMsmc���rp�Ḗ�ö`�{�yE2�kْE��M�D��͞�M��3�N����1�)�E���A���?��N��ltt����hzj��ÍĜd�2ff��hp�Y� 칲Z�N*>L&W�ISU��zwubM�x���Q:�XՀ6d�Y�KP�
l�����jժ�K�<��C����h���!��6X�###e�e2sa��"By$��!W髙�UR�av�<J/�gt+��u��r!��������az.�'��cf�p�L�L��Ŵ-j�3��e��������V:�4�.�í�iӆ-[�\w�5k׮]��!Պc˗/_�l)�Ϋ�	��.&�N̵`zK�o�i�X���)��Ll�	�=P�!�5�Kd�l��JzX
�^��- �j�ߪ���w������*]o���G(lI��j?�q�k���nw:� �P�c�� l\Z=��~�������ZۀBr>�����lL^�YVb6�����<=Ul��t��o_�I��HD4���Y�����l�\��#@��8K��S! ��W ����w���WsC暉u�a݌IZS����#vTVn��j�u���ܕ@Yo�|iv���3�Jr(X�X�lJ���l�2`��8Q����U��O�a�"��Hx~��JZ؂� �a/((�
��Ly��H�{u���,����m��Dӎ���b~�r,ղ����͜��x�?�q�����3�*���R�S���=�s8&�%"+o{������ތdV��ҁ'�Ԓ2�:ZG�&ԕ?=��Z�ެ1�9����D6�ZU�4��.���H7���ʱ� a�,�}e�����mZ�К;n�����ԥ3�-��zij��\���L�ðK�~9L�Z߃��w�D����5���*Xw�����/Gg�4 Kp_�����o�Y@o�Lձ�H���1�S�n���cq����>���5�A�8���*pG��m��B�Vwtt�������*NWZ: ˀ�jy��-m#_���ۘ�d�^�jo�6���L���G�,o:ӌ����*��p\��a`g�坷�����Ũ�޻�:elZ��$���Xx`�u��sϻﾻ��yE���7��t^�y�/���$]M�[�����ҫ��j�;Ҫ�e��3��.�T�N�������eq:V��|v�W흫;a3���gY�����OE�a�]h;�H&#��V'��2|�ᾳ3�3����D���??R�)4#~��S\d#�鑴���z�i�n�w�KP.�iNc����e����h&��z�&�~������Ƹ��δ���4��{6nzp���`4 �U -�A�'���JS�k�B�]<22�$�D,�	��$��?h=��-[��&0�����a��aﶪ�P����s��95��N�_��k���t{��]��X�tr�T�\���h|-�u����x���ڼdɒC��dv��.����Î
ǵ�KAp|[���)8mAhry�ZFT�+χ���F�ό�E�F,�M{)�Q����ːKQI��d��$Z:ҙZ���������v��B̦��M{t��0�mCCVV��N�*#1�_Յ���N5�-��*;�޼fYʢ�d+��RU�dQ�:�Vys�ׯ��A�C��V��l`�I�`;���d2�i�L�fI+�J��p�ou�۴0���rKx�,_���@�/�����qqu�܈5��_�jI���������G�x��O_;1?TE�f��f�?=A=��*mO>����i�$�y&��q�U�utuU�5� � �-@2����h��4���_ ��$�2�h&.94,m)b��!�s6����#+���]��U�5��î�FNVd���_�>���� ��ֆ��C�5�eh����:�D6D����nм�EU�+�����z���H���1|R:qg��sk�qD�1�f{˔�`5T�ڈ"1Z��x��w6>�˲lЋ�`y��N�������Ϡ������u]FA��g�yҪSYz�*��u
K/�OѝOZ�Z��~U.&�C$�K Z�dV[�8;;= ƈ��20v�^�O�!���w�4Mᆀ�	pv!]���q�ٜ�>^��I,WW��T]�2��zj��|���<�;;;�����������yKQ*=2�mPz�����1tW�g�d<����E��'�ۖ�������Zmi˓Y�4��*�
�ȫ+��/W�{�Ӻ*�y>��j�^8r4q��R�'�ds�l6[ZZ�~��� �����#t1tP)����c��4���v���hJ8㕷Gy�?��|4�a�S2�}���B�� R�Th�ۦ\���Z�����ʬ�GFx2p� ~X8���pS�F|;��BCc�V�y#Ydk��q�����[|��y�^]�����V\9�>����O��Ch���)�y���͊���P���N�T���n~Нy�\���W�I���1ᓲ�����v���Q�FX�)����}��l�b�@�����F�:���ئx���/0?��%@b�y�h�aJïp��O?V:��c�0�T'��� �B�
�=zG��3�<5_�v�����'[��7o�dE�q}����JL&�RPU��eV���Ӽ���Ep�5̤g������~���O~��/�\�AVJO��+�O�m�!ElK[�Җ�,-�jK[�� RTS[/��O�����9�l2� ��D�L35�;D�R�H�3d��z}zu�QbTN���<����(0�,¥���t��D�"/tj� �:�m�*�sX�X����$.	�c�p�	?��F`&��<�\��9�H/n�M9���9<=��6ű���1��}��p���8;�%xV��UQ7�P�����x>��zI/R ᪴��������,GhK@WH���/�{x.-���Ɓ����A�rF��$��C�s�8|J]M�p��@�*�}�w�������Am:��Ƙ����V����;J?�q�;M�Wi����������n*�Q/;dcO5�������b	��.@���T�R�T�Y��]�0R����it_un%2/uTOZ1��%63�Z2+b�h\�?׉ϗ�@}���l)����$
l���%�_����֑�j0�! ����F#��°��`�^���K���H���p��64M�S8�e-T8jkk~�?�W6���jN�����O*�R_`�C�p9l"�''Y��J����dB�)d),�(;�hEi�Pf�N7L"�-&I�/��̱���������pee4,mM>�ԟ�aį��3.G�h���T�b.a�_���(ː$53�dP�&6�猨vt�]�	��nK[��_vi�V[��%xs�$JBzQ�{��a�A�sY"�)�Ņ������r\a�m)+�<A��y��!��ʣ���-�,��P�� )
��n�{69f��ꑤ~Q���<{����S\6� �1��i{>�H{����娌u����sw�	$�ic<���7��׸�%�,T!!:�m�0�\W�K�H��^e)�D)���O�.�4so]q�������-e�mQ���]{�^1��M^�c*���cqa/�˄�:׌��.NO5O�G����P��N�ˆ��w/��W=ˈ+�� �Jr7��?l[Y���Iy+eF;'�^� �jp��m:�VOD.vF1��h�)!�#e(V��E���S��,�&�-�L�ǚ����F��%F����l6���"�����́�<�r'1�Rb��p8<88��)�����r�٢�_���gN����ڍ��\kkk+T8N,�2��f �b3`?�I��܄���� ���Œ0܂c�0�����}�\�O1:����{��}���G�Y��S�'��G��������eÖ�XcTsw���Vf�/W�+���:�.n���>b�OR��"���y��9OzӶ��-OZZ�Ֆ�<A�8�R3sqhм%����ߞ��H$��_�%�L��Z���r�J�@��R�xn􆎿��݅�gU`�_L��: hW�&/.���o�Y�,��Hf1S������!����Wp��2�u��QE?�|QK���P�)]�[�W!H��Mae����pܬ�WR�PS=,+ǲ�КR�6;�8+��?|���z�����Lt���*��2dMs�f.�z��O�i�D�ٵ���`4	�Ʉ�6]\�ʪ�%f ���Qz������ՠB���@��}����ǖ�C&/�zYHT����ϑ5�¨�YY�0����S+�N �%Y��*wt� [b'SX�̱H��eDe`�A�e/��"��`t���I��tw)Ȫq�f��n�n��XKүU�/S�� ��Ux]%�ہ��l�F�v1�YQ��6��@�Q�*�u�8q��#76o �D�����<�N&hf��Q���SaJt2,���Eax6H+�, ����% ��KK�@�b>��J�E�1e�7�NKR�^�&gg{��p���
��K�!�n� ��9Z[^��;<<�gRµ{{{P	4u}s��ȰZ�^�K+:"�y4 O��� ;K����� @�$]xvh�*l���^9������xy�"?_Wy�=�}�'�e�S��vA{��|���8��N#�)^L6a��H���͓ŏ=v�8����}�UJ����-OTZ�Ֆ�<Iq�����Ei���`����|\�1�V�pSR>\F����S��R�.kyB?ݰtYg��'�TU��.��]h�>�Q=�����68^YY�jrF �)���Ѫ��x�C������p�BC8�A�@�i�Q���V��g��� �G����8D҇�g���|������~��b>�8�N�Q�L*NL����1�E#�E�G�D�S���V�ʴXԲ�Ño�-]�2���6�gmB�ܷT{�����\��E�?��d��lװeU��VVU�+�!�jJP�4����lP��rss���������T�4xV\���l"�(y�/�n��رE�gE�.���% ;��j�"�.��{�`/DIQ|�l��`5�U��r��Y��e�"׹RڙJ��{���2�$an���m��+�n���Q�C��i(�өt)�`n{�.,�^��_���x7 �����0�ONN�UP'�;���Z�jwww}}���İ1�^��*a7� ��y�mpm�(�PL�.���o���c� �[>ίt�Ura�9�E\���ff�"߸��>E�������\�I��W�9���?�����.����nK[�K,-�jK[��sID>�*�Xu�s_=Z�v{f����Q`��JT�$�[l�0��'����X�l�a�B�>]��S�,[C>�f3�(�-@z�j��ݳ���$��ؕ$��V����$����	�q�����Ԣ���Q�\ֹZd%�Ǳ�G9�,�ZȮM>)*G�xі%Kt�"�L:I��(��H�sȑZ,��GC�*Qv���Ң�gR�jv<ݹ�gK�<>@��e��-��;����],�������0����]B�)L�$�ʘɵ��[2[C�%���+wZ�t�=�<�8����$�����_�R Ҕ�����e�	k ���?��G&2dh�ؘ���8+b�$�f2:TO�O��a��Ÿ���i��d++S��ɾ.tZD*��w��IoiXD��1V�,��?�HPyt���V��Y�P�"'�wjbU�1Q�\�ӫ:+�JU��@l�,�n�Uj�/l6���E�kk�.a���׮�EYd�|:�Z��I�� _>K)�t^h��Ե)�P_F��!�z�*������9�Љb�*�c�(c��X� �zI���[�<��K��.�sr��J�9�NF��:q2��a���v�~�py8°O��l�C�]�g�����,w�(`�A���A&P�����R[aj_?�	I�"���W��$g`j��B4�W�\z�l��6w?V�Uw���DЧ鑙f6{(�[�ȏ�d���>���BW��|��{�rUS� �D+ז���YZ�Ֆ�|��T�0��}Lɓ�3VT/--e��=T�K�|�yQ�*S	
��]���Z�������d�,3!���A�-�#��9Ex#�/��}�	3.ha�����O���_�
��.�������>�W�7�Ro1� k���e/܈�u.���U:i� �2���(u��~6��	��s��������R�4t �Ys϶)�R:�Vi�>�>A�0���L7���!�/�I�.��#c����R��r4���Y����I�S-���v��9��O����9�.����ؘ��x{��ިB�dm�Om���1�����cK��֊sĽ]�i�6w�E����o�-���������Z��ŭz�JNR2�z�u:�Ӫ�#B��}Ɖ��͡at-��(��5: ,
k�$;�G�����f��A�c�;���������������ɵkנ6�r�]�V,��(K�$��,���co��������l�.�t�	����^�vZN��$ ՠ�7n@����p8��Y��b�����d3���Ӡ��/!��|�����9����'Lh��%�Gc}
�����o4+_*L�1<[��G�u�'|�G�%	���MT /�l~�x���%�í�v����;���c��]�p�����b=�Wv][�Җ�]Z�Ֆ�|�R�\HAMa�Ƣ 	�[���N�r�g=3�s1��ݠ�������#�K@�%	��"\�P��eٚ�?[�
n	�ڠ��Qd�Nl$�cJ��@=�rT��:��)�D1Ei�JP���uџ���}�U�US\8��(���y��50�A�i�"�(c�)ɷM4� W�<�t��l�s��|�H�$
�I�U�>�����N~�׳E:�;���EvBC,��rh�Q�WWp;I����ʛ�*E�F�D^O c���A�G��hH�i�a�^J�>�$�5�.|��]d�4Y�����c�!�4�t�,�����K�s���U�zv��3�K�01E�l}���G�l�ӌ�b��9�,K���:�k�	�
jg���\�1�N�޹�X;?��V�F^lY��V@Wr�����m��Jϯ����=F��1�m2�E|�q5"$jMI�'��{R.--Rݼys6?z���ߺuKa[���<h��
'/>::b�^�� �#mz�� �0�| X�\K� 5 ���0�����>�������]^n<�;����3 Np��b����%�/�%�#+,|N^�	�o���]*�HQ�ld~x^���@�A�黆���� ̆h-,4��
�y9���d�Y�4�L5Xj�Ț��qN�6���?�q�"T��Aw#^<�QN��l]�N
T3p,��_d���J�*��J���x\o�tQ�������k/���u��-myli�V[��E;}<	"�[3��E�=�-@����$�&,�O:�kA���uQR��w�nS�kU I!���:
C,�Dj2�`FQE1�L�?�f3�70ܥ���!���٣v8���5ӝW�7��:��8%�:s�y�;��xL8�v�X>��%x�2�6���E,�t��N$�qz"8dM�����c�184i3���r����8y4qo��Ώ;K��qSc-a=D�N!\fꠊ���!�������{j�-�����|�;�)+@h����T��I�6c|��T�`���<+�"�\���l e.>�--r��4��5jꧦ���4�C_��U3�@��t�$�?������x-�����͵����`�X��&r�f�����X&^V"T�S��pM��	���QR�� ��Ե�!�ᕂ!yG�>|�P�ɫ��.24@����~Z�U#�5�,x�lnn޸�����P'B 9�������a��Ys�AK8o @tpdooμs�λ����ॴ������[��`nÙp�۷o�����gP�y8.����z	��6^^w�'[�x!��5@���2T-��7��ps-z~E8�z���o��f��:6Y^^��W���F3�O���Ff?o��7Q�3��hƝ��1��a���Fs]˰�71Y���������
c��\@����ȫc�pӧU����
n��y~J\u�c�}r�㧽hxj\���[C���Җ'*-�jK[_�{��4��jE��5q�KeX3�Dd̀�KE���y���J�Д�LVZ��I�JE�R��dH�%y�6V�)��$���شC%��U�E	��gYj� ����ds�(ln@A�Z�@,J�.V��,7n�s��4l��J�d�$&�'6�����5�{��rϐ���xn�u�],���M0�+��61�D\�R�Q@9�4q�陲kRtPF����+����RdpH�B�������.6��:K��`�I�Q����D1�a�F��-�W� dB�6䱄	�i��ɓ�=��~�H�+"$�*,�U�K���VNg��2h�o�e=7�pB��T#⮔ul^ �7?`�a�+��*��IV�-%� ���Ⅿ=5�y.ڈ=�!�i�Y�ő5��y9 0��u�Bh��I	q�u>�ո�o���l�Fl���W�2�-B�@yGv�t�nr��nN�ȪWjjs��{�b.���8�x@��a��5Xz0�JuM�E�,vs��f*a�e��;}N�V��H�y�2�&�PM��#pOX��<��f��c�	��xI�C�\�
(k��^������ Z���RD8���ݛt;��(h�btX���2Y�)���<�gY$BYh��<r؊L����4[[6"5�I�iѧ13�Y���$>쫲������+c��&�j���a(i��0�J��r)E	b3S�����<Xa�4uڴ�ݞ�}Dz��%�W�u鈘^����~��~�#��/��#��-��o��B���(z�\���H�Ƈ�E�3$�`X�t���Q$aS�q�V�3�*�-��$�|�i8:"���,YQEoV7%;�8��l��B�;;j�']b�����$��������|x����
Yl���-�)-�jK[>�btbmn3
"gk�2)v+T�.��j�%���q�(=�Ew�����ºg٩�	H]Sc(̃�ڰ@F��O8��V&��1�Թ����U,�sH��c��ϗ.�2#�fTڸ��M#��~l3��!��p���%�H쩅��b�L
��=_�A�����;��&��m���)ٲ*0��b�iW�˳d�0�!��#,畂L�l�$�T�:Y[r45?$�K�P����,��F���:�c-��ǖ����5$ȸ��Z�m�������"���2s��w�ސ=M�Δ�4e�n�0-�K��˰�q���-	��X�#{�?h�t�ƹ���aN%cE�t2�9Z	� L(�!�TU���;��2����p��f(a1 �/C&8�&�����������	&*�5�U'''<.p&�ω�� L'�?��X����8��ݻ�ӳ�>�<����G.|��nݺ����5��?�����g>�
�_�:b�ȍ��B�X��q��A�y�s�V�Ty�C��@�5�y��Z�i���v5��p��E$ɶJ��vW��C[�xVa-��Ľyɛ0#����ʦM[HM%��a�]K�:��bl�B*q����?�J��<���w�߿�m��'�I&
�3*�� M#��6E�%^��E�e�F��B���:I����s,q�v$1-E����R���^�.�R�]����BX�����ׯ㑜l���P&��c?��+�+���(�^&�/�KZ3W[���Zmi�'P���A�J%q����A�"ɇ�SI��O:ACbi)C�CS�_�/0#E�F���#ȹ��#�^Zs�����2*%9��<ͬdy��� �7�G�I��̢�(���G5
�I�+����O���؃��c�7�e���:X!__�$���f�=s��"���!��m�B���Q ^,�{Y�I�Hg�1X�A(�A�;�&F;l��X�TEx� x�*D�ن�Y��H�,{��'Mt4��<{��*8I�B�.bθ09�G_.��ᠶ�vX�Z�"��ij�N�4�Ȏ��ZV��H����E~\k<&lD�	���Q�@�����>�MLs�h�jV�s�GmhMVX�PM�"��025�q�1��=}���+R���+fE�/q��2�j�gEfs�Q�����J �4��ADR���},(Qׯ�sA��q5 ��e���9�F����m2�@'�~����Џ�	�"̸�$p	;�/��:w<�L������������'!�Ȳ効d��1�p2e���Z�M1�_�Q��1��}�8b6y8ҋy���S�7�HQV����0�C�@.����&%Z�R�t���12f�D�Ŗ%�Fig�
8��@�����*��R�2�Zi6�W�����ʖ�&�fimʼf�au��l�1�����L�j�ߵs���d-���q��*Lu��Qn���BW��d1&H��,����*�����o��J�!:q�����J�C$�O*z��'s�`������N�k�x��(�4��ݳx�&���:�4`� _^��)��T��xn�lW[�rUi�V[��	�5� ÿw�va9]/y�)�_�'��^��%�#��ؿ�a-�.��]��By+�R��d�U���>f�	�ו��K��x�y��o,*���a��"��� �]��7PDi��l�R �tT�ƅ���58D��R,�pT�ve܂�S4~��SD�Q�T�es-��1e3�$�;�p�ym㎍��ZU��$Ӱ�U��ԍi�����ޢ��f>���]������5W.[�2`]�u�q��e�*�4��xＪId���ڞ�`��{S�ȯ%���VR<��%�c�P���e�2��
f/d�hqk5�vS�� 4Ӈ/�� S��0&�[1^�#��Xe�X,I��ES�o���X ����6eõ̖���1p��_��L	|#6Xq�p�����	�H����s��4�^Č�tQr��(��G�Z#���V��)���.��jaRf��6�����V_\�87(�UQ�t;��P[U�����*ƫ�,��y>yŝ��5��^����c�H+�g_C&FI=��T�X6�Q�m)IW%pPٮmA�ʦhb-�ܱeU���j'!� OdY�K(W������쮬)�(2ŘJ�V��eR�Z��Y�9�������/��b��PU|�8�-mi�G�k��-��B���,l���(7�6d� ��Q�b<�t`�.����F�e�z/\҂gb��9���ς�^͋2����`�Q%)H�a�i��U�HY�KtӇF{AV4H�.+$)�)c/�A�`E��[X�:W/R�J[6�����H[��d�<^9��r{�#$z2ֲH'�`��;��Da���"��sj�C�\��  �EQ��X� �:��������QLT�Kuvi���k�D��3ץ����n��
��_+;�a}3�F.ɏ�GJ�,���bW.t#"����EcQ�Y
��kH���]����h�ݒBy��u� 
�Cԓ
�ߵ�0i�%���Ҩ���z"YșaN�Ly��
K]Z�J�钰Ac�j��Z��������Q�t>o��#\e(s�1��y!K87� �Gt��wB�Y�6(P˒�[I-a��X"9c�Q�Y2O��8[��Ԥ���^��Z�'����NNNധ�z
�ÇA�_ZZ�F���2|b�c)�0��`I�C�� �3�����K ̠��}��ݻw�Z@\���9�=�5�(!��\ɼ�e^�6C{X{"҃���ͧ3��I)d�T >��bQ��iS��� �J'������ w��xu'h3�т}�7���oױ���1�N���[�\}����GT\2�&���,;l��Rv�0Yd�(�g��K��~B;B�K�'b�e)~�R�z݄,xȼhD�!�@��zOf�C]�D�RS�Ax}h�%X��)>�r��0)���i�![�)*�t59=p3���!�X��z�㳥����K:�YVr	�����؄���I�hK[���b����)^��Lf�q�k�(�J�5��R�y��+�y��̗]UH�b�hL��9��4� 6E%�*�|������uX�W�*�H&v������ \�i\�m�a0a���i꿽B$�
R`�P⥺���˹x_DVϳ�p����h���dk1}�����'K|h2h�k��[�V�}�d�HF��c���+�z#��Q��1pP񘑁�IK���?aKf�f{N@r?��y�wᰖ��kk	Ys�0�9��qs�M	�y�rl���X:K5��]R��3͉��� �a���%[���B���{L.)������a-[�y��F�5�LHX���h�b�B����I:'�"]�;P��A�mJ�b��@p��*SO9��  �*�6�w���g��*�h�>~���'d���� ���#��tF�Hp>�������~ZW)�Q8�a��=�&��p#�b�غ�W�M��4W�a���|I
n9��h�\.����J5�U��pHTy���gB��J�p��p2]"}6�޼9��u��m$^ws���x���m�،X��&O!~�n�A�Y*8%�
[0�jy�a�ĚG��Fp��H����Z��*�U�dt3��(X�+� ��cf����.rD�{s�(� a�il��ob���hW�$�Z3�0�K!�"iK[��b����W/d��c�u�&R�t'
v+�#�H�A�5f����Mق��u�in��w�^��Ӻ�$��[P^���a0a��n��^����vww��xK��"��(��_́��'�6�q��ܷأ�_�^�fA�O`���1sm,@�����l�"˶���7���5�<K���.Ci�4�-�A=�#&c��D�O]��dGZi�X''a�e|bvu���f����׃1!�	M�fL������[u8'���Qxw%H�l�9� 8��b����Y)�T�=�����,[�CXJ�L�K�̀fg���w�{�IN,F���\l=����d^��uPF�sN$�Q%`06��!"-`��	��H�S�}��*r4挢�У1J��EϬ0Δ��	ۨO�L�TY�JDV��Z���43cf����---E��.��Q�p�D�/mI�=y�R����k�+�0��=׹��ټ(3S��4fy6�̄�!�a�yo<�Q
�*����0�6�Ċ�GxMp2ā�hkk� r�k9R���,��`��U�P����['�� ��g+f�y�.xis_�c�}uu��/j��z��9м�D+�e4�O���e'��q�&Z�p�'��\�5�v���KJ�L�!M;-bj�̆Q�� � D��B*d��:U��ڑp�i�MXuz@�Zˠ&|�jmy��tm��@��qq!.�Luя {z����{�3�˦p�"E�W�?�~��h�#|�5Aib!;VDhɃi�by�V{)��ZVe��AY��&�&ݐlV�v)�"��.�!"��Р$!�!/E���.'��H���dW�
�y	�
A�A�瀽��B
q3�)ĕ깶���ϥ�Zmi�'P�Rп��AÚ�eE8�:ŋ���rDU�B�Ax���� ���*�c�2�9� �rQI�����w�D�כ˚�����܍��_<F�WV��Q�y+yi�WՐ��o�F*�҅�4�\�|��K4�9b)�h�"�����r���8:�v�1_�p7�����dlA���f�=����F�NK�ֈ�P� !�=3�k�@|���"�SsE P�,�x/Qu&�a�;�dظE1!y^4�Vm>�&��U8�O��-)�-� <�"��:�0�&� /2��@S=[Z8��t�;%�=�I��6��j:�6�Vł@F�(/ɀ�K�#���)~��L���Ns�^x�Y��-�4X1����2c.�7;�2Pa'7KY�8n
��"� +�lv�����KI���ꐲ2A�����o��8$̒�c��3�4Nħ�9��^t+�/�.8�m5������~��mJ9VΕ�\z����M)��/&;��u�m���t&n��C��yck�*��v	+����,B՚�|d�hhB�9f?��2�e��>�NY4=I\�hrW�L �Z��~,�{#�ByO#��j�0�-��a��|�4[�7O���v3�k��\���+r���u�������F���ڏ>��\�2�+�Җ�\]Z�Ֆ�<Aa��*,�I�R�h�I)�mJ��
��2��!�#I�1>2m�0��|T_�M1+Tu0���iv|�(��\9��U!z�̑v��xl:]�d�P�=*�ȍ-�5e�Ab����XHj:�X�!G�4�YSv��Õ��f.rx+Kʧl)��l�zq>�4ܟX�cy4M�*������[�2���$��(LOO9�(K1��R�*�nAz�'f��k'Z�\�0QwV
$Q`����a�d�h�ɐ'�D�@��}#�lPҭx#�S�9ϥBÓViUɃ	�)) �q�z�����%>��@{�`i�����e�c���*ҁ�P�,�q|6��)�:���0x��r誄dVK<�������y������L�� t:��$��YC����f%�I[�A�rD�����;
z���h�	�0�!�F��@��	��_��f�4��H`�����OI�!7�l��1S�9�:��ʸ�\����sU�c0N��h�ˢɬ�Z�����1�E�AtIou=�"����]�!� <�ז��a��c{R����b���Z�Lfs�)���0�bv�l��d'g0�ǰ��Bt�N��K�u��bccj;>>������аO/R8~�F���Ja�r�죤ж� Y�g76����&�	3����������������i>�9��~b�FtLԱDڶpecc�ƍ̖�� �l6G��Rooo�$b�\���8C�R���T�8���A�D.u�,#���]3��p^,`�Hmnn��{��� h�B;�Й�S^)��3\A�QX���H�p�
�4S���A0e�*�т��W���y�x����f����n�f�<_ ��Z9]�.%���w�F�}Z{��ں�����f��y2�y�E��v���1h��Y���I��"a%�� $1�㝰�=
��&nd��~�6dc�v�-Lk��]�}QRU��.�ȓ_�L+J��
�8����B�8��Y`<do �Ͳ�#{�~/������h�c�xA^��hK[�r��X�-my�b)�������Ĺ{5��l������I^��K6[����˗B�%U�Q
E�mkA��s�E�����`w��RS3���r��S6�4��zݪ{���tN\�y�����׸p,�3��,��c���C�������9�v�T�^O��m�4ʆ;�G�XuB��t�'����9�q!��U�B��$$Ԧ���=��������O�VWWݥ�tj�,�����3��hIA,��]b� �L���̳�9��P��Ӂ/ |�������8��#�b2��D���j>8��͕|�?��V�O:�:��G�ņ���H���Q����R<�-����{�C�l���Z���~=�󬘲��Q4�'KKēnt|<��q{���@]8�Ċ�A�!Z�g�
��ZXe{�k��Fd��0Gg�q��}��oݺ�gz���)x تi\H���K0��À����b�g�b�ۤKp烎R�;�5`H�ֹ�
�Y���{�������8�'�P^�7������jg��>�TM�۽�%\��a��2"Fq��1cX� �iS@�&''E&CS�;�U��	��i���K9��j�ijqt�І�^z	���������X.�������p>���'ggg�>�,�>Y�'��O�Ȗ��Ȩ�!����#~�=%��3��U�{5�+a�Z�W����+W9͈8����֭����*�[k[CV[��D��Zmi˓��8�N"�6Ԙ���D7����%�5��D�'�b&6*DB�V!70�-ҁPq)M�_���H��c0b^�
�I�c�C*�v���|0_���[۳�߻����`>�ke���~�K�	�.l^�
+��g�n�땲���(�_�ry�
��Ͻ�Q�?���6��x
���*	)i��N�7�����%Qn0����H�����RFr$s(�hJO�ɵ8������&Dl
����6�^pf���I�%�QJ�Q2�@�~���L���y����ى���zk�p�7�8�峬�v�P���� ��D1�dXN��M&��� �Y`4Ȃ��7�`��$��E����Na,V�^���"$�h��wIj��d@�$�5G�-�3���l�"Z7OE���2� $�G���VV��$����4��G(�4X�P�a�-�Rwfc角�m�Z�sȚނl���,e2�Hjl�H�@gR�:�+{W��`�;[�K�d�w 2�@E�,=�0�%A"
+I����JG�B����Rx�$��r�) H�JdZ,(1q��M���Xł�ԂP���`]�$x�Y�AV�L�R�TP	���N <��9�1|�	 �`��������T����Ϛ zL~��f�og׮]h� �� UA��*8�5s�tf�8����muB�fGz-��k�dzƁ����6��2C|h4z�Z����0�Z� ���0�adn��"[H����`c��$�N���#��%{zz�(�vM��d�@S6�U"xŚ��內5�֘/
Cd	c��̭]�nV־������G�k���q}���h�LΊN����K�N^&oGj:�H���~��ouo� ���S�?L����"�аH2��N��Oa°*kYԉ��b*��W�Pդ�������='�
��ɕ��#@�^��̷ʩU���wE�=0;�O�t�-F�a�N�\�G
�k��-W�k��-OP����nD�4ш��p��>W��0�X
�"T?��ؑ����	!L����TR�dn=#�L	g�i"����i�:g���jBEq�|�O��IӤ�u0���z"8wS�O�����l�o�GG�G0�]%e��Dr%E��+׃�;H��~߸�ͻ_���]a9�DCml�:?m.���n\��#0�^#[�׾�M@ i$O��?�Ϭ��y8��ￎ������p�,���Ű�4 P �,�Hcp|6���<D�� 3��,:88�:�Aå!��Zw��Ç<x�8F(k^i��~6�&� k�%����?UL����������5��h����r�)V���w�����AT.���,rN�h"3W�(�aM=��s08w8U3�#Te�b�����9#Ӭ��q�X��hTr)��ِ����%~Q�j`H��D������a�ʂ:�
��-��ڂ��p�G��~�:7����yRAU��gGDh6�>\��0�c��m^�p���!óy�ݸq·����ojB���P��2�g��Ab�RR(�N�rܩQ��Sj���Lъ;��G�&:�W�ao����G����#t}�E��pu�v^d�桹/I�{�t9����r��@W�R���n݂~�����Q����]_]�����k���h�Ѱ5E9��u��&|0?�j��]c�!t|���+p��_�)��C #���Rp�b=̾Hy��7r�[�y��l`��W��Ⱆ?���rXK3�.��r��Z���ꎒ�W�D~�o�����-OZZ�Ֆ�<q�htak��^Ӝ߈����We#�H�(��l]hx�G�O������ "�$�[R9tg���ɉ����������k�Yyz|pvp���1�Q����?�%����<��&���EPֵ�J_[�Ȇo����"�<@�sDE�`S����n��(ǫ�n����r��H�J@�B2���Z=>>:;Y5�`��"�G�r�� �$��[�|�ɅJI�cK2�P�z����q.�!�$�� �̍��E�uC>a�4�f��]��Ͻ��Ƌ�����wUMN�[���W6�|�7�<�z?���n_����q��B�D�$�C˶�|qv��2���K�5�wE/Y���ܫ_D)3 ��dZ����x晡��NNJL.�4Y��R�
�f;u�u*m!�h	��-�Ʌ-KJLRH��&��B��W�����gG'�O�zK�7�mޔ6��������߃A��9�P�oA�c8H��k�6\q(8֑쨴�舩ҐE�y���E�޻?�	������Y�4�# '�z��5!����iN��e�A��{v������~��[�B��t�Q�+`�v,�5'�e�˙�rx�;w�01�7�ȋ��t#yBW �_A������������W����8��A'd���/ �`��,��jȿ"7c�An� ��;;;���L�m�9���g��-n-|��R4eK��&$[+�rI@)��]1�8����}xj�=����Q�t㥑��ѵ��2�P�Q\7鐺�1`�FV�九�yP��.��­�(�\� M�ޠ\���b������8���'a4��n~��A���a���$�Xؼ&�<	G*�갃���z�i�y��G��p��wv�3;/�0�-pZ�j<t��5�H��i)@T�zǫ�X�M��n��M�e�����u$c
M%��M��E�# LU ��"[	(�lt�1��A��L�����~f�T�ٮ���-�J���Җ_�X��ִlT�š�l���
�w���KH��8Dp��'�+p����bK��ʧ?�iu�&HW{�9�[�]?B'�	��yT#�c*���<A:��ZW!�������U��L�-��(DD�q5�yl����5D-,QnC.��"�EH�_@�
��A�E��YW�x� 5/g:߇��|'�㜰�ƫ�W�����:�#��~��'?��| M������}�����������7���׿���.�����I̅z��goܸ1X[��ڂn)�����?�!t�l6�ÎdP��Y\u��1X�,���Û7o��L4X�1�[�Tm��. `ٰ_1�{�9t�-���\qŭwzz���_��>�>��$�9�g`��$N�O岮���w:�\)MFDgg�����x�{f�`�_2gd]0q�fyP
�!�FMQ7RE�Pg�̐6N�w�����R�/w�8���g�vm�/T��!�����΍����e"�%͛�a���w�}�c��ZŔ�p�������G=|�v�W_}Nc�A8N`��?�Oh9L&���l��K�h*t��pns�&|��~�I㩊�Ų�"����مO���ʒ��,K�����i�ejN�W� �=�f�K����3Hz���7�����7�x��v�.��/.?�<y� ��C��4	�������t��5�lf��|������ ���Ɖm�XA���p�d>�j{+0v�`��G�D���#ZH�����c�]��3.ro��#:uk��oH���O��N��8a���-8fRQfҖ[�W�]���-�<7��U�1b8��Hڶ��-W�k��-OP<����7�d!�!t*	@5��0-2,��)�O1������${���`�;����}���1@�l:E�X��KI���������:=:��֬���!�:�깚P�)�6�Q����A.x�|Ƽ�p��<)sDf%٠f�2/XW=����&�bB�~�2��F�$QqY���L��+��n�@����{�qez]y㾌ȢRa0�t(��t��>"�2�����s�O�_�F�0�;]b��^��3��096G��^|���������(��<���F��h�������G�8 ��<d�����y���ݻo���||2�;;�i�U���0.}���7��,K�}䶞O�Lf��0�k��a/�������r�SUx�%��4�0-��O1�F���)��,���p�>!�a������,�M�N�	K4���F��z�ތ����r�;bЈ�6���U�Y٤�����|~zvR�bFAh˛�H��͓����:�)Z�&�ؤI�n��;�`�w��l�e[O=�3��)W%a�0�3,-�.sZ^֘ X��u�����,�VyJ�ѥ���-����O=�{�dz������;���o~�]
��(���k�"��O�·������f$G�'I�p�Op�dS���/dŴ�e���
0EX��&��fa�8֋���`^l�@�Sj�at�MEa)c��`$�~��ys�y�˝�#��Ф���s2Ǆ����<�s24R%A��7�<�z�0:���CA�9̗8L2��V!�^�"�w0������.}�k_[^�ux|�}:]d�N�3��4͇6�Fz�Łнb*��~��ѵe8|��3�#|�"Eb��mM9<[b|��t
�	]y��	�5��o��Z��VP�9��:��SJʻ�ˋ�eՃ#h�����J$�	��$e&{�=�I�r@$C^�ݒf���.�]�����,��e�?�6�:'�j=�ҖǕk��-��rk��~p(��c�b�B �V�yKY'��x@$���!i��U���q}{{����������L]��Z������T4��l��x�䃻.�255��o��iL ���%;R.�P%%e�Ĩ�(����1�cH�����9�`4�}�ҔA�
�2�],�sF��7rc]������]���<��m��� �7��c��믿����۟���_ Q>g�~��_��������������G#h�o��o��o�Vgmt�޽���{�=���������n�BYq�>Q2&bC�?0m=z�U!H�a�9v��E�jh�M����;���V<"6B^R�}�����G��*=oll<w�Y�onЪf24ޢ.:1!�\�[o$�Kf\�Qq�c��_�� ��J����̺�eݨh
����l0�R���+���/�:�ޖ��!�NGt{(�vz��\��#������$[�z��3����"z\YY��AU�I�R��hqhf���=�� ��Z���9�Ͱ�X��Ç��23n�C%��ۿ��/}��~���4�>�~8�3��v���������
����~��w��я~��g+1OW��S"\~tt�.�О���X ���s�=gB�}�����mh�u%�c����[����s^�І�	 ����_���ry�,��;��֭[��=����}d�?<����>/�ĝ��l��YU��X�\cg��=��dcmuu�7=}饗6o���?�Ӥӿ��[�w���`-o:{��Aap�-����� W�G;� 	ev�Go͜���1Q.o"fd�$�P���P�S4�ƍ��t�*'��>U�pX��s�Le���b ���*Z�sUQ�K�%���)�)�~���-m���X�-my�"CFA�as�I�f:�d���X�ҨD�b�!��!q6�7}�Ua��Ȭ(a�%qwdA�O��#AK�#5T�넨���s���MV��*+�.DS����a/�iv����_|���W��������O�u��J)��d�<ɢ3S3�a�e&�H«\*-�b��;{)GF��'�C�7e�y���y`"�S��ԦNi8ĝ(N5�j)ʊFP��Ts$gĝ�o:+�1���.�ya�YS�.������$;����ϖB
�)�4ˆQ���7��Q0�`i���/0SP\b4� �m^�f�	��+LP�	�oY��aд(��Lv��������*8-1JD0�qhT@���t�ɋz�Å.��������S����vG�I��w�����^�O���does�h�������
2�����W����m�<<<�z~����b��^���[����;�������o�m�Ngټ��9��;�@�����_�o)1Dd�����I����!U�\єp�� !T��AG��j��v:�� (Bǩ�U9�gy�Q���[����糳G�����͛��c\l��,c/Mr�|�-`�E�v�q�K�xN��H���p"�v�N'[ _���]K�e���0�p��<U�2g�����b.����tЌf��:W�⺵�J��f_��gm����Q� n�$Br�ε��,ꭼ������W��ۻ�����Qn�mM�	�m��Z�ē���^`�u���~�~_@܇������5�0�W0X� o��!��?��_~�嵵58��Ν;��8��#�Sh���G����������=*_���o}�ɏ�駀�����_��O���o�n�u�����d�`�ؖ�{�%���fie��.����,���`y�q���v|2�
��,��Q��#��_��O}�S7�y�7#dxW̴�2mllb����wo������9O��Фƹ��G���߆����~�`|�_�b�����]CF�R��������0�)�_hȜLy2:H�� �V}��y,2m��k�|� ���tԍkw^x�3í[R-�<��/������/�:�s~���_{���;'EQy���L����ګ��F�I�W��wogg����0@�[��꡵g�3-TG xR�W!)�
;��Jia3�I�;�"c�=R�Tq�����|�i�ra,.�2(�-�eĜ�'Ҫ��a��D�� ����a\�� m�=`�����+�_E�"��ܱ	:Zw��/ܨC�
�mi˕�]mi˯Z\�Z�ذqy�i1��"UD�	����x��"(Ni
'pD;jF�lޢR=Á.� ��|o���a�q����J���M�^04�S��?޴}�F�+�c�\�����rS�#xd�1���m0	ds|������]"�S�����u��2�9�`�W�������f�h�!�>pn(��o__��_�2���^�~�+_�ʠDkO��Yw���h2"<�[o����� 7�yv��]!�{������pB��Ç �?��3�@�����u��%��� \-F����
��0nD(�<��"���9�-W��N��±�qA��%姊PCj���|�\�"������K 	���	�h�M�-������ 9�/��� 6?��va�I���[�cZ�pΎ��W�F��=ܣN�s@n.b�{䖃,/hiӬ�n��ϸml��`'A&AqDl��?�WYe�-8��"LuL�<�ONN�#]d
A�(���ZL?�޳��nܸh��L����'	�[���T��! f���?<>>��V��	� -�J~��~mww��$)dΒ�W�E���Җ$�ɣ��1�}X��,��Y��~�<x�8D�����������r�ܻqД�vyǀK��o�Cʹ�	��.07���h�-�8@��wצ��761.�7'T�s{� �:좕�Z�ځ��Ev�A-���A988�ޛ�/wjJ^��=���
R�,h'�-P� cd(���,Np!�������J�_���&TPt���p����+�B������Udk�%>�";���m�d���#�:і���_\Z�Ֆ�<Yi�!��B��&g�7�>�!*2������^�,IQ�!���A�e�9�e ������ډH�Bc.�Ұ{����.���O'�����O�w��_5�|�=���mb�
9����}�\���y�r�H��Ԟ�[�P�uP���t�n���B31q��5��O3��i���hvMI)���e|ՒF�_�)�)d�v�� �!��;���6nŠן��9�n��ϾX鳻�G{�ge�B��կ����������������w�>x�`y����õk���<�?}�O����b��??,M�̋�AǬ��!˶X���HA����}���ý��yB°��k�J����?c������Rڬ,iͣ�(ɭ��U��K��I��E�Z�Mq�@���n�t������4�lN �0�%���ܠQV�q�d�� T�%���@����"
B���1���i:g�Fd�La���CF�V�>��t��M�E������ˣ�l�t��L�y���"Ȫ0\��$��tg��{�����wdW:�[E.�0�b>�$���Jg���SD�B�����8��U(6��%��:��_z饧�z�� `�w�}H�V��7o�������!�#���_���_��=����G@5s�x�S���?��O^y����w���R;�Ѭ��1#��c�Yj�� m�'Mg)�;a|/���&�������6Y��P! �`e0\F:���K77�+���=�z��;U���$����.ய���IbT���[ߙ�����;�@��V�@=�IX��)���2 pF%�j:�r(�*���}j��w��ν�6�|��t���?c?�F}�\�0�n<}����7��mr�q�i�~��kˣ�� �^Ouлo��[��6|jc����Z/�ƌQ��i��-����zQ��@Ey0��"���ozn��ݽ"Q��Ŋn��4X�}�!e�	3��jUl���3�H�c] gv��H_Į���j���ҖAi�V[����6��EC�����3��NdNZjtثh�L]'G��q���@S�RѲ���GUل=��*7�!�X����Ft�6���|R�4<��}�N�y�+7O�4��g�7L5�5���o+���h>��"0
��(^H�:o��Z�?}���l>Wmܫ���x�zR�O}"�/�����������	�����=��`0�s�ȅ����=�~%,3�¡�zt���?�<H����0��x'��H̻ S���z �((��k����g�}��ɣ�}�{�+�/��KQd��$f��qgg����Cɮ��@�-��-WJ����;�q��t��k�p�@�{!Q���e�J�}1M���?E@�#�G���� �ճ%E�ho���/���:�YL�%2�+#�S�t�+?�!��(����X掱Z`�[�ٴ������v �6H҂`?|!��uQa��n�6}-ƴ�����+�)�hg#��)��!��b;	\����
�[x�0l��J�lt��4��+�}�K�lv�Ν��~�mk �NN�Y�(��� UBk���@�9��Y��e�`;��'�.~R+bj�d8Č ��uUi�(1^~ewǣ�#�3�-/#N�d����֖�� ��d8]�8A�p�,x���p��jS<��9��OEN�KRmI����1#�"s .��~o�ղ9��YB8:���cB�qb�<�p���%{��k����O��B9�C4n	�=@��T�u`�W�mY��W�)pz��[���h4c�Dlx�A�������cQP�VH�g�Q�B.��^[�Җ_��X�-my���V���^V p�Ir)PR�(�̓�r���E1 9�L$0�eA�U��)D�� ^������w��v[ln�A���^�"�{��L�P!Ƙ�%d2��K�5�%��42M��f�sDM��c��γD\�����E4p�a}�CVr��z���Y�8�}~.���jbM����*w/�c��|��_�y{�s&Q): l�]K:B��RWHqm* ���NN��޵%�����O}��t�����o��1H��Q4X%҂@��Ƌ�o��[����޽�{|����dv��2�,ǧ�����gÕ�yq�d�t{zbًGϿ�ʧ:Y���C-6���������!\�3�	0Y˂�-M���������k�I��[�t���*�",zR�E���<[,"��ݾ�c���\zQ��p�0�C����m0j��Xt����ޛ=I��u����w��#2r_*�JU*�J%	!��hԚZ�``�m����y���`lx�10�X̠����@!4�Kk�TKV��F��������{O܈,��R�������s�v������g����>�I:�&�<@�1s ����J�.`�bEd_��iz���A��c_�t��r[�w�B��S����ֶ��7���{߻z�<�5�
�&Z�i�#����я~4����Gc�K_6w��0-N�+����o���Qb�T���pww.h������Il�{�G`HWVV�A9�����ϧ�|���3��������7n|��߅���o�|��_�����������nJ·�I�t[6!p΀�X��lD ������|N�l��mom9�m�F���)�W]QI�d�6Fg�V�S���ZQ�VO���B�?���e����o>���y��7}�_�}�z懒�lJ�}Q��)l7!
�*�uq��6F��k�]d�0"@��j��z��իW7{��A���J��l)c����xr��ڪz� ��g�¶2����p-�Ŧ*�G%0�tVu�]kW�0#�]E��9��d���^��b��?EtZ�Dt��С�f���%Ic��u5X储fm`a�T����;�}�ߏN�<�]s�ʴ���M��Y@Sq��7Z��M��Q2ME��*�4�.W2�c4˨5+��C�֚�Y�QK	kiHp�5�j��"�)��!أ��I��aKJ��J%RB�,�򯖩M��"�	Q���g�Y�*qD���7>��hJ�-������#Pv5�W�a��"ۚf��UY��d)��uۯʬ1-��y0Jl�d����:Y*�\�ć����.^ȫ�c, �u+�h�$U��% Q��=v�4\	���DO>����}�t<�3���1�����u��O��O\�~}w{���s�ڕ�E�;�l��Z�;�3ѱ��Wo�����Y6��3���!����f$�΃�ZU��V�%�3Ly�EB�D�qf[ſr��O){�[Gnʢ����21l���假�[����>%%�(�7<��S	��Y��3;�j~ɡ��Fs,�}B�MFFl�m`����}�؆!`g7#��ɓ�c���B?`�@[p��Ѫq�����Si��X��61��}.cҏ���o4�Ŝ0
�!����sd�^�?0Ѩ����e�-��x�W`u�ʁf 2���Q��pk�)�k��z`�Ba
N����D�,��]��A�`�vn\�$�c�I�?ا��`$�ՠq1z0b�`����P���,p���������V]�ܢ#�#F� NЉ�*�B ֣E��v��9�;,mϽ�[�Č�HZ&N�L�f�x|L��c�eA*��	�YNf���?�iF��oR\�*�w�?"?h&'a�B~� gibz);>pzcy�i�U���>�=�a���m!��0�}��b_-�����s���=+�2+?f�a�Y���+``d�!���պ���,0%3�OR�?$C��Ը�QU�u��Ԧ�_C?D�v�7=��3	�~��0�m�-���>�<-`�P�΄�|6
��QL���r�x��o��R�+�Z�&8dɜ�&N����H}%恍c�Ʊ�G�l(+��8�B$�^<��K� ]i��,!=F&yijL�,�}����3�7�ХB�����2]Y�8ouF
c�
�57G�X��?��[��^<M��l��]?��~ln~�����F�6�_|�һ�����˿|�{����~���zO�k��+W��wN�=�d�ƭ�q�:���Pk������:q�̅�(�����[���L�[�6�k����#p�bgL
��ศ�©U9���4/��M�P/��B���Ҹ�"�m�b�i�v��aP�d0O���R�8M�����JY�L`�m�,E�'��h��j0�u�m�棉
��J�g��8yF=�$
�6��D��8Kw�w��O%�@6�/�}<�#�*�	6��� 3�<u,ha.|��m;��Aǃ$����� S ~2�0��{��8Trc�Z8�a<�F�g�/�3�����|���X���I$A� �@J��zaa �g?�Yx�{%KKK��+N�������!^Yz��L}��W��e�����A8]]]�ha� �A��z��o޼������b�r�J 6VuG��Q���� O��v�{�w�w��AX֥�/��������w��i{˿�_�N��ɳБx2���3�+��h:���U�Ф'O���޾���P~4�HE�!��� ���`�DYA�8�=6�`Yֲ���J�`'2�vG�[�;���fw76.��$YL�F����ު���#d��,��j�Xe9C� �6.��7aF�G�4�B����Ҷ��܎aY���(��u+�T�I�,�E�O@��s�����zL1���Y����RƆ���ӹ^�ERuk"��H�%&��*�+�sTyE�9�'FIW�*�cx�3ae�����Q� LuVfeV~p�a�Y����x���F�qƠ��'�e��b�,�zN�'�0�ɗ��0��!��\����*T���!R+���3x|mq�u W@U?��e�L��c�#����8�C��YJa�m_���l��OT	#���,eyʥխ!dI�8�=�n��:%p���Tˑa9,�;�XIf�<>�����(�X^48��]?Ln߾]�%�`��-Q�o�EV����{�R�eU���|��ꩧ�$=s�!P/n8<���}�Q0a���yDٴ��3u��}�z�����s�>�8�LMD�j�6Q�c�/`�)���ʒ%DQBà�|���D流������*I�;Q��J��SGh��7<�,��:������D�ـ��L��C�uN�2�Iwg���܁E>�����P��KP�ŀ0z1d���t5ͭ{��
�̩S��_��}�v�P"�Sx5cIb�?DJ*&�؝�Y�)d�aZ.�\j��QB�X3(��2_p%�h��'�d�����>�"�?���ӧa�a�.<��t
w�+��Πa��8� C�D��`7c$� ��e,��Oy���azPR��͈FF#�:�F�uF��YƜ��(��ƍF��֖�h�;:�$�b2e�����xLU\�� I9�T�b����c�YX��������*$V�`�U�0h ��y��g��a�}��B�z�y�܌�C�^��ZI���GY93�C3$� 	���IRd�l�E���&��=f��s��'Obn $��>�Z�3��lo��q�w^oS3jkVf��/3�5+��E�x~��YB�͌jL����<�X)[R�=iaE	�$�B{��7<	�IV=��U6���3%X<n���hg8n,Ƃ��EJ�]T{ZXBY����q�j0��4=C��S�O�����jG���x�ʤ�橌����@uX�BSmZL���<��@N�+��%��%4�6Oqʚu�Y�b�����q9G�p+2����
�زCN���VF�%�z�T�CSU
mRl�(�v��݈BRd��R$�#�ޱ���`�q�������-�
TO1}��[l5 �Z�n��9����/}�KǏ��y5��Yb�q��W6�;��kûwnݝ�[�E�0�� 6�իW{C0\��Q��I��bV1���I�����I�岩g���|��J���P&������a���(�]� ۓ��jS��|�.,,�~���z�%F�A��ىH/ۗ�Qu�&���	�$u��DO��a�k8�r�r'�>��	�C>b��~�y�������,
��2�-���"�Ed�D A������ʍk��0rmg2e*�T{���v�g_	�`��ϵ?���|Vk�(���!CM�~�#�(�	�G�(�0���b�>xj`�yǎc1w Q���Z�V��������ͥ���P ��.���+p%L/1i9�iR$-ob�g������ ��#���-���9=�˕gV�Gl ���c��5�f���z��Q`c�~4�ʊ兖�O���h<uM;��;��P��<�rW�$�0ӛt,	�4� ��0��P$��FR�2a��I~�ת�V��l��L� {���X�N���������n�j���2-	��9l�唼ۍ�h8���6��� �Q�E�UǛ��#maWLi��iDB������֓��S'q\��{`�R���@�Rjːxe��J�E�30�i�1��`,�]j�Qt�Ӭ�� ؆�.�N�J�]a!��E'&H*iZ���NEb�XQ��䒰�vPS�n�ʬ���֚�Yy��J�=��'����/%Y��Ѡ&�W�sB���)}M�:E�D"�_��h������wT��AB��{h�N����9++���[>���
bĥ9��a���J9�Br�x,]�-ԇ��4�}���� �Y��h/�8r%e���%��C��d��F�W��!��ы��6�@��=�ڿ��� %FE7RK�a�T��K�S�W��+u�s��$�%#e�8Ũt6�����Νk�X�&ݟ�8���/^���g���������-�i<����K������W�:��0דW��_� +�������o��ҧS����ַ>��3/ݸB�4W� �*l�E1��^��I� -FFS���Ӱ��8D>S̀�K�tQ/[e�fj��S:���b�������z�GL���W�.���`P�{m�(��YФ��U�G5�M��9��3���c���e�P�*=i�'�������1-��M@M�Nə������g�ݝ�`�������ޮ�`���?����������>�β�KKK�(eiP��l��?t0���9&je��u��l���:Lo�?��4�ዿ�;��ӑ��o{��Xv�ƍ��onn��/�"�"`0~�� ���?��?�7_}�U���>�1 l_��WH�#�`	A�`�/]��<��&J')��	�9����&���
Q�ǩ�^9�O�N�P���p�Bw`��˿��oy
:���OC��W������z/L4L��~�%"��PA�+ �����-��G�q��I<��1^+���r-h�[��3g�$Ҁ�*�&�<�:�R�_�������g	D+n���z�@O�k��"I~�K_��n�ko~nA�W�.�̿��o_X��.�]��*�8u~
��:Q�&�%3\D���rb
fS��LI�� +	)�b����qM��(���(
^���8���f��9���[5�T&�~x6!)�Ҵ�J�ʬ�w*3�5+����(镫$��@t�X~�"��s�DZ �b��\�rɗt�6�3R�sI��y��X��>���(~�:�p'@���g-��o'��}�R�,1|B$�;w�����Ɋ��F��@ԐC
�GP�*�jFK�:�PK׎��veh�K���J{%K^�l��.d�����2Wi�([��$hp(��ܽ���.kK�!�=Э2��6����U�d���ݳB�� �t"�Ci4܊��q�l�{����l2�/,V�n��(���К��n]�թv~���:�rܫW�F�6�2C�7���`�gaZi9�8��[���W�p��Yn�g~��U±�4��$0��,��X��LҘ�]�-�">��^�-�`E5A��$	w�`�(<D ,;�5�@\��"�
w�m�3�� df�2�e�ab��m�Uo�e����۵Ķ�O�?�η�� �K/�|�F�Z�ʆ�i�)�I0��V�GŊr+;H)���aa-zj�Q��m�W���;��DULu��Ò����|��u�U��8x��ŵ�5��n�ƴœh�?�,oԛ�����0P*3LeB�L�bCd�*�
y��xZ�ذ��@8��[s�x��qY�X��3a�a4 �i�[�E��ԧ�߿Ϻ ����������L� c�`F���A���;�>z�~�=��>K��={ ����{�<�ك��]�,����6hvp2ovP���0i�xx���\���4{~i�Dpb��\s�䉵�c!�TC��l��vS�P!�X���H� �8�mt��`�L���"?�i�^���n7[KKV�6�B��2��#kn~0[eq^�*�4�`�4-?IaWR\�'µ�N��³�6U�v�A���°�z�ڵk��v`��uܷ$�SvZ��c�c:u�*�i'5���RR0�BU�`�&�+A�R�ٴ�"�?����R3E��@-�4�a(�ӥM�d_�Z�>�h4�4I����r��*���0A���O��_�+ƭذl���gi�OJ�y�H
3�?(G����ʬ|�2�Z�2+Qr�WJ�m2� Re�|�`Dَ/����G����%%W�� �c �#�3>�t��]�Du$y���)*�}�4�So�e>d�Q�@0�n	�۔��ʝ�â�� �7u��ޠ�e8d���,�,n�9+��`0��j+W��*k*p����'K�|U&Y��h���Q��ae<mPFIבb�r8m㤴`�-��w��·yK����[;��O5�s�w�ޱcǮoo��?�������*\��饗�iv�t���``s�����ws�`���<X�`&���o~��_���w�3�BU�0�P�}��8h�A��'�q!�&�`�Q�Qd`��$�;��N?B��V���������#����y.���?_ÜB�5����%;�����Ν;H&��3TQv��\ZZ���_�[@U@���RP�c:</�7O��B2z�0��u+��6��}�߼ݺ
�`q��l���� �$W���zjnu���G�G�o��%*X��`"�i��|��կ\���"�֐H�.�Ia���?D�Գ3'<��-,,p�+�~�#�a������O���M�s0#�u��݂)��~�k_T�|&���c��7777ϝ;�:��w�w��������e0,�?�<���7oB�s�/��#�ظ���� \��e3�=����?�1챪$ga��$������������[[��'�)�)t
���;P��Y�^8�S�Lm����i���,��0���t��ӟ�4����]���y���������?�*��d	�u�-l6�hR���M���>���/_��g?[k�i�3�a��G�א�ӻ�������'Ϭ������h�������8�m��8�g��J�#˕*q�R>Fx����2�:8M�l�l�BB���88�3 +d�l⩒�3B��Gq/��]�?�ך�Y��TfXkVf�!
�?�~�9�i���('��/V,�LH<c�y�%%E��P��()��,&+�j�MV���^w�U��F̂d�a�q�(	m�y��L�Wm�w��!��@�6��D���H���.��B�C.K>��r%�?Xʸ�A�f>؝�?䡠zSxԔ��&]�T�&m������,w�QVR -����\<�Đ��W�,�8���珒�pܮ�m%/�>�R
'���p��+��p\�݅�:X���j���^�w�]�Z�|8S��kW1Rh�i)���[.>���Xoũ
�c�g���[�v7�k�~ �TH�[H��i��h��	���)��u,˱�T��$���4j��`�������m��	��;ݽ~���Y���x��Xn��$�a��Vm���b��gQ8���&ӊh{���ޮ�zґ��Źp�М���c&��M:� �R�{�B��PEz+�� {T��Y�Sh��H㌦{0J~�> �JuފR:�Ѱ�߭��Z�;{�/o�U�*�(R���j
/B�2���ݖ�����Z�u��1`�$¤_`z�8U���t�3vgL��\<�`��Y	!�@�E�����l��ߺu@���1��gw>I��P	��j�~�;�N�;`Z���2�XfB�1�C��$$Jct�E:%��q�i���w�2E����Z���GY_[�q��4��*�8�`���1<kN��1mf�� kA=�a����)�<���a(����R��OC�ߗ�[�{�&n_�<��܂��f*��U)T�plX1I�ʵ	��6OG�QoTP#�̭{w_z�����\gѫ72�6҆�� ��H��7�mLǾ[wMۊi���w��&~� ��.b�7B��J�-Ǥ-%�A�Of�0]�W|FCy�L� P)�E�n`~oi������N�R�e�|��/���~DѬWh���(e�ޔ������ʬ<L�a�Y���+������_��| ��g=fu,F5X����&>��H��s{_�9��9�xP�L��3�&���9A��E#1lo|x���N�CO��)uH��AX>�7��7��T�(D.�_n�4R���2& Ny{-�Y����##�;����X�V3�'�-�o�f +������H�|[�;[[`+���y�����l`���կ~uxg�����Skgg�1-������!�%����ŉ��*x�����WVV����޾��#�7�Xs�!"4"a\�U씴�0��k����x�
�����߸s��"
��v��$��_�c-T��7������п��`k��=����*� [X���.sK�A7��>}���j��l ��裏B���)�;�����=?����'��p�4R�����؞�����H�!��b�����``�ӟ�4 ��^z	�����"~�+{=d0j�XqF�J��Uy=�{�F�� ���h5�<둅���J	���.hc�;w��L�`B�
�FL���;%�2�F�J�2v� !��c�lkkFuoo�ӯ�k��`�:���V9�t3�L�"�,:��cd� k�pq��Q�ԯ\�r���Wn\�o�L�c�`=���_k���c�q��ɪ!����k�)�����:�
.�����Q����۞���j����}z�я~j�&��O�˞}8�NF��'+��" ������}�k�}��.�>�/
��JK�V��w_~��G��{�BK���o���+P���rBb�*E�i��oh��E�ɝ>�R���{ �Ad�:x\��aIv�&^���>�ЇT��sHG7+�2B�ʬ�ʏSfXkVf�
�ڹi�	��CT
4�?��O���'�32�1�֑취e�{*A���v�g�T?2��"g]��C��,�`��L�N�zD�O1���2�����Gx*Q .]�Ɓ���2J�G� �7���n�|=�MׯJ�a�o�&4�pX$({��������J�Y5�;Rsn��$����������ea����(9-����b�(!7�� 0�[3�i��rlI��g�"��I��u�m5N���:�f�X��f'M%�&�y�,a� ok�;w7�L4����ۗ��A���\0+�%5����
��E�Y���lB�:���{�dXGiDaC �^��<?�0 �7����n�;kK�g���]�l�߻��kM�~ڂ+S����`����:u����
���j̵Q�o���~5�ά-{��i��0�30�Q�X"ƙ �+	N���ڷLm�y���*��ȩ?�,5��J��� �UGQ
��i=�����m���Q��ұ<�D���l����q��B�r�g2
������ᅮr����F\��
#n��x��x>O!r����Ch+�&@5�k�ڍ���0�p���ިA[jN��i�\���^{66����� :� � ���$� ��dȠ��+: h�&������D�h��	"8��������ep�S�צ�QF9�$
}a��p(�q��@�(�)�R�r2�TB�1������!a��h -�n^���K��յ�4��n_�ve�O��uF;��S^iʨz����q�".�����Le�-���ކ���"�Zi�D��jUtǅ����U�5��8��$�ﻶg�!mA�l�*�3����~�E����y��q&>؇t�B���`N>Ï�$U(#S(�#�ǘ,ڲ�&�E���Ή��j ������7"�FJ���zΤU'E&m�yɉxC�ʬ��QfXkVf���`d.�#q�5�:QK���4_r�0�JTLn�*%��o�F����M園L����P�(36�����CE���<�(��#��,b���]�Q[���=��߯y:z�q��ў�(�M#`�c�@H�2�: ���@a�+����,Uq�|0q%��{�(Z� >N�� ���ܜ^��,��ʊ�I<ػ`s��DՄ�c~�4��Ɏ���q��Ѳ�s2��a��#���mll�ə3g��D֥?�d$̂�&�K��8أ�z�*ޗ�V�T���Ȯv~;w�ܝ��n���0����x��g���w8e��b�-m�x��`pow>�/��_���^���\��o|��K��~ky~��1Q��QVv 񒏿�������"��#�j��U�u ������{��E�5�֯���nݺ��[0���жQ�� 	CB��:�X���΁z�y��}��~��$�I��&rH$�ޙ��cǎ�qN�@��9���=	�"\��	�]�z�MgiZ��
�Y`�6���3� ��Y�l���K�G|AUp���-hL',f/DV%��A%��`&E���;���L�+lV(�@����e���4�𢶽���];��0��}鍅'.1=k��
W��Y��5屰m�
Mف�GP��h-oPn�/����`4T$j�y�g�x/*�˜UVda�e 5�(��kmmʹ*/��b�H+^� �	4)��_�~�G0�m<�19y�$�������V�tE��AD��v�� �U��d�&��́�(+��2_l��be[*mb�gA!��^(l�@j��Y��Y���k�ʬ�~)[���=�]�0a�ԔY�%�T�Kdb� 6�	�*���S��F�$��;��#����y^0��H	�Y��\����|n1	P38OW�t����0|���6�4"#Ł?�B�9��(�S�ME�)�,5���\L�}�sJY033��#6E�"�(
#�Z�e��p3�$^� ��"��0���i����ů�6;�B�5I�=�0���a�mK�>L�c�,�Q�LŶ�~l�6� Ԭ`Ι�c[�,r1��,I-N��q�>v�( ͱ�I	��=/��\�_�o'��$�u��1l�V�L>]���Q��t<�;�A5.��u��`4�9^�r����=Q���n�t͎S�'&��0�f8��ҬV�V�s�N4�,v�k���8�������VV:�`�z��'��L)j��\��޸���LD�P�ЇU�o�8�íT+H�g>�O��~�W��$��po	4a��g�������j`������O?q�N�f%=}���w��Ν{�z���B>��S;�~<��[}�$�����
��?�5Wv\S��Zq�Q��i��ڔ�BU�,��T��^m�όh�v'������ח1C��W���B��~Q|�5���j'8|��p�=w����\zܡ|���Qτ�㋫�M'-S��U{]�4��p�,��mdfݩWL0ݫ����H"�*�6�5��Y���l5�!�� `�5� ��`������v�ƍ��%�`΋���^��.\�`Z��^Tĉ=��Ҵ� �Zp�ݭ��o�F�u��{ \��\e6�%r8��1����x'��a�,�u0���a����0٣��4��0U���'�����&�hjb��LFA4Yh��(g����\���<����+K�Zm�� o�*�q����T.�o�lg����0�p��SY�J�-+��gU&�(u�|�'�
������a(c|�º�|�/Ћ����a�13�#1�m�ęz�ڞ�ìeY
$t�2�����N��œ/���;�~_��c��#Ø[��+�?���d'q|j�dͬ������h�3Oِ� ��q���2C "EN�<�4���ē2pb�e	{��F�J�?G.*E�B؋���Cڱ�TS&�f�S���-S��g◓,52Vˀk�j�����p�?��S�j3´�)���+I���=+��?r�a�Y���(��唅 ��<'	9�p8���1
�<���-�"�;��88�-�5��7 `� �HҜ��/K~w������Cex�h40>L��BK�(�������#�I*Y8
ʢ�GEI�O)�� e��A��t���:��1`Kɯ2�?(�x�&�AS���>W	eԥx�H_�߂+����^��9ɣ��]�֊d��'70,�^ӱ:�ZZ���i��00�f����UXx�(p���x�����4�L��2�L˛�{Z�X���F�d�`?���j��kb�mh6��}Xb���|����B��ݻi�e!;@  ^�[ժ��/|a��:�Sow�7�[�^xygg���&��xH���]1E(�`�vw�v�/<-�P��r���/6N��t����|�#/��]Θ���p{���|�'���<��:)y]�G�<�U%"all�p�C�I������~h�Ѥ�L<�`���dee�Cj��Ц	%��9�T�����+W2�6ǡ�̘p8������'��Ƙ�0Dw0��g4����֌�BЋz�
�H(kV����
Qdr:���m�8q��$i���	?P0b��߇)�q������s��A%P9��x�
��<L�,T:�N�et��T�<��Q��m�C�W�����,f��Q:����9��-Z�MPWsuiaee����_���6|���ӗ/_����5z�*�`�C�#�<V��c�uN��&ޚ�Ѡ/0����|���S��׮][X�Ch?�LXL�C�x?����M�j���5�ݸCGE���)#t�h<��F�]�S~�x����SP��� ����Ac:���{�5�n�q�U��#'�{T�.����Md��(,N��2��
oe::W��|�ez[V�fO~���V����z1+�2+SfXkVf�!
��(%(0=#��j�۟����cT��H4L��>D��4T�G�I�!"X�P���Ha�׶�T�a�9"FJe��x���LG�H�����`F��u{����}�"��i�A�Q������d�v���,b��r��B��1g�ťT����|gHG�1dy��J��QR�'q�cUni��8h�Q[B��M����L���TjՐ$S�fz,ȃS�qD�c����Y	�N�Q_Q�Y���I �iH\!��8�l'��t �>��%���VF��҄/˘@�c6�Wb�6�-��TB`��/.�M?��{=ǜ�U��.�}��G_ٸX�;���@h�:�M{������θ'U�����۹y����5@2U�l�Zص��`���y������ٸ9ox2`���������IXL�=��3�Ея(3����C= %���-0ř�cb���.����F�5ڕj�D]u!+s�jbM`���o�^���;/���!d��x1��KX�uϛ���I���{�-SNUR��~L~t��UR�����`��abb�#A��z"x���O��ڵ0Q�P�jc�}� ����w�ԩ.h��,{����
-`�R�j����� 8
���۷�ss�m��K� WܺuZ�)��v0��(�jgXQ �[���2����6�:��J����m��!\���d+����L�uT��,<)�QSdi�<�oa��f���n�v��I�G
U�3��k�q=2Ia5�����3�!}�N��}�"1�N�;s�}�o���͛���� �����_|�#?�?�xN�I8�~�G��i%Q���Xk��^�T�_�z *\�O7���������Pe�Q�Z ����nW/4�b@e�����x~��_s]c}m��G4�~�+$N���9�l�;�̷)�^D)�V�Z����/]�,�w�w�@�I���o�a1+�2+?F�a�Y���(jC�Q�P�"���?N2We�.���'�PQV�����@4��WxI)
�Q�U��)'��'�8��QF���F�&p�K�J6���w��I�����O[��z���4RO��4�1
MB����o��ܩb~�����-W�*�����E�� 0��7�Ǉ?��GNDĆ�k����{���5�SΟS�#_w*y�H�X�< ؚ�M*���d�E���G�kV��k�������I-p�K�QB�+`\>��3�4Z__��'��F���Z0U��7<�W��@T�t�&^[��6�M�Ô���}�gމ�	M�O�>�2�a��O,<��o�TB{�4��?�C�eH��H���h' h�3g�S?��3�%I�T���pFfoo0O/ G�qK*�i�M�ԙN1Tl!���d�ٳg}�8�*]v38ۼ��x3e����9�s�/�Ns�ݻ�~H<�G
�u����J�0>��,�;y�$���W^8â���ؑӦ��X�����p�w���P��"���Nf{8F�>����$s�sTow����R#�.v*x�Uq)2��d4��v��B*7+(y������qq�=RѤdb>+��F=�z��1�d�@���[�;+H��4���x�A2d�G�y������7�$5�a�0&��-Qv�C8?ϝ�������JP7��]Y��s1+�0���虅������v�9cYE��
���ǫVq �f#9�L�O�,�,�o� $QY�m0;���CA�l���Z�Z�w`�f�kVf�!�k�ʬ<D�F>z��/(��>��^v��"NY��M����(�OJF1��Yth���R2<����p�&�x��bL��?�c<0�)�F}0'�2��s������Ȫ�^yG�ӿ�XTMc�d��Mi)e�ć�|�d������47	c�\&�P�#g���d��4-m�(qH?C�T���2��PS�D�V���6�4�>t�L����`nD�ĭaDH�hd�B�ˏ#:,
�C�0��@�0��AH��/�Y��<X�͒I0�]�E����2�R�����tp�Z���Q�$��4E}�7m�h��@WT c��jؖi%2�L�QA��,	]��qE��q6m����`+[B/�
�s�ݮQ�XG6��4��F�n?�;���l�+�Z�?4,g����~�������  T]�ꮅ6}�nA<��C7w��Sg��27Wm�cZ��)����d��gO\��k�`����`����P�&!c+
`<F�`�PF�lOd��(\�z(�?M�n��2�,���=�q$fC�1N��1�uK����d�Ú:y�4��\m���L!�@���$qG9T�����SXq�=�� ��-Y;v�����ˑ4 ��C雀�0�ǐ��Ԛ��Е�´`�2`*a��l۫��
������0d'|/C�3}���[�2yE��(���[ �۵:8R���u�Je�B ����ͻ�7�3ݤ��Pec��~4M�*���]�LiF�u�}ā��� O]o�ۮ5a�w���;���} =ʃ���g�>�RJIމ�zמȦqh�3��`���팾���3��;�[�T"c0��Lf����')�D��9�׫Q��Rp����꿋l��h�����I9)N
��4KY�G�z�)oJ�¿G�,�� {
*�	��o�P��aU8�ʬ��Ö֚�Yy�r`r��jV�|��a���y)�|>�<�4��-i��܎�.5'���@�h���s�� !���vG^|��Bf�(_ 
�<��S�M.��R�M���<�FI�P7�<b�"�M|~�Q.�ޛ҈e�|Fw�a)�#}Ɉa
B�͢8BV�4ǂH<�g� �B���R��7c�)ȷP�^0EƳV^-��� ��1�j2����z(6^���80ǩ!�&ɓ���Ձ�ǉս*�/��=\�-�0T�����A������.̀R�-I���h��F?B��L5���t:����EM
  �r<@%��j5ԫؿ������ٗ����3U��������P-�w�����7�����
�����Z�1�f��aP�>�!�����ӧO��RxЌ��_�}������З�:���]��\y��T� kQ�N.��j��/\� X�ʕ+��yM2��H-v��͆KP�&m���h4��M������'O���o�t�޽���߃�ߚ��Ë������O>�d�����Z�����=�T	�+�&;�]`$�_gΜaa���- rPU�݆	���?��ԧ>u��uf��J����+���w������1B�|��1MZi*DvKF��0���H&�V#���!zYRQ�L�(G��R��*X��"����`J�k�E��&>Aq���GY���ϵ�y�J�?���������0,0��^��ٳ�n݂��#�f�cSs��Z���VG�a����O��=�dX��JY�M:-�$a����(Y�NL7纟��'����Ν��Nsa�8�-�T%^K���ʻ�(��<���aMy�-������ݎ���}E�x�Y���-3�5+��0E���/���c���PZ����g��fH�p��E��$6��r��)�<a�t���"�n�Q[l��G��[h��C��fI�ƱȢ3����$>��W�����p���At[��0����4&��`�+�2��}npV����"WUٗO����S�ױo���#��`q�����j����+��!�ԇʲ`�x��#��*�G��>�yN�-Q�`>��i�P������+�/%L=��yr�2�$��@�MX�I�h-!!fP�ҽTD�Z����TEFՅ��6�f�����#4�6��gy�zzgA��p�{`L�|]=��p߰��6�w��K`4/�7����Z��Þ-3Kd�VD	Fd�:��O����b��!f�k�#C97�,�R����+�(�++u�cg�1??�Ykl����M0����,�s��q��	T���P�;�4H�t~yz
w�s,�i�iإX�m5a �VDjxճ���h`cYi�i�L*��S����ĠL3��cC��	mL~e��	�;mt��� �G{yie�Oa��Vj�W���#�>��~��ݻ7/_���+31a���6l!�O8?/t���!J!��}�P�D) � �������?�]�W ނ ���}�l�ق�y��ga����|���(D�t�#I��4l�4E�@���<�?��8WE?�����x��ra!Qf˜n�H��� Hꖗڪ������%�V?~�d��`>�j�������.��� �@Q� �a���t��][B����<$���f�J���{�KVl��Լ
���`�0M���7Zm�����.�p/)c>va)��F"�#V E�W�p*q"�����P(t�)�4 1X��lX���iV�[������z,��BPz��3 }���������x�MUלѯ
�>�m穷��~�5+��c�֚�Yy��ԡ_,��qQ)?	[آ�(�����-^֮ȯ���w�QV� /�aw�4�3��i��SL������Ζ9Uj���2�>�!��]��G��X����1Fҿ�嚩��>}[Iޒ�Ț��33�+Gh�2v��A0(L+�d)��8,ad�2�Ҧ�fOܿ�3�3(�N��q,Y�p�`10հ���b�`
�X��׵�
����9���~!��6��sd*��)DY�$�=����j� 7ܹs�lί��$�P����Nބw│��I�'�Uٞ�@Y� 	����a� �V>X���b��2��M�}�����p|�-oy���:��U�. 0���GCN�d�b� ��z�[�xꩧ�x��7n��_��իW}?��������c���ٳ��+�r�ҥ���C�	�_��r o�Vh�7��=u��H��w�`I%��Y#���c�a�4V�H�t��)�a�����5�'.'�\Y]]9q����������N�`(��Moz�����%���^_�߯z@,~�9���n݂��:w�ܓO>	�<�  ��IDAT�����w�k+++���'666��_����߇��������Ǐ��e+�}����DoJ��b����L��%�c�(��#0Zo����&����9�ø&@�P�v���w�k�Աg�}V8��=�3tt{�۷66`�lmM���m�W�q
����-�]�x񢪵�˯���G>�AhR45�޽ ��ba̞���Эv��'�'��k�k�]:O�8��c�2b'�T�D�"w���'�߇���:s�Y�T�f��A�	��0�����i�Oy���� �S�Nz�/u�=Y����d���[2��H�P=�����ʬ�ʏ\fXkVf�-h,�@�=��ȵF[��ɹGъ%�ʓB���aR�q�A("U�0l
)�#������):�4��Է�kY䜩ǅ9.�RS�4��S��5��a[�ʳ���(	��ԃ�vx;R�Q�m&2����>rl
��U��J����f��M�،��D�A��<8!+R�j������}�ޠ��R]S�BK�	q�R������Ԗ,�U�~�J��U���[`	���DIC�n�FS0Q���KW�T%��`�XH� ���g!s��R��j3`݁��b���I��K��82*C����Ix�u��Z���x#�cLXN]i6�?�U��Tuh=���ɨV�(L�%u�Tx�&S��"X�`h:8b�%�^�v�(Nx�.�;V�|�
Ȋ-N�qC? l
85Bײ�L���n4�Z-�A��x�:~K�Ks�s����2�\|~
T�"�%���-�-?{bgw���{��w�����4��D����\?�~�g~�6��-hj:�Lff$( 
h"�#L�kE��GiR����cgq0�W�q25Lx��H�	<�0����Ja�xP�Ԁ�zຘ)\��2�
�>��G/�� l�E ��
�u@4�z1�C~�qs�zT[o6��Q�<:=�`���y�����*���z�37�����"S���ɓ�6!���4k4[0_��~��j�j�V���1g)F|��ͤ?��%=����W^4����>��[C�;Ï|��(�٨���a�t�ԝЛΟ�/�\L��;c����P�|�u�ԩ��ݡ7��;������7P��������+7�]y����U �Ǐ����6��奥��0�(4���ZxȒ$�~m������ jq��z�
K/If�1D
;{�b;� :������4��~M ��p��dN)V=t\���@��G�d��)�-9�$)�b1����9��t@�N_�RUB�b�7K���0�	�p
I�!�(��Y��Y��k�ʬ<D)~��A���E)#�\�m�K��6������o�
�A0�Y��/�\�����:H������	CG��^{��&�A���=�/4�`C���g`��ND�G�|�h�BN��Z�1,���0�PfY)��\j��$�#`�h6������[k@�0O���U�ć������5�b4+��u�D	�~})q�)̉J��T�>�Ί�␦H�{](�M�e��#7�ਭA�n	�ѐ4�c4=ũ��ҙ%0Y l��� ��$C�p������j5���a]ú|���`����^h"�Dŧa�R��+W������ȏ�߿�,&b�ц��/,,<�ԛ�;���.]�5#������ ���%�`���n����p_�J\%��w���?��Bm{�]X��	⫅��;����ܧ>�)+PkN)
��X1z����giu����?~��`j���DP��kk�7���/��]^,E\�M�$*��$�AZ���Z����v��@�	�ɓVS�4�f�Imw�.qJ�+p��ת-x:������.��sss���N���O�����!`�LEP������F��9�a���c�hza1`0�XKKKp=���ڵkpG����O~��?��0��>�,~�U�i�`�_x�����}�s0)0��v�oq~����"eg{��F|^�y�=��fW�s�^��DP�{�'���g��vw���'�l~�jeb4���kgΜ�ؿ�Ї>��o|�g�N�7c�DX9��>�ܷ����K�x�ܹ�76���������������>,�q�Y�10���s�<9���$�^L�n�A�*����M�����}�N~����BK�Ї��7�� C�Y��6��fϲV�+����z��@U�(�*�ݧx���yI�VIZ�Y��^���9���t�[@45*)Z���wKbL�*h�Y��Y���k�ʬ<Dц,�K��:i�!�w��c#KUf�_���N��H�' Ȕ���h�E�+��g�^��(�
����\pJ(U��jO8Fɔ��=���Ij`�N��A'E�^��A�o�߃���4�}�,7
��+D�sS0&���%?������� ��AW	n�~�RZ��)��r�369(J)!��K��T�}�U"Y�*<��ae�$'Q-���#afr�P�b!1d6)�/�d$O��E�=D�r4�'VU���EX�������%�t'#���$vL��!jz�-Q�f��j�+�Ҋ3І�t�>o�IjK�܉S�� �؆���F!;��*7et�h͵*�/���;Ϟ;�9s�4�����J�!�cۀ���RTP]ZA��p�
	��ך�7&�ȶ�8B����}��:��,�^��(ڔ͹��Q�Eh&F�*3;C/�U7�G�c�O�����NP�Ԓ$�s':vl1��jF�p7��Ȏ����?��p�0��&1�W�/�l�`?[v6	#�6����w��R��ט
L����Xf(�$NL̓�٦�,��V�M��V���d���A�;�xo׭y���7)#��Q�����W�o���V+H\�[��������y��{�<`}y�&��F#<�h4z��[�=��oP���ŘF�W2�7�X�u��3o�/��,���^�KE��I�X���ҝ��BJ#3�DH���@�E�B�fŁM���D?¡���U�^0�*���Z;����_x�V�d�%�Ĉ��hEfv�����s�3�+ue�4����u�H����i&��8�Pjk����W�V��Vw����� 0��*Ǥ���,xZ���M+��x�$���V�!wW����-1�N��j�k��ۙk��S�����Ժ�����Um&����L�1�
�+�2��bv��#�*��L{��|!|G;f�$��`D�,<����"�,��
�[�K�[�zZDz�o��1+�2+G�k�ʬ<D�??�r���$^�,��$����4��y�O��d��$�uX�c�Ӄ){�P�I ~q���ׂ���vRa�_n}ʮ�8D��~���)�8T"dr��rr^QJ������6�V���ރ�*��9hFQ�!M-~�͜e�E�����d��*q�~�2��>a�Bw��S�N�\\	s������E�[�*Qd@.߅)�NY8I
:t�m�^�G�_���D��1M�qY��i�o��z)��@���#�R#'*�~���ت�_|��0	D��D!r>D�AU0�{����Ra���.����=�	`�L|�Q�=B�P\�j��0ed��k%�a��ܽ{�	��=�R�b�peey<RP){�$��i<��\$y�pgg�z�:����Q/���j��Ѓ����S�W>Nk)�%!�O6|e���e�q�F�]0��D���6�U��ê����)�0��m��>�n�(��z��ȳ���gͲ�'��Z���i�#a�N��{�T�������,]��	��g:tj����'�?�����W)�!OZ
��>qN�qJ�N�6Q"�%NT�����N�:��׿~��%x�j���6%n�i�ٱ`k���q�� adk���������>�doo�޽{�����[�n1��W/�$N���H���m
�c.e>�fH�s15c�h-�u���W`��\�o�>�bPZ�^ܺ����bLi._�oGE�uY
в�g-+�Ի�>���K�� ���%��X�#'kz��2+��֚�Yy��:�CifIC�V��^6)XR�h'(9E��3>E�語��)}ȴ�\CI���*���$q�r�&q�S��dĒ�Qw�5k:btS�@-�;+��N�:����t�9�dD�1<[��S��"�YI���1ʖ[	|��&��4�����J����ރ��-�
H���I�B�#t��L5`bDiȑ`&])�8��(9�\��*�s�j����:$�{�&dκ)��@��m+����k'���F�J�a�&�Hعj6lT�EG�ˆ}J1(6T��%`��I�9ZsDŵ�tLs�
)��[��:LJc��p4���.k�L�l5��c�g��v�;]���h��a&S��8A�����?�!08O�>��ſ~�׮]��5kk������ ����|�����j��5�2��#oz�7k�N���'�(8�i���>w�G�Aemի7`��ý�HF�xoz�-�7ow�ݪ!���_��I� �h�؉����`�_�P�ⵛ7�޸�T���
&��0
�u+�y����v�&i&m�DS%�
�Iچ	�����x6�	ӄ�	a����A�Cz��T� x	���N���G(�(�j���2�L=׮f5t�C�Q�V7pF�>���f�"*��x��ۉS'���/c���/��'�] s�8D9�$S�av{}@�- cl�s ��@�\�R����wvϞ=�Н��`��Z���Yѽʹ2Xt�T$i%s`q&1��ı1>Ha�7S��~K|�������4N���Ɗ�����{��R��sq�č������7�$K�����c�q��K�V[WUW�U�4f�0��A�ЃL ��Y2=`&=I�<�AH62؀dƘ�Ȥ$`غ���꦳�������y�n�����_�O��*�Ζ�tvT�w?�������/v�,�����S?�qas������h$�<h�.�m��_��׾�����@}�~�M���}��~��������۹�Q����@N�p(�iY��+��C0 �kk�,=��;�Fǜ���`���\ɽ^g{�=����?��4:=:z��ٚN�7n�888p,�V�����A":Ace��[������a+l�\OU�h������zNK�	��.�/#���"2�2�O-	�<��CxIJ�%>��V ,qײ,�Ӗ%�Z�ey�b�{���jAPu����8��]0�|����1�Q�x&
�=���D�q��E%K��z�����=�k���sX�	ׁW3����@���x-S��א<�&����3�d��n6�8���/���[2���7���4���'s�'n̴��8�.�B'��W)���Q���q�)��R�����O-Ǯ7�)�"�L#�ކiCCs��4<���8n�6�/.]Yf !D�!dpI�@���lm�X�̀��|�5 �iA NI�fY��vK#�s�A:��T��qu�0�!֢�60�wvv��܃�c���zkww7�Lᇂ�
�v���c ��	�7�6�3ʆ#YҐc��⫫`!�p�kk,�]�u�D�Þ�p�b0:::ʙN�00%��t�>�13�,�$��?᫽�7ٝ���Ik�⥙X�i�ʹːZf��R{K#+�]�>��V��fE2p?l*pN��'<�����w7��^�oO`޳����P��(��'��H?v#��$�_�H�R&��`~3�/�;?<<�D~�g�dN%숛��&�Q��z��Yf�C���!\׺ڄ֕R9�n�|fF>u�h.���Q̋/
u�)?�B&VJ�F8A=rzz
� Ia��(����&������[tΜ�����3�qנ��Fvx�M"�B�	\� �$n�B�![�Ӏ{�_�mc�,��4����o"N��ʡ��8����>�}x��]�A��N#�XFHTR�<)�L�iU�1�)�����NOl��_ie[lK�s	\��uF�T|n-˲,�S�%�Z�ey�®�}�8Ct`�#e�^��?��o,d"���!�	<�l�`��#{�p2��w?�D�a�;w��I�BBG.�`}k2��"Gӑ@���k�qa����,dZPQ-���'�GJ��;�<��'��Ԯ� `;�-2�И0	^�=o����d��'�~݅�q��*��`B�k��<��*���c���s������ uk�\�/���3j��	4]��5'U�Ī�̠��������e[�`6+;�ȴ�X�5Z�v�9���Q���u9�U%����A�`+�R_;�p�o�e���>"yϾv�؅x���
۝�����=z����9FZ���ֿ�����l_�x1\]������`I�>K���]��w�ww=��������G�]�ף�����(n5��}��%��gN]5?��ן��r�>:�6�%͌�t|��%�v����,���7[�������y�%Yn5����o_�����/��g[����?��.N
�[s<�槟}�Y�iܹs����z�մ=ߵ��`�E��m�DF�P.�U�� �
�V�����\��ڱ2a)X
��lh�@z�pER��s����(6��q���ܹ�y��8s���l:�7����&0I�Ǐol�!�M���ax2��w�ޘ�3~`�ް!�_Ж�a�+W�L2���0�U�ׇ׭�-�����A�-3I��*����^Xbl+�*�R�X[p!���Կ/,G:��$<���AN�x)M+��*1���WO[�ۑ��y�ң���f� ��l��Az{�N�znge{���'�	^f:����_��_�{Ǩ=��A�B6/�cZ��?��ұ�ƳDj�5(:�f� tÀ]a5�
��|<Π֣�^��-�U�J�?��?���?7��Zݠ��C�BG�گ�ǀ�����,t Y1;i 5�}6�`�t{8wrr���`u�ef�����k`}�c�GA�b9�����)�i"�Z
.˲��S�XkY�����V3�?�0Q�|L$qݦ�7�!�� �ux�湎"ܜ��p-J�szd�Ŷ%�l?�[@/��9Kf��o���h����[}�bWɦ��=T�π�v��bF�X>�T�����4��7�� Z|L= �<����9F\�n��崏��&��@♮��Oa�p&��!��an����bqk�'P?�Ⱥ���x��me�W���'yb\�S��e)a�?�{�n���xRb<���SR�S,�YRZ?w��`��z&m$�q���c988D�rm��˛��~{{�;?�����dU���8~��X���-�T�&�pnYֺd?+&j�cfVѥ�	7��������G��,o0�n�� lny�z�z=0�/\� Чrj��?r\>*����4-�Zx�V�T����VpS��%Ly/���L� AY�������қs��ӳ�{t$��p���:N�|H�p��dc��0~c�why����1E��
5)fLQ�(X�<Iᇬ�!n��vy
0,��)�� �^C�d0n��	eUi'|�X��iYD���b���"頞*�	�}�߂����6�b�'88WWW��E.9�:[v6�̨gB8Z�`:%����t���f�91Yя������rt�������Q#>?�æS���6�v�Q�onn����W�^��d�H�1��S�e�}h1�ˈ)�|�u��1�l8�-!��,�h��8�G$y�e��
P_s�\�ǬH?�aY�eY��k-˲<E�%<z�o�в�V.l�Z"Q�d�Ja�Q0㙁P���hQ�;�O���sOf�UH<N�vh٧���N��g�{��ny���"�EYQjw����aJDF�y�[�\�X������|O�ȳ�8�K�A��C�hh:�Lu�t��m���y_�譛��9�t��0�E�^����/������"P>��r}�*���Y��G�"RY��
`�@�� l��
d�C�EZ[�PGz%�#��#ga����m]LgQ�&po`�����(ǧ(�
�P�0*1�$�ʡx!Gr�z�ض��C�y�q]��d8t+�p�8��"Kܡ�@ߠQ.*�ܿ<�Wml#>�]���JY���n�m�B²�<���_�\
��\+��xf� ���z{���.�������"M��b;hqq:�EW�v�vw_�yR�P�hf�,��=��qa+�F�}��.>���{�:�n�o5�6<o�v߮�.=���4�����F��z��N���Ja��(:9���)о�'Q�NѾ�
'�4<?�G�����|����`�Ί���?��?�΍wo�~�=8��q��3����x�vh�1l�����+׿������?����ɟ���￟Kï�w.]��j�P���{����Znˍ�'����K�W.��%-�$�)U.�6�+
�'���
���2l���Й�bl�8n��:�:mu­�u�70��1���p�������Ǐa0��}HЅ�lֱD`�AiD���g�|��綷�d
P*�ѩ̱���
��a��M�)o6C��t��~�{�{��[pL�4�=��#��ct�KW^�s���/�������Ow�i!��AZ)��H��JR'˓b+D�>��a�$���Ԭ��8�	�ѳ�b��r����u���h9�����?�����N'Pm{��n㙵��������o|��wo7�v{=Jb�)��Qr>��ٟ�)���+��^����~�+_�O~�?�v�Q�*L:Z�Ϥ�>��O]�r�ܥg�_��3%���\Z[�;�^��[�E�V�	@��N�y,/\��.	��f'C!��z<O ���E �(B�F���͵�i1������b�X����v����-x��,��r�gRN�]F��fzZ�^-)ҧ0�(��P��|�<]]��`\��=]�Q�>�)<n2a4L=\k��P��<%+w�eY�ey�,�ֲ,�S��Up�*�l�fq9��:ƀF;�"9�
EjK�tU�����;�=��_�H���>�	嶱Lb�5F���K4%t����)>.�lE�o����3���?0GQ�@c|K�����|B8�kʁUJ�3�����tM^N��6 0)rz���%w���!)Y�G������������KVU��h�в���'����ǲF�>QY�1ރ���lc����3ʝ%�R4�x0Hҫ��V�f�M3Vᷫ|PnN�-{��P-��gq��[�f��OG`�CNNN.��A���]#m�g`-;gu��^��h��I:��W_y����Ho�Y®��2&�!V|��jQ��	����O��3��믿g ������F�Q7C�t���y��)�f�Ç/_�
'�|���ƚ�y��,l���dtz������ݵ`jS�MI/�F�X����1/����'G�9�i�W0���6�5,�`�ꏤ#�(�U����L���H#!�!�@�G/+R@c��L���I��+�t<�X?��>���k=����uE qQ޿8By�\��h4Oh���l�z�����霞��!�^)����|��EA�y4�Q7UZZ����,��熂V�z�����+�[�?��?>:A?+�{�}�Kɬ���&���G�IQd�O����PxFK�	ȵ�̅�'��0�C���1�Es�L����X� ��5���[^�zS�������|6��5HP�IBxC��E��"y�TR\���]ίUN|E<���"�-�+$��:�pњ\[7xɪOC�O\d))dϡ�[�G��GV�T��5o�eY�ey���Z˲,��J�)���&Ǐ����[x@)�0�Oi�#["�S�k���JU[���p�t��y�R�Ԡݠe~pH#I2�p �X<�t��'?�2��?�;��~軎%2ڙ΋�Q�)��Դ�Nl����g¤�$��N쥦8x�#�פ�!����w��.I`��A�G	�����-0E�%Pv��T��	���p���[�)���u��|��ɶC�y�fF_(�xB���2TɎ�ܛ`�bcg�	���U-і��E�ҭ�g}J>4�{�W����W��ƀpv�2�����M��`����cR D2!�S��B��j?�NZ|{w��V�����>d�t~=W���)0fƍ��+��ٟ�j��:�wZ���I1+0"���-h���g�|���766��u��OF����q��6J���qh���~��~���o�{������nZ��l�[�f����E�RTRR$��Ӧ�<�v:��$�5��T�9/^����v�{9XI�ky��E~hZ�|0��n�5ϒ��v������n��_��W�]��3���I�w{��ݻ�i����J�G�8-�!���8�m���<�FqEq��X��6�ON#��j����d��r�0���x��d����x2�q�iw��No2���%�Rc�v\��C.'�5O��R{�k�����p�koM��t2��V���f����dx��Oو���:<<tt��6ﾋ����}��9��
�\�AL ͊"q=t7��h�]�#�u0l2�����d<�	z��`��	:��-�yo��7���h�'/el�"��s�d���9��x>����*[N.��77ߺ~�7�7�����������{�8I?��O=��e��#������߼�d-���4�	�M�4*�eVV ��7�����������~���Gގ(B�/Gp��x���>�Z�;7ޞM���>�����x��ϼ��b�\�餇�|�B�������7�`p�ך���W��j�N҆�HV��S"|8�sŉ:�M�#r���%4��돤�[��5��_�_�e�s�� 2O��"����⫍~� ��$�6C o�PA�rs�@�-�����ik`	��eY��,�ֲ,�S��&f�'�����̥�9V�w��c{��+4�u����.��9ʧ���x���D�#J��j���$Nh��E��yc\��1A��셑g7b�^�H�

bN�& ��|�g�{`k��N��w���yt�\l�t�~�iUC �4*4J"�c-Aa޸��x-[��|�Xd�y�2s���ǆ��w��>��%9'Z-M�Q�JUj�O��Pg�3�p,��x��9��G��"o�kn�.�{��]ܕ�W�9�h8���NqΨ���m�^t����V�Y�n��'�`�W��``-���:|{���V�p��\ܼ��K/e��ۿ�۷�}�����g������O~�_�*��ŋO�y�����D6C��ȣ�����p�$f�!Xp����գ�utt�Vi�x5�m��s-Ԣ�l���rJ����<~��׿~�����[__?|xz���b���� K�u���J��z^���O�� �жqk�p<��;�݅־A�}���r���o��677îO��҄�T��^�U���^�4\��w�}�:y��g����0U��Z�m��GX�i�����4��(�	�_��a�����m��#y��M^�z���8�i.�R(�1�q`<��HŔ���DOX�}XA����B�̊1:C#��1n�L#��ʦc�����'O� #S�~�2
���T�����k�_��_�ԧ^z�a; X�<���;׿�o~�'$]u�Ҍ�ud^�~�޽{0��N����
��7n *���ډ��y}��0|��r5�[�@��z׭j��[-��>��C�f��9����/A"������e�*h������b�D=���F%���x�eib|��2df����y7�q}�]-ϊZby6�`�������&6X�]-�w��,�,�S�%�Z�e��K�or6���J�A�m�^����0핹�HXLVF�6
a�k��>��Ŝ�"_8E��i�Vf��ãǘ.3.>�QA(K`�t�G�vd�?)B�w��?�2*�ȦW�GEQ�S׉�:Q�\�Oz
�BXG~*pq�:/�鹨e��?8C���o�?Fq��c^�����Ғ��̱���[���k�r7�æU�Uy6�]f�E�����.�<���8��A�OܘuV�CT{�F۰�d����y��5C/��}�4�	i�9���w��N�w��(F�`1w��ۊ���X5�qEȷ� {j���zr����TX$ځ[��
D��)4%J,x�H�I�{�w��W�F�w�t>̺�6g��D��A�!ʅ����7�~����7�aR����{�h6�������54yL,Z!����"�V�`����lX�]w&��_�$��F�l$�b{5�O2O����Z��~N]Խt�Pc���\mP����G7H}��Ȟϓ��F3�GV>����4���S���h#PɕT��gc�R����a;�`y�J�`vlȼFؔ:hyV����"�}���P<��۩�Y�lL]fon^�Z�A������>x����`	+�j�	'q4�dͮ����t.\<������z��r�0�6V��oݺ��V���@�}���r���%	�
���s���b�Q��س������4ln[��K���=�-�8˱�$��ƈGK���²��[�uz��۟�z6�]��HW���n��Ȳw1I@��#H��N��r-������}� ����/_��7� ,�߹��o^����e��{�RC�pc�8��uP�o������v\l�V�Q��̆�������:W� ,�>+�`�1��������I2����vZ�B��VF���8;�������ŋn����je�a4����$��A�Gn��6�t΋�vp�"R��vi�N\����&�$�
 W91]�<Cڲ�Qe��A�
�0�a QzFX:lXzq��}�0+����q)l�s��XP�{�pA��%�W놨8���Ʋ,��[�XkY����Ȯ�����~�kpH���q��=o]�J��,�a����;�Z�J�ظA��A�͚f��\��O�'��,7��v��k�}e�kgDա���=t�H���4v&�ۨ���?��jb���K�!	E���$�Ty�9�7qSE����Q��1�]����,�imK,x��=�|f�Y�#�q;�Sa�0U��2CbqγŪ���a|~U�4���7���&ZxÄ��B�b�����i�p���Ԉ��O���[Е�;�򈝒3�t}M�h�z��f�F�~��___���Ç=z�4�$�$��|\9w�����0�(�U��/}���ĽG{`�N(Z)����o�>[��\��+8ϋn��f���(���l��E���;�cY���'�.rPv���X]��I4d�U��kl@��)��|>��f��ī(~�7n޼��u��f>����rT�``"בRV��c]�t�(���n��p���tr���`̷r�|K2�eR �q��Ɗ8���www��;�ϑ��IJa@6[�s�=�36r(�ŕ+W\��x}���/�`89L����w�}>�pᙓ��|�K��KВo�u>���!��mhR���!р^ ,��I��TJ���~otZ�9�^+d2�6�G4���bW�F(��AYE�����S�b��\����w޹5�D�!�V��l���[���x��MAb�8��*G�!2��#�AkL��f���6���� :�� TZ�c~�p�t��:�u$i���]�,gGh��0D�}4�Aú�E�}��+�>��A݄� �P��yg��t�ڭ����\Q�#��H� `�İ�w���^sX���n�I��:��s_*
O��g �̬�f-2ϰ�}�-˲,�S�XkY����BQ��}�6�1��|�T�U����*�����@�[a�Q&��l�pe7���3�p.�M��EI��w}u%�b|�$����
�*=�4"iK˱�D�_���3��7�*(�j^9ݱ5����$�1�a�z�r�?�pa�׈=��af!�c�%*�9�w�Nm�R�}����T��GH�
Ԓ�@�rĂ-)�OM�^ԡ&�|	�?�0a��AA�K<T�j�Ǚ�˾��;�~o��bmj�fPm�⺛_�p���ǕZ�@G: �I�ٱ/&#0j�x��o"�L�(��HK[�Q��Y6)�b�2�};�
=��ȗ�b�jʧ�z@����ŲG����W�^?>Г���+W.>��m�ƶ��n/�v���8�c�}��_k�� 6��:k�������~yk^��$�坷���A�y��Yow:��8�<@����_z`��"�
�Io���'C�5�F�4�,�&m	$��X�"��S��U���I�q���8G�(l�ٟ�q���ι��t4&}?wkk���rC= ��G� ;���ݻ�Y���[����7�l��`�_�|I��c=�=�%�S��|�C���oO��r|���d�`0:eb
�q��V�Ӥ������c[��%�T-������J���m���{�M��L�J��8||*�sn��Jo5��^{^H{D�͠�8K���=\H,�s�������. .�
���C:]�HA���m�L��M%R '~�`6?Y��<�1���F�~?��=�����v��������QL��s���vT�h�^�G�zK���;<��E���F~n7�p[�\��g�\��g��9a�9Ɋ���W�W�^��� .�����n��(^oݹ?L����H8��P��H�eS�&
 - z�g��1r�N{���L��5����4a�4�V�O
���0�-ʢ�I��|��� �!�[��r"R��&��)I%Uʅd�0���Vw�GNk8�hڹ�yaX�_f�.�4�ᚩ-Q=�x���ⵖ0lY���-K��,��tE������"y��KԌ��uTDͻ�OŒ	V�^˴+>L���MJ�)�P%I2�g�[�7�+�A]!,�8�7>�>y�٨�Y�/�ATb-�X"c�Xmt$*��7�7@\&6I�C�Cn�z��2�/�'����W�j-��%�~�T��B��1������� �~!�(ROTD��b�A�5u��t��U�
��Ɔ4��_q<ayWtf ;���>e�R���op�*�ZV��lV���`�bV���R�Y��XS�� �}�����Lmoo�"�������}��_w�^x�(E��?��?��������z�Ɵ������s�=����෍Fi#���s׮���!��m[�����R�,�����i����>���?tm58U���I��*nIL�c�ѹs�P�N�v�t>��^����sxtʵ�[�	|�4�	��r��[]Y[Y[��H��x����k�`��������U�Xs�~�mW�LV�ט��ZT� �z�Ng�=c;ͺ)|�uն\#�$����	&T�I��mJ:��e������W/]�4�����1�M)ά'�P�&�������'''���ݼy�a%p� eqER�y�a$��ni̼i�bte䰛1�5�I�h�������
]w�ҵ��y�Ч��`zZ�iW|xz�����O��Q2��F2�$Њ#9G��xA�zn9\�%��2�2N��Z����_���\]]EA� �0Z�> 4 |A�x]�WL�Q�+`p·���k��9`-��s���]�q�f��f����h5;�m(������j�/|�U���̼�$�)2ZHk�c��M^�]�)�URRH�)D�Q[�j�� hp~i��b~���Y]3�f���%�y-��.Y�q��^��eY�e���k-˲<E���扣05��MԼ����ߵ��%�A�Z"���.����Z5)�P�EZ�,^Xӟ@�#�p��þq/�hD4ZA`4ɓ��s��S��?�'�B����c��+
*`�, 0n���`�:��kN�ƃ��O�٦goAq��N���[��kA�]�����``	�j2�(8i�0CSTkcXgs�yw�ܾ��F��pQ���'�@�YM睺[��9v���U �3	ؾ���Me 3@ZP�'�D)z����͟�z�m��1����R�69�����s��N��D6���ͭ�c�4Qx��)G����Jى,O<��&P�:�pV��+ЉNb5��G����yv�"�n^L��1X�;N�◿���_��mTW���������6�����'>�ٍ��u��`4�D���v+�Ϧ�����&�:�+U�(Qxz�?��佘dy
�Q�������ܦ�����E������������[�N��w~��n��95i���=��1[��'?���F�r�4M �8�0����4��g��n��#a�+�_|�*֠�Ԫ�����;Mǲfv��Zz�������Ȍ�aiE	�B��.�����X�֭{������=@d���o���)���F���0��l�lv�(]_�����Z�^o���݅�?<<@�
?L�8N���&V��̷����� ��OGE�,�J��I�� A��`8��}tD������ß������:����`��VK�	��ԋ�`xrғ:���o\���<'��(����Y��V`�=� X�tS�Q�]�`tBzv!��d,�����;z�P0��l��҃u76Q�Ñ~��4��XX:�b@����t���z^����=N�@�oB�D�XU�dυD(�GQ��Ӆ�>������p0�g/�� lЭ,˷�=�v��*~���GB)n�L��U҄b�4.�.oZe��Eޒ�k6��6`�v�ei=ć�=�3���et�,��e�����8RAQa��;��^�.˲<EYb�eY���*��Qsl�g%��"�`�c�0a��ꇺ���Q��Mv�B.�n����qZ�.ƄH��T�%���}��~�8�>�H���n��b�@6�9l@T�sZ(��a��(K�\x�|<�QqN�����Z�E�d� A>�GX�rP��6$t���3�!ܛ[5���<�*/�9��]�,����̷�|N#�X$lñ}�)b�ᐿ5#�X�^���4�V%I�+u���2��P�f�-ZX/4Q��.��)�D��� f0��b���Lf������愘��j��{���6؈��1F��������>�1����} y���r���A?=/����wэ��d�M����@��Z o0�Vʢ� ����vK���+++Lk���d� �T���yh�1HP4��pxE��3>[��rH�Fz�9==��p��5��@�c_58>���>��4'�B"��� p�4�����o�+�j`PS�Y���H�pL�<�\
����Z��C���Q����`�W3}1u�f����Č�R�P#��r��,f4�->!�d6���f3��o5��d6�!?�������u���6��E�!Y�v`�.��%0ڊ�2��� [�ȱ�����t�5�ؕ-�D�4;�ව:p�#D^+����6UYM�8ԚWr�`��6�ee�"�DMRD��'���l�0?�R�����$Џ�G:�c pZN�U��%�N�[���A��[�����B�le����]f>4k8�Ft�ry�Z߾}��� %p�����ɚޘ�&�*��#]>��x��eY�ey���Z˲,OQ*���`�UzF�!�2��.�?��W�+��-���-�=M@��?��<��I�NlF ��RV�M�t�x2�3�w���}���^�)8<����#~�qe�b�z��sT��L4�sTg&�ľ����6w1@�����;LP�;7Ã"%	�|�)�e|�lp|_��٪�ba5��eP�K-�l	���MY��"���;�
���%�Ѫ�m.^+0��]A)Q��XB%h��)R��:rF]��!x${y�����" ��mX�n6�t�Ӌ��)����oKWj�!���Y�%�Ղv�5�3�*��p x��Z(>&�:��3+%Un�����p:>>��Xs�Vt�P�^��F҄a:Nt��W/l��7��;d��_�������/}�;�������+W:�&`����>w��kWr��+z�*-�¯~��~���КaTO�B���үz-�F���s`ϳ��Fc��(�0� ��C9���_BGdB#�����:A��-3O�2���
H��X�6���E�ٽVG;��}�����(���y����'C�����K/�4==����Y%�8�Bۅ�ŅLrKI}���4�
&(�;�>f�P��d�@�����ѣG0�׊�D�9%�B �(CCi�\:[_�G ����a4��R���'��&9Q&=Ǒ�ހ�@Q�d2�����qm�nܹ�}�0�tr���H��0�p*N���A���v�ٻ��;/�xmme=����k�̡
��3 k�8D_��g����Vwu��L�s�Gǣ~�ouڰ����z4?x�@��`0�����
����H#���P���o�T�"�=�v�I<�BF�T��Ñ�G�gA��3	��ݷ�_O��dxr�hkm�o���^_�_��G�3V���hx:Nie @�s��(�$#߳W:+�tR�'�����(����k}B�8�P�ª�����?)M��)��@� �7wo}㭳���Ƴy<�I��m7Ӽ�Ex&?��$����d8�L�!LqfVٷ��=��.IY��D,��qE{��
yEE�\/�eY�e���k-˲<E��0!zqV��b1�K���� ����r�S��+�V�+M:��{0�F��9��Jʊ����$K.�Z�H��mn#����%k���C6��a�

��ǜ��7��!�9�9�!R(�O��|�F�W��ȕ�XI��� �'�6G�ёi�jgW1�Uk�rcVV"���x�خ"��U�˕)�j��#d:nqDd�J�QTޏ�&�%8A�'7)�W|����Z.�_m�Y���xb\�е��x�vC���5D���o���jf�4k����V�z<�H�HJH��X���uJ��st��稵���d�ç,���S����`���7�	r ��� k=|�gu:�P" ���&��������������#MAj��d�K��{%J>PTJ0�������b�1c�Ow��ͥ7�� ���C�_y�e�p3�e�ȵ㝈$�����>G��ZE��"�U� C8K�A7JP�d��g�.�� �0���`��aV
f;q#�Ԇ�!���ݚ!��
`|3�ҕw+s/�B��� ���IlI���j�!X�#E;&�N|��}�J�p��<��^��q)XN����Ɓk=x�`k{Z�t<�~���Bp�Uo�χ����T8ӂY;ܡ��}�-� y���.�bҜ�B����,�TU�	 ���t�V��+��(�yGI�SA���$X�L7�5-q�IS���m��lkk��0`���Eڌ>�F�]9�Vz�3;Mb�����DO=�}4���摇����»آ�B껝���P�#�P�Ф�+�2q�Z�"�er@���搰jÀ}�Ų,˲<MYb�eY��(�z��SU�{��*��)�[��=��,�P�$��\m;��k>����BO����}q֘.E����|�E8�El���r���c��δG>3!;��sv�)*�ps-��1��44He��6���I*����6Ǭ��RX�����	24n��-8*˝y�D����rn�EL��]�i7���9��pEP�)At���;(��Q�(=���s��t8� �LLɪ�ذ[��}���jbp6ӭ�pO�-�f"�����+�cSwYK�]����>Q�b�9�&AZzDc@�u���'nJ�94ˣs�3�$�Im�<Xl�^x �g��ӯ��Z�u�s���o��Զ���,dV�#�X����W7�)X��}��l6k�|��u�����������>������L��6}�{��XV/^B�Y�� �C�%y����O�GF�8�f0Ơ�)�2]X6�`��F<�";aٔ���(ql�I*���{Y�EQ�*Gg�<�R��N�o5�x�;w��������677��)����'���o~��Bo}���$�[�.|����k��r ����B?�_��@��dm���O��?��� U��]"�Y�P��ddS�S�ʎ���ڂy�Sİdܽ�8�0��F�<����y��ּ$�H�DGEFK���,�3�;!���be��|����,~�x�w~�_v�-?
��3��t����f�����8���he=>��oݹ�!�#
=�߂���-����x�5�+�)R+�����}�k?����x��� ��;=q-�:M� �\�'m@Z������>���@�w�o)�(�P���zMbt����(�h��4��v #W_�ځf��!��$K�>�a� v�A:	��L��w _�O���W�Wu�ކ?x��|+3�q�N� ���1}��H�KIΜ6�V`T���8˧�4�|2��'*��U@�̅�\Z�Ԉ_�IAc��.]�z�*���y3�R١Q�nׂ��ǡG��Q|��X������-�ֲ,�S�%�Z�e�QK�N1Ĉy-�G
գ��:���&;�N$�Tyγچ������η��]�8������8"�-a��bA	�7`"0e���d��#�Ћ+!6�tc6ޘ�� <3��_��5@��\k
Ue��Y�ju�B���2"��9�u&(����-�3w����$?�n��*���W�����9:�e0ȳމ��u��<6�7��d�̸2�MRVs!��Vb9k�f�2F��.�?D�d�k�8��J�D!�3m�P��H��L^�'h�᳷����n�*L� ;w�\�������5�V��C��mTz(�X6l�a ��gi����GK�i�������� U�m� �x�[עJ�8��X����1{�$�LtN�.��E(��Y�&؂�?à�)�Kn����vww51Q<ˠ�����#�T0���a���ٍ���t�)ST�\�m�����<	��hp�*T����m�#�{��O��aP5rȆ����7����݅�����	y����wv8'�Ç�޽;�c| ���6I��I�s3=yi���K�y��`�V�
��D�� 鵼�*�h��|�.�q�/.V���$S������կ�.���7A(Ns�"��y2V�3�	�"�u�P��	�F��oHjC���N�Jf�O��l�>�"m���2�e�n��j�ub%�pVI������h4��fIѥ��$��*+giQ����6��3�,˲,?tYb�eY��(����j`d��T��� /S4$P��)���l-;`��������QM��.c��Q3�\=�2[|�j���s=��
�*��@�d}���  ߏ�jQe�e���2U	���ښ��ٿ��MX��	%B`���2	`pP8�����'C�00ukkːZ|x��)�\��I0&�(���%jb���
-���-���<Z}�B
�*g#ZIV��	���@��y��Y�=Yӟ��gE�)��,cT�G�J8QT,�]�M�ƇP��G1CN�D#M�DͳQ�fqheo�8+��V`��_��D{���,JF��9Unͩ5��:��Q�HD�&n��������G�����i�a��	ڹ�C�o����r{k`�������y�߹��o���_=�9N��Ť��|����\�t4U�\���v\e͓8��xų���
��^���j{%Q�ۍIT{��0Ő���$�t�L�<�Kz�]�kT%UfM��r�ȑ�.l��**��;��r�f�*RG�������y��w�۳`�)y�ʕ��o���v1�O���^K�:���|8|����og�"�J�9A�@�3��q����ʐ:.��x0�{�s���k�޾��{���p:���q2����G��l`���(r=��0�0)��k�|��0�Q�a����� Pj6��E���$��k�bf}P��s�_8|7x��y����~�߁�Dm�S���xñ`:��z�L6K
O���^���{�{W&'��S@��#����[w��q@G����?666~�S���L%>�L'N6�� d=���p4��Z���Vpr2SYz�,�����!O���W7V����!���u8��h�$s�n[bBG��c�
�䖏F��]g������i�j��>����(Y�#ژ3�;I������kvz����YRd�|1��JF�͛ :��ND�a�码���:�1b�<-W ���٭:+`M�P��y�y�C�`�q춼���y��J�}��l�<�X$�(��Ԑ�$��ɂO��(��.�I얮4	�eY��i�k-˲<u)a ��-�',rQKt[��u�CI�,�6��MZ�Z<iF�7��3|*I��d��j�Zo>ru�BpJ\�1�`���%��»��xS�P�l渘�F��(���
y�@۷Z,�EYA,�q�`ڍ���(u��p���xB��ur���j���]�l��5M�����kWi���7`�Q��S\GQAt�o&협�7TU}㙛�܏��\>ۭ��I����de��1�m�b�)���UծE*�87�S�����C)��g����N(l��{q�D�  (E6���:�%�pd��xN`�pB�����ܫW�Ҿ~�:�\��t��|����:Y�|�ӕ��Pe�7F��4�Q��E�KI� e�A
0������hyȕ�	��4��.ir���.�q�^3YEw�D��t��J��PwQQU�5��X(�g�ق*Gs�%k�aSJ �3�Zˇ�N��~���H�$��	���ײ�U���zB�Ef&�K3BU�i��5qyE���1�<)�s���Z�a�J�g,�,�$)Y,��"_D���Y���Hn�q���G��y���˯^���<������M�Ll�l��P�A^x%��A�X��)���F�� ��T���}����N&���E � �S�d�`�%:�ւ3����)A�[?�*]�h���˜8Τ�a`�r�|/�`�r�M#��dωM+��H^���ݢ,7LZQsKP�k$�aU�<���[������QT�Y�O��S�)r\�D�O��%]��V�n��G/!ֲ,ˏZ�XkY��)�T�F�	�Y0P�X��t�$"h[��������
���ߡ;�ĸ-!X�ג:�b����@���&�#(�p��C�E/�^Q"��fEf�]��(�V��1�����/�in纠dY���y�T=e,�*��'Ί�S��N�� *T��ܦva��?��Ŀ=88`3J�
�����Wef䌽t\Kfp��b�,��	��.O֌E�������
�(�#��,�¯�HŞ���:�:���E����`�7�v&�!YR~�#������jT�o!�׎�����)Ԑ��h:6�+T��|Y��	�իi��mD�n<�wUI��4�@2��Q"e3�܆�r�HG+#�s?�[��`������A��Ҹ��<�h�-�5Y�7�]���,5���B�4[���Dz�W���`Pz��Re��> �yny�+�<�;�8}|�%�N��P�{���j���(�ٸ�_~��$��"�
'�ݦ��6"����tq�r����E�ᅁFYK��K�e6V�BW7Y)H�����z��S�,/O� �R�K�/��sW!��Y����E��n�ݿ�����qrt�<����Ϟ��w��]+�Q�w4ܑ���*نq��r*�"��x���30��sP*�VE�I�s)c�aK���D��U������Z5Ҥʹ3ŵA�ؘgit���DJPtR��߮r�a;xA�Өm�\������r���]=��=7 ��*1�ǁo7Jte��#<�5&�g��u���N����Nއ���-�Ͷ���1zv<��uE�D4͋4I�1^1�N��T('����y"�ž�.�0�Z&�.t�d�F�,BrW�o����Ǉ���<]�wJ�(J	-�5)��x��y�,����)���v�Ftm;�L�Fm��|T���8aӰ�Ա1��`Sf�F���}�G���Cg��-v\���H[ǵ����]g}��k�ЛFS̬��EWN@��-�~�YV6\)+@��V�%teL��ᚐ��� r�&�4�%n���P���0^}�/��~��ȤH4?�����O�?�X�eY���,�ֲ,�SYEi��	5i�'�r��l�$I��_b<S��C ��j9y?ZLR`A~��'��>#���B&�,���,���m&Ȋ7ke�6�߲S���z�I�����U0�p7C;���N9��.5{�'�+�BÑ�8���hǸVi5rZ!(��g$��.KJ�3t1%��0�y*]2��8�0	���ʮD1�"!_)���,hWس��)�F(�~d�E��*J���0��1(�Ҕy	3B8
�{�a�Sy/��
b�d����O�5e�AT	 l!𵩯u�}�Pc�rr-J�lA��HP)��D�j����4�� �U���3Y�+
�EsI.���	��K�tVg&����ٹz��w���x8��}�x=߹����f^��l��� �U�c��a��Ͳ4�����#w?��`㫅7&GH�U/P�pÖ��-��\���N�ɱXx?Y���}�ܥ{���%~�7~�0t����5K�Q|Wø�#k49=����6%a�t��!�0���n	�k�/G�ڒ�:{�N�8?W�iJQ�V�Z�7Jx,�*�����r1h�yx0p~-f<d����)��x��PM���N's�3p$yGH�7%1Oz.�U������h�S~γ��矇#���s�����kI�>|x��1�!��"���GGG�����M���Ҝ�c!�.z�><9�Z����p<�Z��m�Oᓋ/2�����9��]�{x�8�)Y���}zʙ�����]���(q��4��$��>E@�~@����� �lТ��^���A0}�ǧ|8�����cX��=�V��0�Zа��)���=�ia�-�8�8��ô�\kaWa�9�7ǧh[�����ii���Ur�חM���>�Ύ�r��=�T \�e�Q�k-˲<E)��A����
������Ѕ��n�� �J�%�I�ǽ̈3�~���p0f7qH��Ο��~_�S���jq���{���t\�]��`�"SIa�K��#~$s�V�0Tf�\�b͊��gs;I1�?I�|<>)Fcd�F�<�9�~.�4# �s�.��g�C���`W���mw��B�ʥ���G
\�,K$�NlO#nq\0��2fBj�&�f�(��
c.�0y6ܨx	JTÚ�|x`kc��j�%��ЩB/@�U��l����~�|<��bّO��Q=�1PV���щ�9CS�"��S�)��)��` �>�Z)Dl�uE(+ d��'��D��R�Y�%8��a�>�,�f��- ��(�Z.^$'�|D5�l8$�p
�G��st< ��7۫~x��}���4�P�������y�<z�w�T�˅���6 ��� #h�h6C�7@sb� Ӝ �LJ�J��v�,FJp
 �SR_�+4���f�
d-��d@1lv���Q��\�r�t�̯���<�}p��o�y��9��H�f��fs�z���<֢ɋ�q0 2��;Ċt���ϥؤ��G�&�(�%d�		',D�.ɝ��syh���?�y�@e�:�����̆�S�<8z`�R:?\b�$�R�^XAp��*�x>����PA��<F�>�6;!T'˳f+D;>@d�ڸAs<��Nz͕^��zacg}�~���7o�N�pC=����	�b�
+(t��2w�~��*T_l��3�{E�HiXR��i�L�b{}�mvB���t�e��d�;��H�w$,'�'��:[y��nV�GÉ�{V����&�����,�"wa��L�n�kX�NR�p��͡�	�P���������{����D�J�Fz!�_P�g�4ST�@�2�.��vp)� s���@��Լ0�[��F)N^��C~ϐ�c�!�K�%�,���?Ή�i��k#�2$�"&�Ų,˲��e���eY��0���e�-CO�+bL���O����L��KI.($��B;l�1���%e������|9�( �4�L��E�����N�Ccf�~mmM�º�.&�j�9�*+R�����e00���ՈB)� k�6�2��1�$*�4�!.5���Chga��E
c/^�v�|���1T��8�p�"�)�A�(�0��=!m�w� �RuC�'y�̙����#_H���H'@Զl���9�k��0	E%��q2�X����T�P#4�̗��N	�1h�V���k4#�IW���-�Z�oF��mt���7x�YAi�jz�2�u��ԯ��L'4H{����0H��σQ��,؋�lJ�)%�Yh�6I�?���{�B3)y�պ�WF#Qf_��mc΀�U���WVVn\�paELi����<O�E�Qd�>6p�^$z�={K���ƿ�+�Z.F���� �F�s2�G�j����������o><y���}��i�W۫�w��������ɟ4���Ō<T5e�)��deu�}J#��_��9wWH��������o�J0PVj��;�2Md(t����<��_0IJ����n;�!�Y���v��|E���p<�1��
�8���=���Љ������~���o���?���7��00~�>�@>�A��I!��N4��<R������P*c	M��0��9r�Tw%��|���5�Bj�Y��NG޾}��e(�ynk���e���f��D�qaĎ�#l.�1��z��6�`�Cy���B��W��-�B�+0\L�Z����@����ZgIf�hςtu���N��#c3T�Ac�q��,R�2+N���}�(*J�iiF���:�_-�XkY��)�k-˲<E�S����fl�X���*vj�3|K�-�U���	'�w���!hR�M4�D��5�]L�$�;�R�f�=���}̸����6;8::988�ON�S��:�P�{����` ��@��֒�W*
��xm�Y	�TA�Iq ���o�Y���2�&*M��0��"
��x@�D �TϕTn�͠+�+�*
�'�p���)&`�� $���j��Y�(��� Z�e$+��rػ�����*0ᒬ��q�G���25)Y��4\��>4xLԓ���T%NhpN�͜����$�6-E�-��2�w�]�Nմ�-��X�R������9�K��wmC�|�ˊ�����vx$ӥB��e�4O�F���xER�m�X��h��rIH��8�!������%IV3GWQ3:�s eQFxC�Y�������Z�d6v}wckMN�F{���i�%z:ڃ�_i�ʒ��؉�eN�zd"�%-"+P^N`d� HOޒ�Of`%b�.c����nqZ;�/���k�@�E@,�N��NS����h��S�h�� �d2��o-��ƹ#��E�y��`-g)J�d
)n�Z��F6b;R#9�C�-�0�$��:�g��AN��cllrgaU�p�c���y�����%�u&voč��Vf�U]�ͥ�-R�J�4Z 2`�5?�۰a�����0x���hLk(�F�lQ��koյgf�����^�x���FE��.��̗�b�[��|�|#*����m=(+G�i2%2��eEp�@�$f3�����O��"YP�tS*yi�B�Oo+�.�(��v&7��m�gK�*���<�����lq��gI��ʿu�&nw~J���8�H��[M���3^�60m�ahR�.T9��*M�ً�E��0:(i�U�be��:-�s����J��p(�^���"/��:�ʕ+�ՠ !-���Х���^`hC+=P��=��e�`�f"ރ�&ה��ޞN�Ϗ��O�}��]�$��s����Ш�f����C����Ãɖ�=	2DFWf# ��ۀp�_aP��%�
OnyC�% �ۄ����=���@�:0�
������r�6�d�u�M$�m�˵�ڴM�i�k���Z�^iB�x\�͛ZQF�I�I�>G�����|||�ގûw��6酟p���	�IX�T�_�b���#�r��^�]-�!�:)ňU�W��"v�!�O-��㬚$o�qb���K!���L%�Y��t�hҥ'C�����������N�����������=88�/�fC@�p��|W� ���r�Lv��AQ�c�ye�P�Jhe�����aZO��k1�]���k�/���ߺ��6�M~^3I�$��ef��O����O<�k7�������
q4щ��u���L�*���a/�����ΟMH�:r��_�%�L� ��8.�lam%����:�nC#y#j��E����NOqXo ���������h@����G?�����w����?��?~�/����c�Ba���X�uΪe���L�m:�� �!������Y΋{��\���(�O���i��GGC�,��}��Ǆ��x�/��\�גE�&6���v�^C��`4���|�'̳j}�k�ܐ\)��[KK�5(H^&�pD���B�zt�T\����#s���]�:-�V���`�A�;���.//����cP�"�iJ3����ClA;�x<_+�uĽB#���*��0Os�RZXJ����U �v�qe�"k6:[ʐ��=�񋄗�f�o�KӚ�m�W^y���;������E��F�j�\�̹�K_Afj�����[��s��b,�+;�t?��S�-o�y��u�{ߡG��@�ci~������.t�����ΙѢᒱ�kV�m�5�Ea�v�c	KDtSz�1�Lc��U	��q�ݚ�����(d>����[�ʩ�7¦mڦ�C�kmڦ�t㜉6i���S�X�fߡ�=.���u�aǧ�� ���R�X�Y��Xԩ���^�R�F*�ʅ�?Q��!���6I�d3�'�\��c���3�P��V����.���ä^��ھםj݊0 �buW �;ac����`�b�6����6��i4�{�E�!I��h0��oAp�.��}L�X�E���ot�Z�
v!�.�ҥ���V�yhJ��uu�މ�_3��P'��:�?�'�!$um4����*6����BIX����YA�T���v"���`�~w}��6��] 6X����Aȑ�*���u��gU��5)Mgj��t
ų>���F�V�;��L.Ӆ��^�s�ȫ��<0��ų�$�t��d!z&�΄�-�4쇕��:����� g����o�,���/~�������^��^���Mbt^ۑ��W��i��B�%������$k�)��kμC�T�{��C3"���_)�!�Q�*�:\(C�qR@���jQ�Лl���gO�IJgX5t�%B��h5�*�.�I��2�D��U�u��m:f-�]h�8�62�g�5�
YN���x%�ړѪK�Z4�t�dӇ��L�*��I�BoU�F����	=m�
�zMF�k��d$PE>8�j����Y�4�{ҹ�y�����F�N�E���h0���>���O�>;�M//��T"|��MX��	r��y��;w��d�$M	��U����ң>�%+��zQg��s�2Dv���A�3n�7�"m��ˀ�P�"2-S� �X8��3퇣 ʀ�{[;�p�hg<�J����4M��xH'�&��ѬL�0
	F/�3C+�F�3�����Y��ᘞhw����0&�=�Q�> Ne�H'Sp/�a7��I�Ya ���x��e˚�3ᎷdyuY�M�h�ו�s<�����c"����4|\������V>893N ������zaU��i����kmڦ�DC��j��Oh4���z�Ww܂�,��㽽�yqB��&��3^~t)H�c�,�rN�ľ����%Ẏ��Io�Y�DI�Jƍ^�C�y�;�8�T��S�BVt�T7����!� �_Y��@�K��Eè�
����N�G����$�����N;�LD�9=�4Y6�^pImM�&��S�'�y<��d������u�Ȯ���u�t񇮭�>����Ҏ"�*�YN˓^��a�']G����nvu���Ҥ�\+R����VH���:Zέ���Z����e(}.�tz����cI��lkkKn P� K2I���U�Z���)���*ZV��TL��>��h>G��*I��������g����k�х<x�$	!��O�"�lo�(?��VB|���	�d�}�jp���i���5�iZV�b�y�%\��?ܚ<z�0M�ڳ���g�9R��c�Rx��D��FC�!���*YU�������A��y�L��)��ܭ�vb4ju,1���kV��ri����d�8�nzw>�v�S]�|�fU��u'E`�'O��$�V�^���chL�rVg��c5έv���}��f��u4,���J�q`��<j���f�j<R�Bq�����ȥ�� ��D2�=#��4�<._F#���C�F#���"���NNN�m�6=����7n�N����2�Oh{��7�ٵk��=�J=z�~�������������|ao\.��;j����t&>&/��j�il&��r�VY��U3�U%lv7�?��,�R6"�b�˺��S��u����֬��ڴM{���Z��i���6tM�ɜ��p��!K��,m��nQ���1�8��t�|�VQ�ţ$
Q������-I��\�zU�𽦖���u��mq����ͪmVV)����f����N�w���6���)[��3RŌ��&՚�����\�m0X�B�e!0��-��0"������ G��c�X��.3�,�\F32���v�#�D�1��Ȉ���E)A"��d���qA��C�P�[��DX��%�>�@�õ�{dle�:�P���B�IfP��[�R���.�R,	c3������tK֡���+�s�gUV�E�����H.{g������u�<b��ގ��a���/:�xl�֨Ed����Nb(��q6�$6� ���-[�������+�'��0��UU��a� ���5����
y/!Mќ���
��"�	�� u��jh"�旊 �6+����v^�եr�D�'_�����z�?�/�K�Z�2O�$�AE� HQW~l	�@��9Xmȫj�Z]m;�H�Y�U�\2)��馢�x����4�S�i~�yVW��ԅ��xp��u׋/{�E:������a/KP�v>K�ܹC]Iֹ)0�����w��)�:2�AX��@b�" /b��T�d>���x0�xNH�#�lE��-����YB
�T`aw��6(D�-(�Ͱ�MӄJl�ѭ
,�y+���31�<ZY�ƕ5�O?����I%vP�EAHK�>Cw� ;�, ^�uao\�U)b�Q���ȸk��q \��˒pԲ���Y0�����V^V���x�zUp9/�l	�,��xЧ)B�<vaLK^c�9���)LO��9T��|7����6�Z��4����ʢ�-y�3�S��
�QU\��a�=�<;}~���}�����{�x{L;[���0��d]u����}T�;=zv~�|z�|4�cYG�/��5BkAm鶓){C�Vֆ=x֊��J���<4���~��-����s��OYq�Y@A�9pZqE���6b� �}�."�(�`�aZ̄3��4:t�X��t�"�E[����}x�S��i�����ڴM�i�Z
���᷼׽�:���$��Τ؎�X_\�-��-1��L����k[�?q}��^N�{����{ۻ�C
֖��� �*�:�D����&��� ����|�B�	�PJt`eB׃����Q#��X��d�,�$\�d�-X�Bq�0y(�(����)��Y�K�Ja�J�^���m�ٶ���.�3���6�C�|�<�$�wy����S ��#����A�f��O"'�,d���E�,w�8�]�f#��命�`�����?� ����Q���@+R�ͺ�ؑ�%�M�Z�j�%��s��ѐ���q��;���W�a���n� f�e�:+:�����aϴCh>TR�zG���gg�?��|�k_���G�������ӝ����.����.����-n��1�U���y�%�ZQG�%���̙tI�݀�G�����pk�ꫯ>��߼y��#�oQ��-r�������Er� �?e��,�{�=�c��q@[˧�\剈��ٿ E��AP�)Me-�6��=@"��|K����|��ǲ�q�A���lF�E�Ң����O,c �H��ɔ%�e��bY�8Ď��b�Ch�m?ܥ̑q�9v���~Y����� :��P�[*�� ~�ģk׮ݹ{�����V�>���z��{�gXf٣G��u��̖��dR1K&�$�g��&qyD1�������G�	�e�iK9�m5�S����3'g(�Nڐ�7���W����QC�m ��{o�%����·X<y�K�bMN^��kW-�)W�����A�����?/s��'�J��6�]u�U7ɻ�y}�kywu�J�S�/	�[��]�cEoF�F��SV��i��2m��6m�^���%D+�/<ɴi"�ܺ�����e��3Zsp��aZ%��T�d��1�#�=��12,l��3�eӨr�`���s���N��J�`��&��dG��J��W@�bƑ9�ɖz����L3L�-��|e� �.���f�ne������D������}� Y�������oV,$�����ٙ �������}>���z�!�ޖ��J��҅�|톻d�\̦���h ��?�k`tr��+3���2�`Εgp��8O�Q	�C4��`�N�@�g��Ik���xΔ ��izȼB�9l��CׄKMj�*�n������T�m�.~�)����)�)@ҮnҬ�b)1j�����ϳ�Tn4�xFCaO!W��,�f�&˽o}�QřN`aK:��Bf	M�Xy1����)V����|��[�Q��ݣ�r�����7���'��ֽO}�����_�m�w�֭�`��f�%:ᛞ��P�F�P�t����j]:�\��,R�h(�\�4�%�փ�'C��WkHB=R����Sz���_DȤ�5����]��
"����p�
4@&IQ���arY��n̋�=HQ`�A��[g�V�I��G���06n�0�g�T~Fl��;�P��+Eّ�lͣ.�Tk��sSl���4ID�:�GC���Ѐ࢕�ߢ֜�'Vb�}�l<>�}�ْ&��ˌh�H��q�?�n\�������svF�L>���wv�{=�����*����	}�;�^���S���%�z~t��3�s�#� uV��07L`=��cIG ��-�%v���4f�%*����Y���E���+�3�9>��>�8�C8��ܿ�|����'��_�������ϙw�}�.}wv��D����*�n��^�4yХ�c�����B.�Q�	mȴq�c#�ʁ�y�u�#F�J�,��@�Gӆ�B:+׻�M������%q�M�p� B����@�0��X��e�~U�{�ae���L�E���Xk�qݻo�6m���m��6m�~ڶ�$J�֜�϶�U+���wB&����%{s ��,�i�c�իL,'�^?�� d�6�D��NE����Y�>� f�5`1	�_p%�J0F�Wm�O�GYN��z��z�ag�w8M@�8�$��ESQ��UԴ�2�lߣN��O�̾�O��/�E�	[�3sE2��jɕv$V��gT��#B_].
��%���N��#���fUkU��3���륉�*֏@ �B���C�7H5�q�)�9NJ�������Ѓ��dV`%��B� fZĨ$	�!%���O�<��fWL�gzdE\��8��áU��ٙr�W��4moO:�	Y09[�N��-�����Q���E���$���ׯ߼y�������Jto��s��W�f��/�����_��� p�c�$t��^�ѠGvjo8���AJ^;�8-ZV,y�e)�j��E��a]к(;��m�DY�ͼ`��PU�g��ǔ�Zv��Ag �=��ø[���<+��9��\��$�8G���%��$fBP(|:����3,|(��)�c�	��7�ܚ<@Y�^��ⵚ���I��FY����r��u[_q�&�:ֽ\�^ġC�B�4z��qg�>X�h������9�*���tN}�D6˖%J����iC[\�&]3�E���Z�k��h��X�{�myw�=>)v������Қ\��|oo���o��oi'1����s����� ��X��p0�m��ɻ��U��]��՟���۷�ق��Ͼ��[�����������2�g�(6�8�j�K�,7V��UW�4`-̹��v,S�����k�M�N�\
H�m�$�V��9��\���O\Bmڦm�˴�ڴM������
� ��,�tV�Y�>��Ժ�MF�CݼS�@{1�ylK���:\C:Xa9��h��G>~f+�*�O�o~��qϏb�e	2Q�B� �V\L�.ŵ%_U˷��UpU�k�!K�9�H��Slه���jDB��/��9�P�b{����s���w������ynB5%I��i*!i�ncۑI�V����e\�0kL%���S�9 �<R��t�$b6�����;ؑ�S��7&��� �X��W�of�kޚ��X�(a�"�U��6��la�R%�4�zkdx�:���iҐ�z��Zt�\=�|����X]�j�䠖@�U����A;��n��l�BN��Ϯ
���G��v��d�k�7��@8�ZEVO�[&���?>W�
�	b/�i���)��F߄��a��g�D�X/�2���n����{����?�����6u������.|��Q�CC�v1��N:����X��,ɫ�Wk�	Q V'귮�Q�p�{,˨M^�yq�=[o�<{��=|rE�7 ���訪�pg��ޞ�4�	��*,��W�mh5�_�a�,�ǔ���gx^����mUR�GɌ"����5K���2���!T�������l6G
�"�"�V�(��)$j�J�A�:�n�}ʗ:$ᯫ���C�'(�N���O���҄�8���h�dq��4�����ۅ_�&-b�3����1Ç�P��y�A�BǄO��O���������EY�N~]�)b��h+$�,��it�����xq̓hP�І"�����(;�<�� K�d���%�����v�
��}�"a�%	}��0�eB;To4�rڀ�_׋Y�F�eYĵ�⾚g�޻���G�ߘ-i�z�����L�,vWV\銣�銊�`��ԿU���+��JU�u�'Jζ��g�(+{u��_�ѺU{w�������Iʯ2=��8�	g��ҭԏ��d!}��M۴M�d�`�M۴�����N��[�$MH
H���T�&߼(��g�8 ���Dۗy7ϖ`��\�������������%P&{*�T�s�w�@~S�5B�UtP-��,xU_�!�`� ��wG���Ւ3R�k_�C��
��
r(��k���$�&�7��i�K���}�xuc�&���"c���y2���WX�p[��g�L���8v���u��*)���,'x�n��v�&|TWK�oU�k�L�䬯E-������C���7��][૛nj��R/�8~��D�ߖʐ1��	�5Նj�N���e$*�a��lpyyYyx�Y
d��Dg��A�d�8F���s�5.�J�豂���O?#�]W�L���t����+����o�����Gϟ?�O�����o��'�`�?�`##��B?�`&���P��-'U�S��Z�s��T?���y��䂶�����:��N:foooƸ1���Tb��A>����,�YR�
6�W!	*i'�m���i�I#����Ɩ)-�#+Ky�����A��]+�'����DЯo��ϲ�H��oRd�f�f;�Ӻ]֙1͹��mE�9hډ�.����x�!5&F<ˑ&Zr�Z�}��07S�=~s\�M�����ߏ��~/MfO�<Y.�sGTdl ����IșN���hL�y&a�O]!�x	E���zd�<4�i��磋3I('��
�ps��&��U�V��h����Nބ�y��)����E�b�h2��ʘ��y���r�-P��2X���l�%ړ��V��~+��ڈA�2�a-l�<:�H�;�0��Jn�
�GÈ3iyV�L'tr�smN�<�'^d��i��i��i��ӷ�"�.�1$'�j�Xkr$�
+�I��_Sa�U��a��`TQEIԚ�-UTl#l�I�v{G"�@��CzRoh��;ׇ=!�'}�F-C���Zd�

B�Z�0�3��\&��A�I&�1N��ى�*�����U �E�XNK,`D��?��K��d*%�[��
��X]<c6^ք2*Q/D_q&�����!"����e�(K����+u
��֬nWٶhX�Y:�v�
�P3�Z��խz��Fj+���^VT��Cx�#t%1=�m#�}�*��-��b'�P�3�<�O��[)�\�D�"��%44�<��LWk���Z4����u�Pzb{���iB ���u�<.d�U�r�7)j�����\.O�0��
�A��q^@OJ�h�u��1kֶ(T<��z5!l��qN���ef�~]�����Qo2���#�z��5 �R�˙26!X2�8ۯ�A�U=�F������V��_Z�����x�0�9ta��`�x
�_��O����*��k�*�����L�2�&~�]��IFƕ�8|��r��9��v �UUˢ�2Ry���w��iUly�-,�W1t����5�L�-6 vg�GQ��
o��^���ak�������*魊���dhFG��ߠ>�y=���vlx��yg�l m�2���Lx�I��f�iY�<�9�'��.�w��G/k�w���i�
�Ҵ����������p�]W�&��t�3�ZM��Y
5YUU���\:�<�O/.[.�E|"�rMP��aM���d1�ȧ)�\!=����wyZg�J���)���r�ƽ�(��Ў�[!d;<�:� ��,P�d��J4HU��/uTݰ��պ�"֟�����-=X�UlO��yi�F �D7�9�i߅�Os(IhR�:|��d#�ۢ;+ɳi��i���Z��i?m[��V?���"��5�Y?M��n���G�Qj˶�k�h��W+�wպ3EP���z������_~����1��,���KE��"��*��:�ɺV����B
U/��]s�v�y N��@W988@��hgg�.$����DB.��///��)�t��+��j�D�[l��֖0i�ኃ�Z 	���z�(ic���V�S�#�|�	�/�r<�[W�1�Z�-�Q���~ք�4�$��kF�k?�:�0�bF�y��D-��Bew{�J�{mU%����m��%��r���	��Z��lȲ4�ڤ�'ԗ�gD*��7�h�[ӳ��gGs���PP��ilB�\r�qHcT��pgkwww�������������?��?��Ͼ�����/�ֵk�^}�M�����/�_����"�rƂr�6in�h�e	T�>�ࣻw�Z�%3P��[�Z +&���Y�ĵ*��I��a\�H�󃘶0&�Q�������>��σ�;H����O7p�A!s�4uϠ&���6�0]%bk^��dhR$�f�i��u�1��VK[5�K�����"?H�wDY�� xǥl�m�ě���q5����2d��&��|��|~<�����$|��c�l)�=��a��)��6G���]z���	��1�l���.˂��rNSfF`��8F"����݉W7�a˥{��a;w�І�m���I���˺��4K�'P��DO&�z��9��8�P}�8�[R�u �"�����ÿ���'OQq+�#���N+�2� k�+�����u��V~���ПM.F�k%|�Q˵%�˲���Ɍvࠇ�L)hv�̐��q�;t^�Ⱥ}����\˽����k�6��m��i���e+��j�0�M���+�M69�ʇ��C�X� pR�3��k�r�W�h/�?�iu���Z��g��9����W�2=d�Ԗ�+l�}5�>?=����(,]M���<�B2�pb:ȋvhY�b�l(�?c[YB���b�1B��@���>u���>X������ʢ��S����dq��?����[٦� K�$ �^��6�=t)�w))W懑&�U�(*�J���8�XY�!��d;WuJp��JW���&l�U��ܞ��Ki�+j��@�G,��t���oi^�?�;� k����VL�Py�mc�T���-S���Ke�IlI6\2��,���j@a�;��E�R���Y�8[)�J(? T�� ��$���B����ȬX�^�H[�s W�� )��>����LT{��k4�*LJ�7�sJ5	gZ����}���K�Y%�dgUhB��W��\�����A��$�d@�Z�^�7BWmG�7�R�"?-�z��n��ظ}̠�^�Yz�(&{�blz�����${��d��q��7n���^�����ݍ�h�����F!+L�d����k�鍭�K��6up]5�����w\Ϻ2��������
s�9X�Pq�� ��4WY�q�*�s��I�8�m�g/��4��I��^LC�d�"����&͍�c�U�֫^`�6OL1d�Ym!:j��O��r�q����-�](=��㦬��:@U>lC�����TJLUeB�v(K�~���b>���(�0�kI�[�A�ݠ2`��*#�0�̠�˼7�M"�u�����0W ���pa,�Zɖ\����!J1,p�z;C�d���T͕�8ρ�)bT CN� ����p�0��_��C_!��+�w�Ta|M��6�pG!�	��Co��������`/�ԏ�Ϟ�{}H_L��ߘAړ!�ii.��T���%8ikỴ�D���2�����W��T���\"��k=˵ٟ���p����@�D��U��Z7 ��4Kk��xp���=C�j|��Q�`��믏hI��u�� ow
_����Fm@�gi�4"2i݄�AT�r����8�^�ٵi���kmڦ��j�u�ղr6�
]ę����+�t6�$N��Z$�8�K�Mb�P=d�̘������|v1�+W����P����FOK%+�N:Oܥ�H!J'�B�D_찖�(;�>l���Z��V��쵕G+�r��YS7���E{�u<Y'�Ӑ�������S(�I�g���F��3�\01+�I���%C�ߒ�J�Y�)�vw���ް/�c� c.�E�T"2e��r*E[�������_�����-f�B+)�쁆޺�故l	�3��9�F��&<c`1��:�5Ys���E�3rkˠu��BF���5y}^�B��/�D�6ZU���1-3y-=��ũ=zTYh��^���������߼6��W�"7C�E=L�#�[��������>���w���%�*�yr��͟��_{��������w�߿�W�M�#?υ\��wyyY��[o����%����w�L�������V�x4���l~F�B6r��
�%�0���U�I�I����L��\2��w�e�5e�XD����)���Poiު��?�%'�\�*���9��_�\�ʧe�Ӕ��I0M�I��8+�s�Q��X���lwZ]�*겕���^�ި	g�.V Z.���)�fُ[�q׌g��(+�X;16���/����\ö��޾��W��t��ׄ7�ϓ�@�ii5�C��!�4du��o2�Ǚ�A��E6t4�ߓ�P���j�Ϲ���g�m��#\Ԝ{��w5|9�!�,˓sP������<��NI�9j@e+ލE4��!='B8t,T��4H�C�T�wk���dcK�9at4!#��0�5K��5��M%�6`�*cu)_&�fW�M1�O���G��...��H����B-���|ߴM{���Z��i?Ec�:�+�o�f��;���U��zZ���;�#����h%&J7��CO�.���U媥�G����4�����;C�_�֫+�=K����A^Q�l��)VM��-T�˜���L,u��Ǳ2Dr�����8U9�O4^���>G���<\�N0���)�<�ML�6�\=�W{}�6���9��S�GMsF~Y��GVu�Ći!	lH��qaOC�a�ǽQ�/Uy}���~��1WߪY�����'/D�#��A2��]�7������|�cߨ%�Γ�*۠��u��x&Zd
?LB?����bM��}�O����\D]�TM=d��a�Ʊ����K�&�zA�RUƧ�)?�}�
٪8��z��Rh��^��;]�y*��5c*v*��6��(
����=}�������iT��Pm�l9]��nfa�F�q������./N���i�̾GqxV�C����|Z��zZS�.Xe;�Q~`���52#��ܥ�����lyqq�����I��=��Y�f�9�ؔc�P�8��'�NC����j~�][������v<|�W�u�r9.M�\��՞oz!�T��:�=/�R��SE���U�����*+�fT���=i�К+� +����,�
w�+1�FA���N�G|�ct}���ɩ+�c��q�YXne�g�
�eKރʓ:lp��Qj�2��<�R�*`0V.2j��X����3�X��9�M.9���R�YQ��S���/��N���^�7I�J�*Wn��pM	q峸�0��Wt���S5�:$��).f��o�(�9V�6�i)�>U�_��h��r�0�vh��r����ӄ@d ٠^��|>�����v\kB\��E�a�%���7�(C�C.<E�;OsvA�r�L��
YA�!�В�9��r�>��8�Dd3�M���9���Ȋ�q,Dx��(�R�J� �9���T��Gr�8~��xvD~x�`���ݿ����|��D�0e�i��^p�)o���<-7���i/�6Xk�6�%����w��wM�|�R���Bn�-��?�r��[Ch��p�QAVT^C��a���n���{GGGd�\�r�5�$���ַ�E�F���s�DA�^�t*�2�hooo8�ٲ����\������IRR���kJ��f�ʋu�3��L�x�w��ZѼj�1Bs�d*��X���/�r'�~�DX�= �[,f�n�/�C����E���>U#H0�͢"a�zTFZ�8Ҭ�B}�h��魭-�VT����k��`�,�|3�r��)r�cD�aFj��WK��`����%�������k�o�&����]�������>�������e��4�\dQ2k�u>o�o��Sd��b������ �X���3�$~USK�Q�	��-ҽXL	�\������ ����YdE�#u��RY��E��,�c|N#r����?�~�98���p�`�/��/>|H����| �M3��CT���dr�ߜ���ٙ�>x𠧽W^ye[�,O�d7GN}���4;�甧���Ʉ:��LI����J�9��&�-��Vq�
�thб�^ĥ���yPv��^�����r�A%e.��}�B�B�-$�ƿJ%��D�s�8vy��8Y�ԁ�	SMJ!;�:9�X:��Ύ��sk;�I��AaV�Xr������h2�XX�� ׋c�v˫���2Aݲ�y5���/�LX}D����~��1곇{�]^ r� �:�t]z:��6B� O�V�d�[=Q��
 ��Rw�#{��-�\ZںUﱾH�5���Ӡ���ͷ�|�;ԟ���A3�����s��E�֣�?��?��7���_�՟��/|�_^��d�~Iq�������c������RްP(���崽��V�V��ْ�F���V�����left���.�&E�"]�$@�2�t���Js�t�v�Y�ӝ�]٥��կ~���?�o������W���~�e$8v�6m�^�m�֦m�K4Ǌw&�׸R]���i�k�Oubǎ�O�6���OU�~`�8��5u��X�
N˘����ꩪ���l�u���y��bH�բTEj�.\Y�w�n���6qm"���G��&[Ǆ0Z�l�T��?�r�.�����x��m^vL]٦�3ҰO�%���ȷ!IMx���H a�
IQ5�$:�F0� �g!w����^W3T�*I%{fM^YM֭*81���
��B�r�ڠrW��y��=<�������,M�	�,ȶ��B����:ʫ^��A�(q�9V�����YC���\�Tk��iнh�UZԮGX����Z�?w���m��}Da�`�B��.�J�j��E��KgQ��]0X�7��<g�����P�
Y+Է��������:�aB���Ĭ����RP�0[X�x۷�y:�`�^�����r�`���g�������v���ӣl�a F��w6ݛ�>�{�(v��޺���hpp�v>��7�mTY��z^o��Y@��`�2�[�UҨ�L��YS__�w�n8&P1��g�A���^]�'cw�%�=�*��ɧ?�x��]N�]6;�{��":q/�z�������e,�@��PW��j�4��j�'Z,��3ئ&wQ]�b�jPYH(��EEڣ��尬�_D�'(�n��zs�[iϠ�ZN�g}�c-�2��$���u|H�.�
�3@l*�8F4k�J�4ƃظ�K���d��h-�pc7cr;��g%n�v-_�,�B�]`l=IKZM;��v���^��+��ӼO�h�]]��z���^��#_�t�I1Wvb�y�#��3!�0������#�?����*�H�\�B^��s�b5y�H�Il3�|jA�q��I~<�߿�>Z��eJ���v ��>r�蹱*�#l����"Ϗ��YU������*�nh�W��Fj#? ��(�$�lŹgʫXRx
�*�Җ6i7�L3%E�R^�?�^i�� �2��4W�V�F=�D�K��7��8��kЗ�]���Q9��gb=�ڬt����+���-\R>�����Y��~=yj��E�A����8����'�7m�6��i��i��r�5�����
`�vՉ;+��r��l�����R~�\�ﻁ��R�DL@��!Դ�g2���
��+�<}�\
�k���V�J`�p���������#4"��1��}�U�d��guk%tV�����R,W��X�Rb·i]�Vr���ca�<�59Q�����+�҈� ����3�"��+�(��t���1����F;64����a�fxj?F$�	�>_K�:���M:���ςv�$�Ḩ�z�|�@SR�f��a��tz4?%��Ƨ_�7��Q?��!�;���,�i������Q��Dq�z��;J�#�R/�����^ѥ񈿜�]��q�M$
,��<ۤ!�)w�3=���v��|6��١!�ϋyC�'O��{��S:�ա+n����;<<��N���)�[�b�9�ћ�M@��8���W�J������Ç���Cĝ�[�n�����AJ��|����o��M�lϳ#h�y5�ە[��r�:��7��*��?|*��KV�}Rw�yj��s��!��vr1_�C�؃����~�}�k�՟�)��:�+�	K��w�VDQ�y^8g	}.���=�jxLkFCY�r<]��zFf�fm=�|{ͣ�b�\�N�"�<�f��,]��R��]&��TV\\�:�s�W�o�w���O�I�,\�d�mM�.��cߚ�X�*��ٮg�~(ʕ��$��8�n��=��CqBhXf��������3�DV��<OH9���(M �U���R�U��f�c�����J�|�᳎��2�A�:����d��X�\�cy���#���� �5{X���e#Z��ι�/���bza������<�q���l��)�	�e�7����i/�6Xk�6�%Z!�m��m?g��F-�M, qz��xOy\,v@��޽����$c�_QuJ�k�p����hʫ�?Ư���/���t��o;���'A=�	�'�B�3���f�s2��2v6�(��F?��������L�7�i�;=_��C�%�P���@��m�TJ��a4$���1.�JV5lt>$�Ȥ��at�z��$d����%Y%�X����0�R,����F-6��^�?#�p�,�"M��U���Si]��Tiz@R3�btH��}eyE�$˺B]2���MF����}������}��UY�L���ᄟ��,f� ���[s�!B�<��+�Zz</�B��z�����ߧ�/�A���Nq~~����|�1�F�+�<���@��!��0
U>W8��t'�(�N�Z��y�ա��s:PtY��ʚ���j^{~�}��pg�{=ֱ<M�-��C�ϭ�ぷ۟f�RC�c >����A|��%٬#hQD�>N.z����_x���{t��������^�,.'�I�6�ܿ��G��������VG���'���1�*���F����Y�V��Ǻީܓ��~�׿������׌�Խ�������]�TI��O��c��w�_�������m4���~:��i�|��{k{�^#s��Pz.
��e��Z�3	�-\HS��ivqv^��]�%��-Q�A�Y�CP�t�5��;U��kZ����*4A�L=�bt��F�!� z7����i]Q���32�kx�ހLgȯOFQ/��Ik<+2�sF�����"�6�t��,zQ8���2��;�vG�7f\g8R/D�1 Hq�b�sh[T!j�84�b��4��^q�g}�+7�>]������e��K��:��"���*�j�I� �
kM7R��*�B�w1�&\&.SZ.�fP�@#7iN,��(EY�y��h�,e��3F��_�G�AȊV�<IkgΦsB�a+����.�$�g���-�۷o߸vh�|�&\O;p�%!?��"��uA����+?���zK .Qv��gi�1>� ��ڤ!hk��I�C�:N��U�Z�c���s�������Ti!��+
�U�����߸v��y��� �)�;ޢs�����M8��%5[�դϩ�k�	����ڴM{���Z��i?M[HnMcJx�ծ[Q,��q�I��#ݿ�bIǧu����R�#+�
���5��rL�*ɲ�1��VY���i��[ُC�3�b�yP���
��Ո*䟅n��8�&�B|����j�@Z8\EgB�ɢ�?��ZN�gr���x
��T�E��*�>  ���;���4�V���.�����d�u�{��,ɯ�ؾR�+�|�|T]|��|& �p�U#Fϕ�>1��1�����j�p��v�$d��'�g��*)����M�O�T�3c�wv�7�,gT��6��j��s�'t7�t�l�I<�%fU+��Z�I03�م�u�`=S�������/..@��hG#H����(
"��n#3���H5J$2s���I�A2�ri::�^R]��[S� 3ZҝNdeN}rr�/�/4
�+����ґo~��L��硯9��ɻ�;�<|=�Q��ϖ��� �!@�*I�bK�/�J����L�\K�h����t+S�H���\�i7:�Gr5�y��F�����X�EA ���$2sD�]V
?B)�@1q��(%�(�9	P�ٵT���nE��6��"��!,���s�Z��ġ=~�x<��k�����&��Γ��$,�S(�bhe{�v��>��9��t�5	���j�w��/v+�I�l����9�J5Xwr���ɛo�9��n޼iX�!�tggw�7
�MItN���g�_�M��e`��^$�&���j��|�Ӭ/	Z�#w{���y���O�����LRo����9��<�!�'B�� �8���a<�r��F�x����ˎȒ[�k��6m�^�m�֦m�˵�uㄐawde��ڦ�"V�j���5{��p�):���im(�7+}���,���2�E���*�����>����G���=2&���#��4�}L��b2*��k�7�cȁ�Lp�C�:����7��YH��I�"�����V� 5�#�ܜ�{e5���;�'�ݍm��J�
�8@��K��;�vE���MV���V�����bG?�ֺp�C��<�|�����aQ���ȞfׯS&��^�(��Dy�����"y*@%��Xp�ߕdk���s��[������z��>b�zV��Y�uf]�5��&U0A���΁�*U0��z�_h���A7�z������ы��+{;���?"���كc:l>_���yz���& ��n��҂	=έ�\#�UT&�{q	%7���*~��aa�F3�a����B���r}[����R�r�ʋ����ɝ+�a�b�W����?����O�X>B\�Yf��x>;;��g�7�����%�?�_�����w��+������gOQ��~��)g��_G��}�6u1�Ͳ� ���V�_.��7_��(�y�D$�9�2�8>z�[_ێz[[[~r~L���o}���~�������v4������������ݻ��_����������7����5�G��'L�d9�GaHx>r���	�fy���,�^|�$�g*(F�}J��� �p�*�\d)b�r[�ܦ������u�Y��B9�v���,G�6ɒ�Ӥ��M�in�<�����޶!~�����7�,�ʧE@k��LOb!�1����t6{׮��&Y�5��c��eHf*�ط%-����t?��Z���	�L&���k�ӳ�'4N1�\'���CV��M`<H*�z��0{
�ڳ^�B�\G�C���k���*(�s�9.;F�@�����K�3�#���g�0�Շ�����Z�gt���ޝ���SrP�j��N��W�⬀�I-�M�.���f���1�Һ9j�,�Qq��?�[Z)YV���a�@D[�XW{��'fU\Ϛ���T�by��Jkx����S�G4K�F�5��+A]D�|t�����[_�җΓ���i�f�~?}����^<|����g�wI�MW*h^~�w��ul*kmڦ�{�kmڦ�t�k�aw�F/|��פ%�_�֬9,[Ρ����.m�&�]��R��
բX��7�#�)�(�BhP�a?-iIR��_E%��ƍWɪ��g�/��("����?&[���'MJ��f|��nᵚx�DM0�\�^���(���s���X��A���ƦZ�i��ҭ��_� =�%���\Ē9�m�BVb��JrN�t��h$A��UEa�zW����IR��go�V�x�u7v���r@]4�kV�W�����Q�����g2v�}�!p���������t�G}Lw;C�-�P��x:-��
7�UtRQ�Oh������[�V#a6��P��1�%��E��Ν;�݃��>�����߇|"S(4CT���ur<����7�|���] ϼ {"o�����Q��IT��FWM�'C���������Hޠ$Au�jt��9 �G���H�8.���+}�p��E�O����''�W^qW� �pf�����ޘ�OPwuT�t��P���(�b)�E�����F`3*�7:�<��=��m.?A��2��U��8�w��n���@6fҚ�\�	�1�<���ZV��i,��$e����^C��*�봧�m����+�״�?�r���WU[[��U�ףn���'cZ�㩵�X<#<�*���ϭ^k�ͮ���6h[���݇roJX �R ,G�&O��� J4!i�#�ҏc�NWG�3�뺚`�F�[/�N�iw`��ҽh��B�N�Y�LY�^�P�*�5+Rf�L�[�K�<�)�=���7�$���{|i��h8����U�%R@v�&������+���w&���e�C��.-��
�gO�EH���.l~mK��Z��i/�6Xk�6��[ 0�9Ӣ�~X�L�E"��u��((��'���4���e:ÚR#Ej�t�U/�a�[���4W�b�b�b3:��?2^�=у^=O�%��?/���JUV��J<�'z�.�EhB��d<�ԽW?����b��w�S�)B��SX�5W��>�T�~��c���Bn ��+���v�D�QߥZ�`�5
:���Z��(f����{e1�������QQ��ㄤ�`�p�{�!��֌� Ub�~�t��a���2���A��*�U�x�<O��[����x�̰�ԽW�hR��0v��8';;��o�:y���# Ý�VS�������.�y�1�A)m0[T��K��o9����"�t���6�:w�^��럟���^V��쎞L��l�Lv�u ���,�x���J�"&��+�>��K��կ�(��k�vbbB�:�mI��,�Z<`Q;���i�r=�:	������u��k���q��X�'��%�e��w��կz��>;_<}x��wޥ������N���=9�<|�Vt��Ӌ��?�.Jhև������gg�`|���s:�~xpp��\�	���0���ӂ 	]��2Wy���3�$���� �@���Y��/��߸v�}�ߨO�ONN��'K���6_�^�ٟ�tP���ۗ''�G�{'�OG)j�����[����ݷ	/�O�P^?��4.��'�YV�Ӥ���&�pooO��9�>)�xԏ��tWY��L���	"g��Dږ��F>gZZ�n� ��W�r+N�k}.�cE���dL;���6路_�U1��ֶ�_���|eg{G^`���Um�n\��>��]&��]=�r��)�i]O}:�H�+���o����C�@���h?��s[�4�~ J5�l�������d^�L�ݻ��l��aw�{��35ڪ��&/��}o<��ԝ�����k���u�A�?�N��;0=�s�J���k],k��֚�V��~�������L#�hbB����R$"��wCD^�E�.%б7���j�uB��*�O݋�,C;��}p��~�-�����m8�P6#�-���Lm���+�P�E��r!-:'u)*�.����v\>+g�G�ShJT���Gn�������h'!hG�����>�d��CW����������0��O��s��<y����[[[Q��3qQ�5�w�t���M۴M���kmڦ��m��z!�G��[%������'+���܋���j-�C��\���'�9�YqEK*5zY"�:���+����;�}�]4m��м��;��	�����p�� ��F�͂�8i!��e_����3��vro^�$"�!�\B�v�t���s�j�s�����{���k��l4�W�p����?)�� SRQ
,P�a?��0�lj��ڪ�mP�Ià�
.t�P�˄��W1u%�+�r��'l B杻�I�`����.�C����V�#l@_�z�jrzA�P3:�ͤ��T�B�M#'����yk�횀48�=d��J~.�ʣ��'B�:���a�`� �"�.AE2�}�睝��?~�qk,����݋$��D	i�=�>��ޡ'�&�ַ�E��r��p8,�Y3o�PjXQ�]���ݾ��DQ_FPs��u]�P
�r�:�tZ�Z�r:��bJ�[JI:�!b�ӯto�_������p/=�,���9=ce
����6G�*� $�=�m�f�>�&��жQ�%�u/� ݊nɵ���(iI)erL#�������ԟa/~��A?B��A��=f2���ѕ����a�'9��%Y�߇�/I9s��V�G�)�4� ��/�:\.1�-e\����b�eg�+/y�I��A|���:BO�mz� �+����������\�T���u.*Y�hw�&��W����~#p�aGu\���[ iT�M�t��H��V�`kL�a��y�,�}�~κ����)xr~I[%�\s�wɊ�2Hm˄c��O�,K���:E����!��O��]=?9a�U�� H.%=�����w�}7�o����6�9�ц�iv��������ڴM{���Z��i/�֑�+�oq�
�`��ؤ�Fv��!��}?0�U�-qũ[�����-��N�0��<�_L;{4�;Uj��E��_���==CW�T!�̐o͞Q�3+���]�-C��Q|����������ؔO��R���U6����[��?9:~|q��H������U)�����Ò%g<9_��	B� J�NI��X�,���`n�dI��7�L�"��Α���53~U[a��e��#6VMV�%h�e����8�B� fʑ΀n�h2>>>���(�߾�����e�XvgsJ+�7:G��+pB�"%C�����扯� $�"���r�T��	_5lnBG!�L��x��8��b��C�܋�W��-�=��y��?+�(z���x��Ȑ���A����9Y�.�J5t�6~9�����Ė&
�ʾ�^����"U�w"@SE#��"E��(�{�0���a?��w2=ug|p��;�y���a7;�$+m8�࢘^�߿s�<|����fM�$י�Ǿ�=����ګ��zA��ƾHp��i��鑦0ҋl�|лdF%��f�(#A�HB"	@�ht7��*��*׻��=\�;�f6��zՅ��q#<<�=�w��#+~q�4��H�g�G���������������>��_8{������g^���p��}��͏���l�M��j^hr=�˔$V	���);�V݃Uj+c��?|��'ߦG��[����0��~�ӟ~���~�ܕ�W��ܸw�Ν�Jsssc��������_��O�7��믽�:=�S�`��w�$[����P������3�я~d
�wܽ�`���5��1�{V�(�6<�@�F���vi!	�T,t�ul��o������df$
0�9w�����յ��~�U��a�\�x�����𐦁H�z�}ju�~{ߴ�8��lci��y����R�jwM3�|%����ݻ���g���_�Ǔ�w���>�R#}�ӣw���WZ4�g�2�����8��,#�Wo��nߨ{Ͻt�iQ7¡cg�I*�p}�{�$e!�a��aX����@N���XPLP�f��Q��Dx[�<�RU���y��\�
��a �u�+�g
�u�(P�)�F�HHr�_� F�D��hQW%:��TŬ�����'I�!}W9�D�v���G^�r���+gh��+©NFK��������/�`������]��v����Oרx�rUd���Hq�k\�mJ�������������g�����У#������?�����|�Lʰ]�������?Am�(h�Ķ��YV��S+�E�A�!���8���P#�r�h�ۼ=u�c�y������Q�?���ʘ�q5��;+���%X�S��yf�C3��L�kL�K� p/��TL��.\���[o?�v��c�޲�d�]�ڏ��ed�H+e37���#�x�O�,Oqu�~!k@9��]�
}�^O&���C�RM}Ʉ�`��f|f�+��u�H�n1X�(}(�������QG�˪/l$�'x����11-wѬwZ����2r�lds�sfY�آ��\Hwt����Y�d9�bRΜf��N��@x�~�Y�d�����)�z%�[�B�O?e��Y3�q`���l�r�V�	=OZ�SS�n��u�����>���U�����#^�>$�h6�����v��%G�0>ny��zL�T�t�8}�4!�I2��7-ևE`D^mllxށ�:Z�~ћ�E\TJ:<<���@���X�E؉>'@p�~��H��o��<�y�ԩS���zk�����ߦ;��C���tw�#�wm������$jH�se3��4_˃�tf3��~rp�ҥ�9	��1t�F�������(�x_W�-��w:�T�)7��<���:<<w�4�v{O�<A����V�W���?�����'`K�y]�ؔ��\F���XL��DB�(�Ш�ׯ���4�t!lz9�vΒE�aĺ�"���{=����FC���J��K��/K���z@���NH#�OB=l�}:���ۄ޳8t_x&��s9�� �3���"�W�@�j���'�g81�D�dee%��:/0����c�4fq�Y
�v���3٪nY��9�c��]��_�.�3sV��3u�I�*�ZoM$,u�\y�ј�h���3vA�W�6�p��$3a�"����|�_8u�-�0hli`A����5;��|�#��ks<Y]]�g���|��t�V�9���{2�T��Tӽ�ȹ�q�ףp�c���@piC'�ꦭ9�-])����.�Ҋ�JKr�v6�4-X��ح�51�<�5o���m���mޞ���J*9�*>�J�߈J�V�K��w��ũ���-����I��9�R�Y�zC�+O�&�B��*�Y�pl2)2eD���6^��x�����)d:.��qZ^�B���q#���Nb E��3Yol�w�*��a�1߱r��wp ѭ�ao8��B�^�&�:јBQ*��*8i���(�Oj�&]Nk$�!�(S�c0�r% �<.��	��d�AW�E*�2N�Ty����Ɋ�)>�Ś6��VaZ*/-)��,����+O������Y�nm4 ���t�t�ŵu��T���.���m)i�YYy�sG�d��q�vB����~��	�s�6JA�f*z��"J��f�����yM�AC@��� /�+!�Ӡ$���N^�\<v{0��ĴDX����:G+���P���՚�t?�,���<����\8g���-A3's�<G�w.͓"�<�h�7��W�r6,hJ�����m�h���dP���W.?z���#��*G#:����5���<N�K^����0P�?讔�卥#9�K�rx@�e}m3�d7JG������}o����<�:M}�uW��h��642�p�������)�j��]�T��f3��̴�7��͵����T����'��Ѱثooow����n� �xx�G��i䗡�6�q��k���i�Ŷ�^9�-�ÒyrsiY�YϹo��V!���t�R����{C���c��CK�!�=�64G	=UY�T�Zs*j,�q�L^�p-km*�$:��$���=٥��^�x�(��y��J�ô;�U�r�L���=d:�T�^��|��6�.J(e�V�@����f͵}�Y�[4���B�Ȇ�IX1�hL+t�2���hU�E���]Z_���J�3�.t�n�,/
���o�%��P��yk}*��I
q,�(�Oi���/a�� ���l�ڦ�o���P���K3�ꌀ
<T���� )x�yEm/�X,i���t$}�Ц�\����-8.��m�P?W���J,s�n�]����J���������n��o�j/~�#/�c��έ[��F7�_X�|�Q;ۏ�wP�L0�:$$ ��A�z�S�e#���h����Ԃ���w�o=�����[?�1x��N�B)mSxʴ�ı�̢�=f�8+[�Hw�'�
��V��J�ҩP�Y�]̹1�mޞ�ͱּ����f)BW��~%~&�O���.�cw�W���u�_�ZU�`�n��iĔ�V������c]d����B��'?���v��n��>5��q4�މ0]6��M�*i�6F-�t��mBe�8fTϨ�^�Bə@M彶-s�]cZlWM�f�-&dPhJ. <D�t䊰4j�c��ʏ���q6D��O�`�)C�����L�f�C����%����zGv�����:g�y�@wTh�.m��	��Y�����#H��z�#M�ѱ��U�S�4k��I2;�C]��eՌ2���V&���i��1虶?���Ϲl�d}3]��(3�\�<��-i2��lgXShuqquu����k��TurB(z��o|c��n2��W�[��w���W��կ������stt�Ǽ�l�2�/��N����Ͽ���ϫ7�ɾ��Ph��I����3�� �`wa-̙�qΑ�GI�mqCe�K8��h�f�,�y�[o#�e4n���~���[o9z>����ғ���7��2x��҆�~�t	���x�9���;w��<����<DuD�|=E1c-���8OQ�����n˘��M}'��bF��z�⹈�hO�g,���\�s�4ͫ5��lH�Y�{h�'=��a�V�`3B����A�s\T8��L��tv�yP��T!Xrxx�,.cǰM�Q�~��и�;�Z��z��w]�E����
@���B��Ĕ/T�4�O џ���p1A�LG�p�'���;6ct�l��'�vF�o�8>6--�as}�J3�G�1��� @պD�������ݻ���,7Z[7v��+����@	��G���1aѓ�=WOD���*x��0Ĩ���L��ܒ����e#�@O!������Y0�"H�݆%�W9�
�t�)
����l���T@y��m�~�6�Z�6oO�J!��f�$�� qP�.l3��L��o�S�]����P$�k���]�(*�eE�Td :��Ә&���a�
bi�XŶ��;	��/�\�;{y���&���aB������s���x����V Q0Ȅ���%���T���d��M�M<�@LG�a�`��D�Lf:�$uLR唜ed�l��P�$HQ�B��;/�ƕ�� �!��k�-�_:W  ���5@	�Ř5��� �`���a+E��2���K�|е������)Y��U����Bg!w��;��R��d����OYcYpԎ�>���Nv�a�[��COs����z^.;��D�Ʌ�	W6ݖ�����t���4N�����u#�-��GV�S�s`��'1YoKN(�P5�+�����u[�F����D.�"2�����!Yg�ї���,/�>Yґ388�~����:r�|�kxd���S�5	����E� u#a{X0e�X�;����]^�r���E�^���� W�е�`w���}c8�'�R�j������0^\��kѭ��o���Y���頗�7r��~����{��Ý'O�z��|�q��B���䍥p!���SҔ���y�V���[Z���V�WZ���}��I 7�������]_�8v�$�n�pj�вh%���fp;gvrS!�
QG��`JX��b\��h�f���n��L+��d����mZ���U��Px���w�T���].�*��[�G��.1�?`���,!�Mk��K3��DY��XV�!������l�R�xDZ^=.c)�oz�|<�%jd�脏H��ɬ& P�MǍ�Ĥ�G�+/:O\ ��$��µJ[����Ħ�v�5���H��(��Ȅ�\��52�-;�a��j{	ͫҤ�Z���.Ği�$�G&��y�qi�Qd[	���2wlf*9�~U;�ӧ�ȢUC�ؚrP�e8K�wN���s�hk5hO����${�������N{�M��Wɗ3�,Mf� �+��rC�5��������N$s���;�<�^r[�㝺x���6��������?��w���S���'�yaqq���K�$~�}_�=ȡ�9�뙅S:�SШ�my>���ܶ�F-w�(�4�t��fM4[^͛�e/�cKe��3�B|9��_�e�F�=��ƀ����-�Aґi��f	�vj�Ue3�:?�3��b��m���6�Z�6o?g;���Nű���٨�JM��?IP�`�u%l~ss%�V2�Y���0��?�F&9�.ɠ��p�����@�z���һ������e��%'<V��ĤSL������yB��#ra@UN�Դ�D�S���K��5��$�E_��2�hb�57�n��e�fJ�1 W�li̊�\W`�V����w��������Vr�6������rh`�h��Q���f���A�-���Y�.�}��|�����www&B�T��@~N�*q�����4-���Mb�7�%��9F��������y���u�H�ǌ�􃅅ǲ��׃� ��.G��"*H+xO�΁�I/��p�.�󄣗�=CI胎/��s=�gΜ��_N:����\r������n�sK�D����-:�5=rc��)���Qn��_�U�����4�����<�&5{mm�����=׼{�.w�d�w�݈�MG&�ݜ�\�*g���v��U�Xn��p�F�tuz��=ͺ�@���٤?A߲�U�@�V���`�C�v17u�H��Ŭ���#��r�:O���uZu�J�ױ�@�z�t8�cZǉ��"�F0�\\�g�g����8��4���T�d����*@UU&�v��/��*upF/��v����Iku�*�5]�6�ͽ9�5�\�e��:��X["���Nk�M����ף�WS����u��3ʰ��.�'�L�F�R�/g*���<����*���YU�+�������O`?�m��Wj�?�\���O�f+a��[VΣ��9,-�u��'�1���t�g�h�TGF_�FxD�(�&��L�&xz������̇&��&���9' `l����iu� =n��qѯ@JI���#z�x"��B����iw�B�_R�SMs��0j���_��Xk���)�!�b�Bg!?���, �	0��o���4��y��
3Q���L��4��l�j%A�� �ٸ���Y�Y]�@Փ��^з1P�o�q9i�Aa��$�Vi�^�n��!IG�L����Oe��u����0�1��L�f�n[j�qz{O���
k�,mj���'̦Z@ptj�A:K�*��%)��CL�y���U8ͅ�lOX:�R����w������AV�B�J!  >H)�d�#���+�Ih[�ZN's-��K K�!�g����%�Oہ�r�V<�@��+��q�l=ƥU*�z�@��l�U�7��t�<�hE�� �5%7��47��wݮ�vd<B���[E-�֬̓"E��5�O&�J��Uk���,3������vE�n榻���|�^_���X8u
��E2k�:��#0S�ٟ�ɟ�n?����4WVVjM�����G�Q�{6=��(T���@��ƪ�v�a���/�Q��e�a�\'A���<~��~��tŗ��������Ǔ�]��$�R�M&����x�|=��/��}��Q��ܻ��.Ϯ©-���wv���d>�M72I	QHyj�n8t�ah�A.�{��o���|Pk���?��Ps�"���܌hLb#��d�?xb����0vO9x:N�]�D�[X��$J��� /7=�iZ���IB��&T�9+�p�Q���}�Y���2�~�)C��[��@�Y��CK��9�V���2a�u�<j#��t6`F�ӵL�PH���Sw���P1_Y�.+\#�N�������Ї�`���aC�Y�i�Ĩ�L׶\â�2��,0l�謨脏@&�@Ǵ�茥�R� �Gێky�� �=��@X-�(b���W%h�ȃo�6}ۢ���F��Qn�ÿS�DJ�Mo��Ii�ʬ�b *�t�aP0��O����v�0��?�5Q��^Uv4���m�<ւ�tf��t���������:f'2x̕ �Ep��0��K�'�>M����?�ܳ�v��M�n�9Cʗy6�y�]C�]x�����%�����pУ;��︞C��!��R�%��ֲX����Ȩ7��~?Ndr�?P��3�<3�E��а��2�lv��� �y�4���6�Uȃa@�|�%|D��Cz�yr��^�s�5o���m���mޞ���B��ٍ-N�����~K1�	��dW��)�Ob3�uy,Yh�dU����Е1�훑�]�����\Դd��]��M9��6AM�X��o�E5(��{cL9���c�r5c�݅u�BZ���I<;���t:�OKw�4Hpk<Ax�P�n�c�5�rYUY0��`�pm9�H����Y��T���V���9�	T���j�.u��`Ϻ=�o�<�E���`��R @��5u�CÁ
l8�a}ss3XA�V8`��I4���M��D�پ�����$���s�9fZ&J��.�&	"-u�����J8��i�F���J�o�dV� T��#��1U|�l�{7nܰFE���G�y�2�EŎ4R΀�x��"���YY�)��PW8`�`��Ԃ�a�p]���A�T!S:f!�s=�J�y�9�����hR+�F�훈?rәZ��F]�����$2倛�1�$� ���*0]��z@e��]=C�L�u<n��</x�G��r&�A�U�3�IZr�q*��.`Es�l6�B��A����J]MK�zב���?����8����)g����SQ�u�U�'?�R�Fx��B����**Z�YlP�U,H�'���.GԹ�Q*���D���J�N)(��.8x�B����\�b��b��ը���ji�̖ǥ�z`tܚ�.���q <�h?������4�g;�������d1���)���g��f}3�˶�RD�6=nj��3�(�q�~��ƍy����P=���X�d��w�}���haa����ZY�Ɩ�N|{��,�T���X+��9�C���Ѻ��NXY&�▗��x��I��B�e�j�.��xs����I=O�]� u���9��;�A1�Z�6oO��Xk���)�4�UӨ|�P�"�%�D6�SehAM��%�#��܄���ͼ�L�t 6�Ԍ��Vp��+}1ˍaHgl��7��]S�z�<Hz!�V{���7��S��$CL�4���� �6���K�dQ�!8�uF�ㆰ;=�(ٵk8x���f��\<��LƼT"�lM��(;�]F#U,	��㌯4h!����K��>�ΐ%��?:9Y�ڶ�)K7�@���<ښђC&S��R��
��(ص<K�a�3~䱑l9�~圮���U��y k��}�m�2k�V= ;�h7�Z.=׳���0t�'29�F	��ܳL�~|M���T�Y�ce#�O��hlmi7@��F�J��\"�R�!���E"������B����7o&y�[���P'(��,$��eJ;Y��M�J�����d��\~�x������2���o��{�'��]��s��!��7�>��φkW�~�Sm�Ig(#O��X=��?���j��RGe�?�d�{y���f���� 3]#�����=s���:�;�fѸO�Z�[�������l�nmm�=0ηj�u{��A����2����cg����Q+t��Q�ݜL�$K�zF�c؞O�5�"C��C*@%��*�g���<Swdq���m����^�z�h����K�Z��;��s�S&4�0����E��XB�(��,6����t�!�k��`�Q�����Z�Gp@�Jf�,�B,;�i����=���(h�KǤ�Bv3R[eAs�]o�3�}ģ@�NX���m�
�Bu�2i��1t�	s(��})�q�y&8`�3��
��)p�(^�¥�Y8`��P�4WV��3<��"mx�K(���<J�2��� v\pZ�]`�J8GbB�����2���u����bD��������O�q�{R���Vf�L�ذj�(Y���(�]���|�pI���2�YS�,RB��U�
65��煨�y;P�%
�t|O0Ը��5k�#f���5S<4��j�-yg7Xt�U{�Ɏ�� ����U���!%�,͢���3����O�ϋ�^�u���y���_�6Zw�Q���᷾��'�^�t�嗮=s�B:�����4��5�v.���Y	�i�j��g��QBF��`xL�g�\kq����[w��n��X�qj���Z��p��6|�Y@eb��_�f�����O�*ڻp�%�����axsd5o��/os�5o����GWTq������B�A��ԙ��1���>�����&N��[��Ŵx�������\��HY	Gx��m�cq}h��Baݧ$rP��I�8�	�%�I�Pi��i|�l�����i�3���𕲘�'qű��*P���/,�^ d4s?����~�F�x<��+�ں���tIM�t5��Ϣ�]��Է��lF�V���S\-�s�ԅL="8�I�;mbS��W6��AΤ���pk�'�����d!5��Wvj>�';�u�Cg������BT���^b�Z�I׷�}u��i���Ϭ\�Q5V�m�e���-:�z%��������h��LHL.t|�(t��J=,�]$|���:S�*��>�=y�$7��1�uiv�߲���,鷄�ht����^�A}�Z@� �@/��f=��&��b*��Y\�nw¦H4��2�� ����E��XYY�3&��Ug���~���$\A�"䥫����p��3#*J���s^O���&©&�ĈΏ���T���,���֬��dA�F,��IB��5��F��,`"�A���Q�~(5 Q
I4����Q��BC=���'x�	Mc�ˇ5hY�
B�)��f}fs����#]�I�`Qb����-^n�#qL��?��� o�z�2��fsO�5�D]m��A����~��W:�r�Q�L���9�?US�r��.f���z��{��:��aVL��0׬ʋ��*�id�����k����z�*sf�tl���޾�>�祥%Z���������O~��+A=pt�ײ]���@�QVu�Y�Xo�z��,�wj8�ϳ==�xu#�ѷx"�L�]?��(��-�ojV���;���y���is�5o���z���G���9'�A�+�3ၳp|��]���^��xI-j1�cX���9�}ϲ
K�1t�ױ��N�c[1�M;h�[|���{51�QR�~{���sL�S��s��\z6k,"�Ad6
/q��-m�(Ԛ�Bg� [$d�O&����*[�3�t�~	�/5�)׶����8vdIr�6�E�}�w�ˬ�҄�c��C�������� Jbu�a���+m%��М���t��:�F��(L�6"�S�8��cZ�QZ&��`�.�Ҁ�>!��/���lG�B�əZd2+����ۚӼ	_�#-G��d���B��&���T"�'���lnnn,,^8w~,��q����I�ۓW�~�d._���k��{�r�8r�8Ɩ�fj���7�|���;t�8����U���,A�%�����`h��d�),XA�'���nG�����3��)�ܹ=�,k����]�hi�ƅ �F�Q�Uz��(�De���~,�~|�w���}�*n�B���<��?��������J�=to�������K\���ǞL"Kn��-� ��莖��i|�G�?�yK� a��ivb'�2���wT���ӕ�iw����WU	T�E�����A?��pV|�DcWF��zj�n����^��z$�~t�j���F�e.�Դ,z�1%W:��Ua��'1�P��H�p��HDc�Xd"�* �͒�x.ɰ�@�5M~±�}��5	E}	T�qZ�*M�ı��*ߖY6�c�¦�4Y��}f�^HN��f�N��^1MF���J�_ Rr/��^����N�"M�ķ��џI��0h��d&a���ߢ��tDN�Q�L��n�����6�"B����1ݪ�9i.G���p�&b�����焦p̘�*�����"�)-�T�LL�*�9����%�D��-�Ӕ�^)��U��z0�Y
!� �,�'R����p��p0%\��rp)*�y*�d�N�Ѹ�������[����<G���G��ٵ�"�Z�������������!n��[��gίfDJ�����v��:wj���#���h��*�u#�}�p�G=[�s�g�aDX�5��|�U�B1`���[4���LP�J(��+�ꮍ��E�l�2�Ɖ��y��y���k�ۼ=E�ow��)�M�]����r�t���.�N�Ɍ�2�`�U��M]�-���]�=�ګǈniaii�ެ���<Bɷ�)�*@Qp�_˶�K�g���n��l���~Q���*Zj�����8H�:��Pf��1+��߰�O�%kCsM�溨F��H�~���t%��eW\�C�Є�����̞��GqZ�ϮɀX��B�x�`}pe2>⸁Q!g�:��3�JA�q���-���˗��E��s����v��������Ƶ��>}��������֪�R�R�F���]M�gpY=ֵV�>!`Ƭ�+�pʐ��t�X���=z�P����}���H��U5�4���U0�w�-2eAqvx�t���Z�p�{=V��}���b�0$!�<�\ccc#d�n�O���������D7����d�&��	�N�Eh�d�(����r�N����KWoM�t�~�����	V��:j���۷o�Q�n���:}nO
:�Q
�NctD�������f�������g��Ѵʙb]��C6�n)^�ё�ph�8@��c�>�ϊ|V�b1�^�T�����3��8Z-:nI��ha�t�t��Ѳ,�;�N��9Lm�q����(�����y�W:� �beD�t��@)��"ȷ���#�D�c�'�{ZҺЊL��q����n(xC !���cY���U<��h׋��~�1�*d�;�E�25խ2���k}u��U��gc�����t�:\VN��St'��?f'?�ϫ)��U�
�	p��:���ϩ�-�p�z)��4Jt<�8M�H�K�੔Yg�`�`�2#��j�z�K&�H�6uHS����Ѧ�Bod�4z�G`M�W����3k��ϝ�mMr��T��_\�xX��ߝ��M\�^jb��m��em���mޞ���	��B�y�:����-xL�i-�1�x����4Á`�0]�#!L�����M9�֡`Ah;���JF>��җ����px�/~������?�3e���ť���=���W������DY��l�qK�s2Y&Ya8R�������LS�6 ���e���t�ֆ+�4
��"�`<���FiA�A�Q�u��`KU &�fd�f��Pe�Y
���g0x���C�6�.t����\F(ԝ5ؿ�^ҵ��31l'/��Lw-��������-c�g�G&�T�Ij�&!�4��V6��" +ܞ2���]Kڦ�T��48�ɣ�j�}FȮ��2����0W;a@Vk� �'k:�^�Kc�����>YT{�1&/_{��w�~�O����������S+�k���/ȅ5R��~�P����w�x���C�t���]���{���.�[P~�\鸩t$m�dyo0�U����z���3�g>~�T�VF�e}q)���T�����2��#��X���G�ѵ��}���{�Tp�_�r�Ժ��d~fI���7Q��/��\���<����������������h�<�l�F$�����")h2����;��@�R�7���I��o^y������۬g�q�ڵ���[o�%�qX��uZ�9��������'~�Z���p�҅�W���u�]��]����Q���ҿ��{g���ի�`ZS�&d��tNeȠU'�����h~���l�X&E)��P��S��=.z�E�D��3�3ӱ���B�L�uJHӚy�x�݂�{�Nm����>��s�E:g,�A(<���"¢�Ν�Z`�,��^:j�s~��_�{�l�&�=sB2�'��Ǟ�r��~���V�����a�;�n������ܹ���կ���s#i��
=��Ç����7o~�;ߡ�q���B�o2�������Z`�2��p��x�e�@�qN����0#?�X��E�%����}L�c;^��-���0���^��w�s�*2�B,N��JVX��ȉvB�{��
|���,��l� �,�G��~��as���R��cs�2dͦP��e��N䀼Of�,�e�H�\�6Kxn,�t�>��6ͽ7�-brp�h4j����4�S��(��%?/NDaԃ�c9cÊ�xW���"�{��f���!w�=u�ԕ�S����>����_X>�����VP�,��fIe�t�$���x�Ƅx-ϱ=�v�B�L�����7���LA�Q�!M�*4\��t��y{�6_0�6oO��E�J����7�Nd����)��E�*0Vj��cǪ���_��Wذ�uP9oeEнi��f:w���=�łk���C��Af:E�N�a�e����П��SU���x�E�y��j���+�/= 3�2���h�$�Z��2�Z ��~`���7���tdIMY�ĴN{�UŮ/�~tK;��'.�%���������=�����|���w-�[����)Y	�V�9�b2�5p����L���4����ǣn�SG�@�W2�=Mz��?�Fƫ״��,6�k)����8�cq\h�G��s�l�;Ұ�~��T����NܩG�_2wY��A1}>A]�,��}d ������Ƌt�#������G\qggl�����G�f���;<��u,�vi`ɬב1�����w���N���~nF���=�}��s�cN6�����^�|y����\�35ei�����/^�bww����+�fm�mS��y���B����3��	����1y17f�R�3{Չ&~&�tx35-=!�9�!N�ju�EϞ��+1��n��8�`���`���d{O��@z�:4C�zCL�4��uA��M	H�e<¡�&�LtZ���h�P�f �I�Iώ;ݸ���a��)�[ �jR�&MT�V�5.Xy�ӚL1e24��}(G�L]�5��i��l{�_��`^婘Vl�V�Y��Z����&��Y
�ј||���<��y��b  ��IDAT�	r��d�"�0f��'�nJo�X��+_��`2>88�{���;��+1��p�A(�e����k��#�ÎȪ�����׮]K��F1�f++k艥h�[���~Ѕ�W�O����є�^�,���,����=a���uB���W��8fc:n<��Y���ۼ���k�ۼ�<͘��L�P,Kz���S1��T�'Ӛ�Zy�Q.��;i��JBT%�d=3�2Ǻ�$+��\M�N�_����FG=2s�tm��ZXY�Cw�h�(#�کQ�D�XR�$���EF6:�#o�:15��b���],�U�=���}�fp�L[��%��$��\9��]f���t��.�F1�--��
.���)�	�n@���2QSLy�Dի�J��_�r�|E�s�'B�kY����v�ҳϰ�H��Amb��K�Y�4�Z��do8,�5���~����"56��,���0Á�I�A�@��,�<M���>�!Sy�(L#���13!{�07�[�����d�;�~�ҕgL������%i[�,La�i���v��j������./n�x&�A`�K�rOc�ԥ��X�j�r��Y��Y�e6������M�I�D�r�1e���r`�d�?�ƃI�(�?zt���O��q�u���i�"�J[��n�,5�XX��#lK�,�~� ��?)v��ݿq7;:*iKuz�M�h���L�3��W���*�����h,#�!�CR�t���������[p�1��:닉L�YN�o����/]<���F���������Qs��3g������n�<�O���r��ۍVb�U�ޤ�Q~��6�T��H�X��z4���izx�}������E1
Btu�
Y\ҳm��s���Qo8��i��l�u��@R�9�i>�;���';��{NgѤ�t��r&I셁��ɨZE�-�[mP2�J��$��-�1����r��l��?�&�礎�;��6�E���Q��`=���t�"4P���!D�\�����\o�N�/ԃ�F�ݤ����Oң#��Р� ��T�k93��E�-ɴ1��䠱AlȦq-Q�86!UZe6��WÂg_���އ�\�%Ff��j�B�Oj�q"������Vc��4m��ޙ���3�g0�[�dK+pɜ_ns�- ��#��:���������Ǐ����x����j���1d�� N�-^��<払I���Hx^�4�w��e{e���iu7Zt���)a����h���N��u7N7���x�$�E��{^�Dvh]��t�=�)K߁�!N��Lb�UA3t}�L<�N7=b��mޞ�ͱּ��S����'�������[������[������_M!�9��V.U��&�q���h��t������2���������~鳟�ܭ[���_��<��3�o�~�����l�)���2Y�HXVF�FU��5���kL5�;��Ϛ��f�(�+��YI�v�k?.��am͸5G�R�m��G�.pe��(��s��	]]�߹���4�5��O+��9s�����ϵ�˻���7�˙��*pʊ�5�N�?<�2�l�RE��<���8�Q�J���
���h�s��d��:�}E���ZOݻw�|kiee��x���}�ß���?��5���b;� Bh�Õ�=�uk�ι��NO�v=��Ã(�k��������x�+Z��1%I�]���/�y�~���`t a��v���������
Ξ=���LiͲ4w�=B�:ujss��ի�_�h��M�rz�zH���]��ڬ磊4��t�� :Ù�s��}]�E��$��s:��ݻ�������*��+W��@D}��t=<�~����~0|o@��Jf\�pA�
ҍ�>}zx�z���,%˞{��h ���v��^x��7�y�:���E7B7��v�ܹC} ���>�1
�P�Xj��!�I�xXt�r���w�<��S���� ��<�Dz����_��_��\���}���lll���_�5���/�k-�@��J����~>Qojy���p=g<��F����}��C��b��_nv£���G�n޼��2������9#-O3���>��K:~Tc�[/t�B�CI���/�:�;��6���s�h>���b�TԻ���*���&��+�a��U��������9;�,�����-Y�Ϝ�UsLF*#G�u4'�^ň�z�SZ�Hp4��B��D�lՆȮ5s!�%��L̧O���6}B#���t��m����[���}�yki��I=�xؓr2�hUZ�]�4��W.�s�&́���G=��s/��0C+�9W�@g����q:>�i�������Emi�CW�FXV����΃������zQq�4�=f�5��Zn��y1o�6o��6�Z�6oO��=4��'�
�b���������������2�I,���Ye��k�0mC��P���}7y��c�f6v[�%�_�v���q�!�k���"NC��a��wL�bI�m��ÔD.b�^����;��Tr��� �*tU9-�༶�� ����8�Z��L����Lл���^�m\ȥ�4�F@�� 1���P�@M2�WℿUםÖ�mz�p�8#!�C0.W�l���%t,,R_�W2����T�5q�Aةw�y��A�da�,5���K�I��"3|(�jf�W�9�S��FýGq�Rz6�Ŧ���5���Щ7|�w��<�s{�c��#2��Hn��zcDI�ޤS$���a�Uw{=��ؼ^��6�YU	L��`�;&���e�eO?0����n�kQ�'�h~Y�UG���5��b{q�m��n�V�t��N I�(����M2�6��4�G��9���|U��Wf�J��^ZąʜI٩�	�$�qg�F�`���7I&�o<k��4}\�X��w�Ih[(�Y����/��?4g3�kNaH�,z��t�P��ho�}�P�W_Zk�Z���Ngq!+�3g;K�6Ȃ<ُ{�]�L�	��Sx���S���������p��Cc��NeM�)WO94��Bz�	^p�)j7?
1��
�GsW*��aV�!B�e���RI��u[	{?4\S�nn���3��d晅S�vM��pk畫�L�[^��wv��<tjk��7��:�ہF��L�N�w�t|R&4M6�4֩3��N��FШE��ڲ�y~���J��Y�Ag��kk�-;���������:�vK.%M�lN0��4���$H~�pǵ��B� +�;1sH�A\٘�L��cITH��kgȥ4!�9�r*,�z�'�	nI���$��ᦟ�B\'*�OL������)���&6�S�{�{I[
l�*?P�a�Y{��齥��N�@P�d�+4��&���hE���%���N����+�S��Үg�jX���,�_TK�9$��������tZ~��w�d`[a#t܀��i��ŕU��~��4�� 52�k�i#�؃V�NG�iZ�f^84i��ʍ���8���a"z]ȇ���v��:�]��f�<�5o���m���mޞ��P�Q#���YV�tx���r��������~Jch�j-���y/������HҨ�1t����[o�����?񙏢�co�~�ۿ��GGG�����`ּU�TaF���<��Y[��l��"S'����P��q\�@?��P�T���kv4}�k_[ZZ"�I1�"}B�Sߢ��\�Rd
p�k�+��V�r�b�W��T�Zd�b5�d���u�vLMk-tn*S�������ݒ�X���kB�:��x�֭[g�_>}���O'������L��9�ƞ~Μ4��c-}�dy2�����1�,WY[;��W��U��q�����}�s���߿�����я~D�,��L(	-����E?�o�+y;�����Xm -�D��(����,��ݻ��ܳkkk4OP���d�Cڸ(.^��ꫯ�w�~��
gD�m�H���ݥk-_�<{����s�=��y��t�nH�ԕ�&�bd�����F`0(h�v-��ݻ�ѭѥu-MNߣo����+o߿u�ҥ[�Gt�����g !d���d������|����Z�G�s�}���J:�}��7o�ͽ� ���ع��^�-}H#>�я�4����&���x�,/�3x�	�ʦG� $ل's*1��Ă5��Ȣ��T��'�:U�����h�ut�~��������UhV\�v�>��?�C�ʯ��W�H���{�x&h䥼v�<��y]��>ZJ�ёtS.\����-��|饗����G��o��6=2M�N����[��[�Zc<Ӵ'����,��rt�\�<	.e�Ci`RX[At���oR21&�s]�9��$猿J���A(]6����&��/$'�9ZBJo��rS}�l#�Q/NN�1�M&��Ξ��o�t4a�>3��jY�kJa?�Л� 41���V�\J}�����2����������,�'W?�"=���5��_��W调[4�<�O;L�J�y*Z�(����a�F��3Z5�;���ooM� ��1aFx/�ѲM�Lg���aXC�a�
�*�w�z�ơ�d�Y�� �&P(��f
֢b{1@�x�1�N <���T�ۼ�ۿ�ͱּ��S4%���t��z�*!�T�WJ��)`T]��g�kz=.��T�d��Қ�V0��,��A��,Ӏ���p�<c�D�����d��G�p`<y|�<��8I+)m��	+�Q9�(.+�c�i
���О[1E\:�1�'���c��K��'���T��<��߭�M�ɓ'�T��q�1*G&d���u�=�U��
�I(80PYQ�x�%x�v�z���9�dU��ch!-z� Hde��¶e��,���I�^'�d�l2t�w6`i��u�-�d��Z #���6��fXr�9l�21ё<�>�ئ�3/8+ؘ`~�2���T^��`�{�aۉ��
Ĺ���xԯ?�y��g�6;�F"�}ñ�B�Y~V9�LJYO/�GQqp �9��d42SPH�b�qux��ʳ$f�Nm���H�����z���&��rG�,
��;:�^?�f��DurAO�mC@)$�������n���Z���d�G���V�/+���8��'ʆk�����,�	B�V�6+��2�]%ʶ�¦I�!��/.�{�k��;J�`��ƃ04')�+S�e��p����R:��Ԇ�e`�,鏭l��;[��XZ[/��d��hz�m�B��&�xh%�~��k���:���A��l��Q(��4r�� �󂦣������*H���K��������԰���I��Ks�v[�� #ꆋtJc��Y���i:ePk������a�ܻ}�S��,���hW�L�����K'I*Q�GHf��y;ah9������:�⒑��h���d����GS�oԖ��iU�{� H)I�4�҂��8�w�YV��-�߆锡+'��^�@Ѿ!t����Gہ$$P�U?�uZM�Zo7O�z��vA�D�SI� �_��^�W4�Qy�ГQ�H��r\a��q�T��C�#L�ũuf�8�G<�ݚ�?8Vy[Ϙ�^�!uV������B�Ҫ|Lb�2���j%qR�c�Ӭ:}u�J�a��Z���Ч6ʵ��s����v2];w����t��,��&c)�L���'qL����t����Q�t��T�m�>r"��>� 
f�͋2�˵�)����.PqF'gX�Q;n� �Q��b�=:8�Z^	|��`�Fꌣ��_'q��Kp�q��y��f�c�y���h�43F��ݚqc��BØ�R��dY'x�a��b�����ۚs򇊉�U�t���舎o�;�����������l-�4M�ͭ��Q�L���Tc��b�siL�)mWuMUU%���*���Y2�X������o�a{�F�$;�p8��SA�rL'^��r&�e��gf�3!b5/�¬nZBP�UA���眦���Wh�$�}vҫ,�e5�u{�u{ee�,PĠ��Z��L^\E�P�`0�t����.�6f��b�k"XqKZ�7Q��m|R�&�{��ޛo�Y�0���mfP�u�ֽۏ��=�J0m�&�laa�,6��������o޼�m��(��sDJɀvl�G��oG�P�5)���h_^�vqQ��ײ,�"!^2��!�E�D��4��8�O�#c��Ri��H؋N�E=9ƍ7�T>|�0�-ㆮ�](�枍J�q��,%�E�2 4���х.dV�y������/�@��ؠ�]�@���fڞF��a���K/v��Ӗ�����*�]�,t����ٳ�������_���ʙ3h��Ӎ4�����z��4W6�Ѐ8�85�K'������I���d%n��B\єJ�����8�W"@i8-//���+��qQ�����K���k����l��"�җ�D`�ƹˑ�jڞ^6-�}N���7�N�_�*8Y�[[[t��]Aҵa9����h�����ַ^}�U]ΤCv4�q��fT���i���L6-Φ�@�� QF�tmQ&��!�����W��LN��:z��D�X���a�(��	�M')����\Hvr�g{�q�$Str0����=WG�,�ry:�8{��V��a�?�~��-?8�vG��k�)Ϙ�Q�f���5˜��#�;wo�ϯ���S�V��B�8��s����r{���&�>�ysN�c_��a3X�K�SH1���E�p��i�[�u	�=#*N�]˵��iN���BX�4c��4���#��x�]�@���;�����|���m�~�6�Z�6oO� ��+�Hz/J�,2*�,-e��#���~T	�S�
�{�LJ�)������6#7f�k
���-�,�'��	K247l�%�R&I���uP6��Ā2)����@�S�ʴL'Q��*/�2,״J.���Q/eU�u\{fH�,�����a�Y��d_�2/%����.?��t�W�pQ�n����n�qQ P�-�
�n�ʒk�l[WO���8J� mP2G�S��-Ii2/>ݵ�@�P�-%̾�u�I��NR�U��(��z�Q7��k��J&�_��J#cҰؖ&���p�YC�~6�G<O	��@Z��X��+�:�2z�Y	f��0z���dK��q�a��0������'̱Xo��?��d�6�� -�lB�*v��Q�1�n�
�p"�"K}i{��PO
j>��dW�a�.RG�)B.�󢹴��0/�������YZJ��D9����{�XK��J�s������&�U%K*�HI�Z�H0H�!X��[?����WpȰa� 7�0�ې���4��HZ"%R�!kbUeVΙo~w�9���;"��*��2�y�J�7�q�'��k������v=�gP�3S��A��M�E}'���������1vNX*I�FN^Z_� �5���bF��`R>�H�ҵ�upq�𘹲���[.'������h�,=m�����F��z�}���{1��l���,�$��{9���'nfM�Vۿ�=�J�mE��Z�b�ױ"Ē'Gg�>��F~Dk�`�>�I����e�����SG���	
�.�xց�f�(/r(�T�k�Yѽ�#m��J�^(�{^�"���F7��G�Bq�����4�b�3O�س�<����
O5�.�!���lJw� ���Þd9"Q�Q���oS;%X���p��"��5�:`����������/G!����Cj��Um�Φ`�il�����O/.���x�s�-�u�R%4�to��9���QIF=a�*��]��]�^Y	�a�\��	�?	Ga������U`q�m�h� �0��%$I�U�� u���r[W�P}�τ�tf˱G��Ʋ<QՀ"e�:"�)ėp��A�4�h�hj؊����7H�]��V6�����%�nI�A�#���zV{��Y��&��u�>��E!�����}덷���\,�I�iz|��8^�̍�{�a}�t����#�������֨W9!��7���z\���������/h`����t�x:G�C�d��O��5$S�J��<�L�d�ki���<jz�*Ƃ�߭K�"thX�w�� %!s6��+�k�V퇷�Z�U��qs��l�xvS����c���_h��a����X��;AI�L&R*GR��H� ���@@"13 Jh(o��׹��P��̴�^_Y
�cd�`-V\, ���c�2u��Y����rU\*ЬH����<,D!���	[O��]��_{~7�˲ͦ�)��7,ڈ��,eó�6\�d�.��H!�>�woߎ�x�5\�wL8���̑�GJڲ!��U *hm�y�O�s$��s�X�n�N����O�'�@�rl�p��xA}k2R��v�Zv�F�An������ni��dLf"��U�J��F#z?+`�F�p2����2��k!��t�������(���$D%(�Vr�$cg8�������ۃ_��_;��mT���cB�;f��@�Ę8" {���<%P�QC�����j�7Ql�޺5O�,y�[t��5���x0�XͲ�˄z�5�����OY��[��n]�Mq+]����������$����/�P��Z�͢�#����ͻﾻ��-��z�{�.I ��|H[s)[FPU]��]��ʔ��d��սue;�І�!�K3gz����<����;��{�Y�M�R��_��;w��b���F#&K,	�I5�#���ww
��޹I�
Ѵ}�
��{>�RdQ�z��/�L�����Ә����76�tz������1
����-�nX�/��X����J��,d!N��}8LB/�����(���u7l��6��9Wq>�Xb��z�A^�������Y9���bv��#'�Zޱu��8��d]��a#m�����Z~
t	`�mҋ.Ш�r�l	K��*�/���x<~��i|��k_��'?�ď#g�nsZ��M��`��k�����6�����:�?y� �:@�����m�$�K�ߒ�5,BN�Gv 낻��|�;�M_��Z���X;����3�V��j���֪�ڇk�G!}hC�&��n�<A7]w�M�%Hf�x3u��V���v Abc��2B<���رu���;�Β�F����*��u�(�#S`8
����|�uu�&[<��*K�,e�k.K4<���,�[�\.�lJ��`Zj��ց�ֆ�(f����׺�FM�.lm�طD+ݿ� I���>u�|XU������>g�u�Q~�2�gQ  I��<��]�\�K�I�r��D6,��������<��3���[l�Jt�$]��|�@V-\�K0���P䈌r�B9�<5
q\�q
|	<�)jS;4���hms� ��u���$�O�1B�ɴOV���.��S�[�`1_�2�����0I˓�߀����=���"���,���B6V��1�*}�������"�z�o�qJhN��������c���O&o��,{��a\2��*�T\�I�������6���_G௘-�7www�7������l��}4?���{-=�5a�>��A��8�0����d�^x�2"�:=GN��h��:I]���E�w����<���{q�E�������������ϗ}5�fI��o�R�.G#Zh�_�FmK�'76?��>|��wL޺��y�c�X=Ͷ��j��ܝ��E�A�̤�:����i�E�hn�Z]!wh�R���f��� 4e^��QV[��Q�sj�QË{�[�^{������[�T����G>�o��]��ޞs=��?=z� 5��gO?})�P����Z� �1����l2	<s�:ޗ��o��?�'�{[����G3�t��/_�J�2��+H�����eY2��B�S�29���|���}�*C����붯q=�i��]�rp�Q�L�2�T��j]�����m*T�&�@EB:�,*�����-D��F	R�\�܌f��JA��n|[�Q�[Hł1]"K*G�R�.JY�X�Ii�%7�0vλsX)���ʌ���B�|���w� &Ӝa���}u8Z/�����_}������^x��?u��aV�~� �X���_�ݒf0���������1�~}ڨY�%�Y:/�֓��io�z;����ӻ�i%`o���"�=+�ʱ7����6�@n-�M
^�p>��C�R�pY��p�ls�+�U[���m��Vm�>D� y��T=��ģ����s_���er�I���;���^�C�������^pC� L=OI{�:r�X%�ef	��9}Q�qM���Ng�ٕZa�xV���ݠ��6QC�T�jH��x!��N���}*��gĜ��3>�_�aOH0�F׭X�(�9RS��w�B��c^"IBk9�����<�z_�-��ș��Q����e��Bq*V�qF�g�46Yko��vD$:@ߜ�5��IC�P���@���$M����k��"�E#�h2��M��Q�O������F����p^g�6�;��sƕj�*�	��p�d�,���I�p��43���/�#�;�!�g���akkk2�P7������8�-��Y��c���q͹���71�"sz�t��nܸ1��_U�����=���|>�qtC� �۽���4��KC$*�X9Q_��K��F����Ϋ��G�A- -S���]��E�'���2��,�X�E���>~Sb-}�|��HT{���M=� �1uA��$�d��t��N���� �>^��z�/�?a���i~:�)XD��yX���)��~��O����.�Ͽ@�귿IoR��Ƥ���P�� �>�Q�0Dj]u;�ۣ��3(LZ�2t9��Y^}�U�ι5��dBX�g��ŉ���}Q8��a���+_���|�.�N3�:�i��&a 1�8W�s�9��3sդHi_ndF�$��:W��ɗ��RW�_d��jdH��u����nk�	�N�i�w{E��^��bm�
ɧ������>,�z"�aCfʭ�+t4�M�����X��.�q��a`�M�i}���������ʗ����y�����߾y�&}�sn����C�+�V��դ(�
|�+:��]{�!��V��Fy� ;7�����8��	���QP\l)�V�<�z	kv�j�Vm�>L[a�U[��Y����_E�M]�V�M�����L��k<,�..���NC��j;�-=�Lk�)�����ͽ�`dj���sԘ�(�T�=Z+���ȅ�Gq���_~�#![��<������񄾓����Q[)�!��d�-���|~�lCH���3l<Y��*�	�^� �)=ϑr��._&�X
���̲P,6���c� V��V��6A�bx� �y�s�Q@��E�z�msHn(	���ī�Q��D�� �N���^X��;�2E��؋�X���8S���Cϓ�R�o3ϋ�\�Mr�皓m*�Z5�0�}_e����F3S-�Y��d�M�@�^g`����5eE�����7�f�Їa�UI�y*YL�V]$줐����N*�'�YRjBK�׋uR�K;���i	��,��}G�<TD%���`uD>5M{�`� �Le��hh��+G2�<�z=7���S'K���V�Ȩ�t�؍F��ü�V�����a���f?
&Ev:�Y���4i/��5Z���o*��t��Q���w���|� �cO��tƏ���	�o}�;��dS�nx�訿���x\�U\ƿ��K����>8��QO������ank�:�ɔ�Ϳ��6O3U��4�*/l��nI�$?;F�����Y�2�j�"̌V2�Wk_n[$q&�g�r�\@<?#�S-,1��]����T�@����_�Kߺ��4��|��w�޵g�4<�mąZ���o�{���{�I��%S��u]�?�;;���nѭ4�"���
��~��_����v77�A��;�ܼ���>�i��G����{��t�ɟz�kOB#��GQ_޼��?��Pڈ��k��&����D`�[�0T��?�.t]�\"Ԡb��lVp�ewPS�B6-1��Ē��;��Ƭ7��t[�v��H�v)(`�}H����v��T'����4���mS��v!����[;���*��-�=[��]��y��{C�e����];�q��i�(�i��cfyyቫU�����������n8�;������᭻�v���эI[���p��U"������~XiU[:j^g'ɤ�U�ֳ*Y�L�"����.0�>�y���-�:�]k\���:1�xdJW���.z`��ꤶN%��+-*Q�J@�Ҽ+�k�V퇵�Z�U��Zc4�BP
n����y��jI&��	�����>mm�s]
���P�B�JU���\I ^ɩr.q#��-�8�O�g|z:↼��'��#�clU
�a�=�d1�6GKB�E��iڹ��F	��\g75�X&.����)���6�|�2b���8MMD����Lw%#Ŷ89^�D���&YPF��S���(��/��r��^�W.\��`)3��ц>�ħ_Ee����_�>�w��1%d��K�a.Kx��������	Y�q�,��QV,��m�F ��,��ܔ|��ل&��'f���x��ȍ	8]H�Pm��eG�#��z� f��G���&���k�+��[GP�X_���i�z\�z=��.&�7n\,�wvv�<?==�
!I +�4;88pXpm}4�~pt�L�P���A�jZ!G-�KƷ,N���9��x��UZH+T���U�84b�kCE��~���qo�� ���/R��-z��Q�-�4G��]�f�v|||vv�ۿ��^di$Oߺ!ii(�4���"�g�I�03c�h��E�rimϒjo2� E)�K�f�?Ń �w�6��DU������Ϡ�h�T�u�(766h���G������|d�����,C6�'?�������1�p_��\��ŋ�Хq@����g�~�biФ�H�F1ᷓ�������]�F �֭[3��H�G_��R�i�����?���k�XcyAk���l�/~�tu�n���������4V�ӱ�J����x�'����"�4τ��
��,�A�����u ��0�Z�.�Sx0��}XK�Ǩ'�j�
�u���\�P&"�ŭԅ�G��-�F�q%��k�N62���]_Ok�w��>��&xWZ�������4�J#�r4t/]�d�	�$O�FE��� ���!8y������.��n�Md��U��~�^�̦S
�7GMs7�p7�4�x���'�����&lR��Z���&�K�ڪ�ڇi+��j��!���İ����E�-�IJ�����|�Y@��� ܪ��k���o���n��ocOq!Ny��sܚ� �X��D�J���2�#߱�^T�"3:���}�k��uК�
��I2�\76��B��9���~_��������0��rb�V�
���^8F���Ѯ��`�5bkYο��&�,�&y��aV��d�OU�j����@^956KX:r�t�G���"�]^�z���wC�u�C��am��޺{/?8���q`��o���Q�������h�&�O�^�\���P׫C7�r�%�޼�
�W��l�P�66���x�Z�S>����L)r֍+$OT\��&H� �f�Z�M���jf����{����!b7i�N칁ߏ��G���ŬoT��J<9��`jl�rj�]��3sэ6���S�F�ڃ�<O�E/w��%����C2��^}(���ί\�RV���S��L�X%dÚ�����Ӽ�d�������ަ
m���ՍK�{�m(m����#GWa�ѻs���^0 �Qd��d��i%.洬�t�Í�{h���e�VY]�j��g��*\����{A� �j���E��a	 �.��ٲ*�F�s�~?0VB��y��b'�R'�Bx���&��,�YIe���izB�����T�<8� ���x�#k����9�P��m^f��4W��>�
%H>�I_�/��r<����믝�xH7<��4�c����;����,{8>MtI�t�&uY�b��j���r�+o#��֪��g>�__�7��߄���������k�C���*��?�����՟�	J����W����9�l6{�ҳ��o~���"Y��v����lB+5]�~ ��.���N�N-Ռ��ڨ�sX�ޘ�<�	�9�[ʖ�)Ո�K��,�8�@�s
밳Nc`�ut��k-��+�]K����v3n�@�h����ڹ���Q���(��<G���O~S��'C�ۘL�hIҧ?��O<x���;;;A�hli�����z�����}/ti37�tA��0U&��L;���O�Wt�)�:�F����R��&yr��t��ɟZ�^�s����� v�R��@�6:���(�� ��Z{x��sײ�����h+-�2Blמ�'�k�&.����c*���j�ֵ�Z�U�Ͷ-U|҅��F�<��vN��xB���翝oU�9��C�6fGw��q$Ӈ�Zr�SHš�U�� ���yD�Bܙ.���u��r��,A�U!@��z��:c�u��?0R�s�r���$f�4��g���]	�<u	�Ԏ�������k'����ʪ8o�*��aUY�$ �!��xxxX�	g� ��v����3U�h,��8���wXM�R��3������˦�Sz��!�"���z�ͭ��=:�9���p�%Ƽ�Z��3�yY���և��|�Hf Je�J�b�-�L`)���WM1���bJ�h�I�\���@s��=bR<�i~C�������Y�c٫M��s�":~h`(O����(�C0iu=������<h⅑�Ω�"P�����,T��ZЦs����	�ooo�C�ڵk/>���;o"�,��ކN�����
:�V�kL�� �
�fM*2�Y�`��	����d�M)d�`�n�V2s0�y�+-3)��(�^��b�`)˲��1j�3Q�>'��{���)��2%ұa��X�ZR ��i����ᜮ�5W����K�|����ٻ�Z�a��o���`�dB���666�
�;&</[Gǧծ���|k���彟����W�����������o� pH�����h�ґ����,�5�~Ҡ������Z9�)�JI�)������ W<��ʢ��'2r�B�w���Y�oVv9��e�雁��%ae$;�j������r�n^ĉS�J�˼�0�rF�[�m������6ވ�b���/��� ���MU8pz-SF�L&��w|Eׯ_��'	k�\���t�M-x�D�����zq ���c�k��j��B��2]t�٦��Vݪ����0)���|��EU�ﺚA��j���j���K[a�U[��5@H
-q�?�򂫯4~�_��be����8g��GW���_�\��=����pgdt�jI�Vpj�u�Q�D�B"�ل@{�U�pVEU���C�����M��5s���A��C���0��s�sX.�)j�85A;�YLV�YޒT��2�M�
�t��Y��ی����`@��mKM4dU�V��r�V�D�Q��y�Pi��ݨ���akG �r�+�@K

��7.�P�Q���7��d˄�۫�f��}'�`3�  �22��� 1���>�~�_H�º�ɣ��x>�N�:s	����mE/�54�C�a��[=�䰞��.]C]�t8��2�S��]���TYo�Ü!��B�W��T���J;:,�rd`�����7.<��<?.��	fE��j]��yj]6�Ҳ��L���_����%ɼD�݇n��ķ�u>�zqP�-��d��s� t�+߉������B�2�ɨ4_'��8��L�����d�f�ȇ���Hq�$�[x�Ј�X��]D>uvs�YX��-jD����.� �)��F�}39���7?Ɉ��E4�<8�Q^M�6%;��^�rx�k LS���)k��wsU~`穢�<D��&�1��Y��J��ӵ�%��da�5�p� �+��)n\��V��P���Z�$�J�pq������n�IX�tՓ}&ɓ+W�\�r1����x^.��}WU2�ga���]���������x�?ӎ�������~t��pG�OMG8:9��h48>>�.P�5�>���~�8ӓ��L	��|�GS��SW/T;:���z>���Èi��Y$jk3�6�Z�]�4�b�.W�c�]w��j}U�������R��i�K���y]��mwWyQ�:݉�~̕ӹ��)�4NS�c��vn�����㹦Ȋ,�k��Oʑ��ǩ��ݮQ<����m�^�����~�>�QӰ��g􅻏����s���*���J�ʩ�1�9p~DWmC�+�Өe�f?+z�����iK��ѝ���̞�鎥��_��n3��N��W)	���X~V �w�����T�_ŅiGCY3�*���ҵlX�j��j?���֪�ڇh�P9g�:��N���y�ǙW%(�q���:r�q�r�as��� ��A�J|��M���$��z*K�D�3Rb3F�GX�Cp �m\�ld¦/�j"�XN�π�*G<����.Q���R��m��>0b���-�gL��fV

�|��j�v��̡�KZ�H�b�R�UJkg�o�<��T	�h�'8��3Q�����k��C��"�c"~z+R�џ"�&rc������^sr.6�X��㩤�����KF��ɉ{e�W^qSw>�{w��&�"�9O�+�^�cQLj�jKL��|'k��TȾ�0��t:%����&�����i��~�_M3��#v�͡I_�>\}�
t��W�}�#���7�>�^������������_���FӽmrY6QA�MI���f�! .��`�K���]����������\���W�)���m�!�Ae���¬��Ӡ�t.t�j� 3I�s=V�P��F�X D���21v%�v ����ms���4�q�^#5^�"ʗ�P7����ˉ�(R���,��nޖ[hXW^E��[�M��6�)֙���g>���_��_�����o�ǿ�������_�v�g���H.\�)�3��? /�"�RZ�E]Z���ѣ�%����P�!�Eב��>�Nn����E�&0�a��� �cYЯ�9�K���ΠM#~X�jh�3(�_�%9��(ad��ڜ���Mo�����\)��g#��kT����F�CCA��Ce�z�橖��ԣDJf�DM:YA�(8� �Bb?�y�A�/փ܃,���� �vωP�L���Q��cX8�����bF���~�	K�l_�>}�{�7����_��7�O�\����F#bj�Z��=1Ӝ�9�AHV
u��'���3I�T,#ٹ�4o�H���b!��hqm��=ǫ��z�x�4w{�
Y�ڪ}���Z��j��S�((6(��B�?z��V�0`a�+^�Z����d%�a%�{��?ݍ>7\���_�b}d���!s��֮�B��8�;xs�D��EZ���ت�6��`ap
����Le9�&E���,��J�l�8~`\���j�
���]��j����[����[]��8oT��3�������k�4� 2$\$GB�F:2�,��W�� aG"�D�ʃy��
j���|��(�M��&�[gִ5���R�#r���Yΐ#��3#�f��U9�׶.3K'X��WSiT�@U0_�r]�y���>2v@yx�d�xs�|�S/ϐ�S��0_*k-��f�d�k�0���R�}c!]nTP �)d���O>����Ri{��{uRe�^�����P�=�i����T���\8��ܼ��\�*�k�?���.^�L��;;9Y�&;�Ƒ���t�6�C�W=.C���N��VXs��nR̼\���9�j�f�l��ޣ�'��LM�`<�L��nE�D�I�����0SO��uQ� �	*�P��n�{9dkhaӸ�t/X���𔓣|��9��]ch��J�lv'��֏�&�s2@=+����;��f�Jd��b|�%T4 n�X���%�,t��%�]�D�������~���/?y��ǞIl�yq��>О�낞�{W�~���@Fb����cW/\X�2��d1֧��|�"M��F��iZ][�ml��̳�;[��ܽ{w�o]��ZL'Q����|�Hk�(��G���$�&�y�(��L��E�В��g?�b�[c
�����2�e��EmY�7�
_�7E��n��5�?;��Z�?J�'��8��lv�Ti�m�J�1�_�k[�Щv���6ì�}�p�j�`��2Jq�Ū��f^feQ��>�d���cҾ.�?�����{W�߃���7o޼����'g���^��<�m
l��*��.!�o*]U!5\nʱemt����i~��F��\d�,kژR����1�:�ȼ���f9GX��w�n�?����N����K�i!Sj��ǵժ�ڪ����Z��j�Y)��M]�GJe���ɊpFHδ��<�YCK6��k�HU���[w煬�<�����h�GE�K4���Q_!���8��e5� <?���i`�h �f��d1����x�D݄y��(��i�t9�鷚`Hp
��*vN����=ϑp��Z��Z0�H v#�$��sv�i�w����y��h`̰o��^9,U�Ȫf���VCC ����sJF�Y� �;��焮�1¥���<>����V�j^2`	Ӂ���,�b7�K<+b�N#Gߕ5t��tl@�ܣa�;��kpYj8�o�*��%�/�pU�@ߥo޾}�^o��>ll(�L��f���gfI��w�bZ�� �����y��->�Niɝ�������ڕ+�k�9��g��ȍ�nYC��fcP%9x��
�U��1�d��nF��X,�������]�� �J��������t��ڀD6�'�
zyUJ�*��mha,�,t �㨇�i�P�N���!�r�70��ň��xM4ol&7�i�?�Ë���Ϲ�G��4�G�'��˿�K��K4���x�������S��7�9�6=�8�!�~F#�u��=oQD\���hcc���>��>��;���k�E�����論��{�}������{�:y�������O�����g��;;;�nܼt��W���$�EQ2O�hei��R畩��8W-�}�/����
�7� E��1��ܗLD���y�\&>��)��p��K��^���6�v>��%���n�Ȟs.���`j�Wz����$��q�	v�(-�wD�>g�����O>��+?��h�ޝ�/^̓�_��_���oRg�{}T�r�t�J�(�*��	g�q2f�]4��B�t2�xs�2N�I�$�~���f�<�J�L?���j��}�Տ��<�Vm�V�Gl+��j������$O�e(���d+<f0T�k���8ֹG��,��}�=�$&DsHO�m	>�Q�� �����z���"�<uG�F|YY5����c�wXңx��.¸�+Z$H�
�&C���oĎ�쎄�۞�!�%A�i�&�D+�X:h�9b�ŝ�aH�����Έ�]��M�$�l<k��h� @�@����k�l��3��ʁ~��mZFNd+^�jrS\F�����*嘢,�:��(�d�F����R%�a9����� ���T�<� :������z�c+�5����e� "2t��q�:�K��"�R��}�� ״t <��[
L�E��:B�Ԩ��Ne���t2/tB�d�Β2�aD�f�(��Ql]�J/J3�	��8dl���"8ڧy���- ��c=�V����d�*u�$4��ݭ\��K�FS���������F{7����{�*ٚ����/�q~rrB��7�Y��_�2H�V��H�޽���_����P�֪��xf� ��|���Q��|P7*Y	��h����jH�q���:�Y)�2��G��jG.�1a�9_(��hTY����u�k�q-B~8�N����uuv�6z儎]H�̰�V����"�Y��iʾb-�Z�i��@��Ҏ�iz�@;�t�������{4>�Gǳ����>�oYB��s��v�!���эΖ�}tR�派b�E�������^Y,�g�H������A6ϋ��͛��O�����]u:�f�����z���������ݛ�����.q�.֡�A���/�h��N.���rm=�P�AYt�����n}%Kȧ�%��ĴI��xf��yM�"<4��'\���/í-�޹�:h$��ZJ��z�n��K�;���9"B�ţ�Z�ɰ�:s[�J����(��B����1��eTD��$OF��=���[���kq�N�`��U�����m�Z��%y��A�-b��u���z=k��h-g���<b���x�~o��=�R�i����ioGz�[�Oh�1>N��i�
�Ր�D��Z5����;vs�Vm�>�VXk�V�C�������B<=B�/�������x�6ρ-���f;�҅͐aJ6�d6�w^}�U�`�'�x/{���ݻ�ٻd�H2ze�Iy�W�"�#�z��N����u2����JfY���B�3əw�<�Eh��J\K*d�����?��C�E!v���~D���,��<ȇ=�u��	����+ø��i���S���}���[��$��8����R%	�4N�K�^^ �"�����?�Ǆ�_��p����`�P�Z��I��1��#���E� $�%��0k.y]*���C�f'�l[��AH��,B�֩���s�Ic,Ѱ�]�1���	�hc�I��\#��9��U�F�Ji�w��]��ᐰ�a-ZQ���O�����G���@ZA�����VO�Q��ho=x��\ڢ�߸q�z����)�������<f�Ga-���j����|����7�#|��ﵝ=:�����}w��*�{˶1]��]�����
�7�i��B�=Mõ�5�����ͻ�����ӝ����̓O|��������$B��R;ۊ�j�nT��U˙-J������A����,�*�O�Ɠ#��m����fY�4z�=b��F����!����caԑ0w]%	�^m�ay�$Ihi�
ڏ*�阄f�_���W����i�h:������i^W����Z���l��g����[�n�u%��
�k ?�ܹu�6� (���|6^��n �!�L��WP��������Ǵ��a���7�nt������F��z��6"Ө��n^���2cS����@WZ����e�e8��c��cnt7�-gu������.��s���i��%����=z��������qpP���C E����)}�⾞��3�a��(�r9;�ὲ����=0�a��#Yp�8�
�/!䑯������Ff͕:���r�b+���"[��j?r[a�U[��쒛VI��Ě������c�y���a-��y�ߞ(��Н��C�&	9[}��e�%}�H�O^��#���;�Q9��\/���BL=j`5�H� �`{sc|z2�g0(]O���p��È�C� Ⱦ�h���^�Fi۔��`�r@7C��y�|��Ja+]l�&z.�do�C:7!����h�j82��Y��Q��9�G8.6	<�	6p`_���m�Q�����E���K��j	k哅UBΕ	 _��ځ�`mj͉yi��_�c	!���E��ǂ n�j"���.�l4��v���#Ao�~�z(��(Җ�b8D
�
1s�\���P��i�������%MVRI�TP�֎���u��&�R�D�ʝ�L�Z2�2rM���=<��\B�f��
�iU�Wj:��˞Z�,G�Wβ���O����A6�v2���tл}���E:��n�u6XO�ԾaQ�r���F��\uML�����ׂ؉�GӳܘA����DB1����$K0r����k����c��KZ��w˅����@nh��YS�7��92������K�Z���3O^{���4���3�tlޛ�]W9!�r~V\�\��q���>��|�36��\����*Ms[X��F&";��Pw�C�أǝ����]��Q+��y����'��F��á�%G��&��s%��eV�˦)�-����7��dJ?,T=�'�B3g�'dRA,�s��+��AS�d��0��ZZ����rZ�$���/^z���|2�MgLr�^�(��Z��X�E n��R>�7�P5�e!.��t�45�X\�=,���6������Y5Kꂂ����7g�h��au��z�ΒGC �\N�і~u.D��%j4`��K���~��j� [����{���.]2F�o�Pg�΋tcg��#? �ָ�5Xz~6����ǵG׬t@7o�WyQWH�|!���蝢��)+ϡ�U��t�T��ϛ��4�LF�e�R�M�j�s�+��0~6��8Hy��E�(��B$�sL�x��ڪ�Z�VXk�V�C����P�mS#Y\�qidrU�w������[g,�I�3�#ۅ��.\���r}x:/����߿t�����E_	E#լ+��A��Bj���涹�yvv�t�AT� ZU I���q|�+}m#vڲ����2��u-�?��lVBD���k�dI!��RF��6�ˊ�{�4n��N�D���M�c�%n�֝�����*:�Dh ر+Tc�u�6��(��5sA3Td�
ǅ�X1Vtw]�I��E���m�.փ�%N��wlW(g�
�pJ"?�`����
Xc2�c]��i��'ΟwSFΝ*03􏏏0$�p�%�7�[��i*�ܑL*��"�����8�A̪z��?wg�~���p��zt�7n�u6AI?�u��j�Ar8i�}��n�
[����%39Us������;::Z%�Y�͋/���I�I�ԗ�f��LμRL�x����O766v�=��n��V��G���`p���d�(��&~�ш.���f59=��rr�b��h�LG2������k�;*^�q���)+r0K284��QІ���d�[J�;͹yhtc"�)c��/Y�	�A�R�7�p����Us�F�@����裲�\x��OY�NT�|���B���J�b��ӊᴛ�jc��J�Ӌ��R�}W�,�J���B])Ѻ2`�� �̅
��i?eu;g祲-*���Y��Zίk�u\/�E?��Y�oȈ�\� ?��aЗpGl�<�3�����FĄ3����;=E���˗��>�^��
�&t���'|/�<*�!����ڰd�,SoT�e*s�� ��Dgd�4�4�?����e�*Ō���e�h"���lQ?0�z�Vm�>d[a�U[��Zg4��Ou]y $(��9�f|�'�-�����~�հ�s+_t$[\�m"���B�uQ���8��y�"8+�v�
��ት�/����7Ǉ�,ܽ��ĺ�����ɦ�Ǩ�-���gY8��z,*��aT89�^e���/m��	��^T��v
����e�)�7��>b��g��D�U��T�--�'���'�G����YF�hcTs�[�E$������X�*ɖ�/��p�W�J��1��
F3���3��Y�������h�I(%���"S�%��W*� a*ժ��G�@>��+;�P�΍�W�����s��\�{4ў�V�Hy2���sC.�03�c�z5����hT����uO`
���P�p5��f�#d	i�YOc]��J�������*U	�/\�e�Bd��U��C��8���鍁K8g6ڀ\Dg_�bt�hߏG�iҨnX�[�ǟ!����ߠy|ᙏ=��s��]&�	vrB����h2�|��w����M�����������~w�W���=����ΓO]���}\�Ŭ��s�l����*���\a�!��:�G��\�h6�s���}������?��St�d�jZ�����6�]�af�>
���a%���б��=�ј/f�j}���^��+W��g���}c�@�ƌ�'^~�L�N>���}���1��Ͽ�e��E�mQ�2�p{oo�7~�g�0~��3�]�`TԾb�vQ��Q%�E��3�1dNo�%@D�%�2���p^
LmQ�}�AV��~Q겈�b�B�k�Bϋ����3˼����'�r��$����#ϧ%��.��h��\I�v�2�[2	[f�.GAC��_���<7����L��o�hCȧ37��}�J����u[��iAS�[��\,%�^6`�i���"e�R�l�W!2�W#5ĭ�448���.6,���?ߓ���VTP�UW�Bx���޴�8�E�вN}�9�+p��;O���. y�X������p@��eu�u����/~6��p������~�@4����#����7�E[ȣ�v|`�*-s�k��3�AN�W�j�u�b��E�ԥW��P�E�&�}���������[Ve���*��#P��
�_�JkǔF���e�0~�u�����
"��jEj�ڪ����Z��j�5�VK��ڵm��:���Z�Μ�'�m���ѴxO�6�o4O2�6x�{��d���wR.�7��(�t�H8J���{M��p�TVa)��#t���z>�DxCz�u3�8~1>)�ʛ���B����߯Z߰�C��ij�����#L��$�(o��]t"��JF�m8��ؕs�1�T�Gl��^P-=E����|�K2���v�g����{��c����\v��ʢS6�e�T[Y��w.&�jV���|%,;I�dk�5���Z[2ڶ�mj�P�K�.!�I��8� RG����W�T;{�4���o��f%�e���� ��Kq��?����W�DX���K���_1�h�exz�:��+���t��{��򶽦ӛ�	��B�������`P&��B��~`�Y@.�+���uV���TZ`�aA�����	����t$��(�4�JF9/��DV�����N�S�`�2ץ����t˼������?�s?��������[o}��5�������~�{'PG�`#�Ǆ��0)AB��u!���]�K)�2˞{���V���kaM�P�VSM�Z�u��y윫]�햓�aՊ�Ɋ�U���RZ/�^-�߶&_��E����C)5&Ҧ��.��-�-_��n=w7�ji%����Ϛ�Y��-�{.gl�KC*�{�;I���qn-o�?�q�L��e�J����.W��R�j�K����x��>���s�!s�U6Em����1Y>4Kk�.�U�~K�r���qN�n��>G��?l+��q�[��HRjݥ���m� �:ƥ�$i�y����]l���u�n鶡
ժ�ڪ��m��Vm�>\���.���V��l��xj*�������Ny��^Bn?���+]������O���~����󭿿��l/�b�T��D!�]4�՞���������x<%+ys��tP/)p���/�l������^��\Vy^���,/���y^���9�k/O�QYWR�K���t�w�A�#�A�\�HGR: ��y�f�͕��3.x����djI�_��5v��(�SXk���($6!���t.��A�������2=�e������&�fB�A/ʒ����

���ˌ~���L4���Q�������"x!�v
(7tؗ�0�)J��p@2���_h�L�C�!����=�W;5\zg옃�#�(����r��.������������+O_�J�:�y��w�=~��$I������l_�z��w�z�������?��j�߾����?~~����KW>z��x������7ߠ>��K/y^ts~zX.FƋ�F��:��YQ�6��޸��/|q't���������+�l�0�SdL���Y���P7'���CZ�J��Np ��{1j%�L	��'��db�W�yQ�JU��:�]7.��j�����;U�:m�b�T��CS�n}q�§^ycz���sO<q�������?��W/�2�^�y��?�+�=�?���0�*���YU0�C`֣S�}<��������D@�ʵ�8X���� C�j�ӛ�2K/��--�`(��/�*�Q���]�OuK����Mx�	��.tN˯�P=�V�
��oAtGG���Zm��)`6���;MĞ:WfO�2�޾}��KK�|D�B}��䢷�(��|�t8	��v0�-�x-)�<����c֜���x��@���XP#3_~C(������쒇�xl���#h[�㙺>��. հZ�ñ͑�{�	+(�xIyi�ṕ�����ӿ�4\ǞE�.�p˖);���G��
��*��n���&;nN��V�XK:�O�9��р55�5ړ��b.�s�6��t��=a�9�+��N����'�>�rC+���w;�2᫶j�����Z�U�pϹ�S�M[
�<A�͒RKnT�ZB�����eܥ:�~���j'dW�ǟ '�R��Tǂ����x�X |��I$�F~��粬"���jSǛL&�/o��1�F�,���� �O�D�Z�J��Gkt�j�g�8�%mF��J7.a��6n{h�c�q�*�D6���S\��G�~�\,�����s%���]�$���Вe�O�T�j���u��1a�7�q��y�]��|M�onY�P���E�����0P�*'�I�Ҳ�g� y��ㇰFU-R�+5W-�cR���R��ЯЇ���	���}2�e ԄX{R{��f���@x���ٙd}�2������Ç�M�F����`�,��M���	]odg!J�ʩi�	��]p��!� ��ǈ��L4���>W3<z-u䢰�T��;;>B��x��ѣ�aD]��)2�D
KT��LdR[�(�AB� b����W(*[��F�������W��Gt]���:�����;�󩏿���v�����M�����>�,�XF��g�	��CK����v:�&kkR����+U���f��p�eD��Q_��D^��v��yDR�`,-��d���R3v��(�:5snS�6�*�1����I��m��NQfI�S���4���$9��9gfÄ���w w:���v���aZ�:�Z�%%�aÿ�q� n�Ruw��
��YKF��"��7�2ۣ��Sw��O޷o�%�\v�$7L���v��y;���MK��cѼ�^ Ibo����[w� ��
���X�!ɾ$�$�aE���� ��e���g>�.u#�-6I��(/ۦ���Z>���>m��u.E��\�2n+=�U[�o[a�U[�њ'�UN�Ğ@�{n�����Lq�w����0��}�����+�b�'�G��Cׯ������8	}8><{�(
�<�w=mBDn_s�FY�g�y���Dg9(��
0Wu7��^������><=K�T�o1����dQ��ŅU�l�奂Q튪t�j$rT��z!	�UEF�V�z�0�5��Ҭ#R�1W�O�˹oKi#.�ijpyUMS�EW�t����nΡh�DS�l���"Tͩ�`�� 3;�����|�-ư>C��/��L��9�PLZl��E�Dɉ�4]d8�6�|<h$�V&�
�pEP|�����SQ��Y��J$a��o8�?���]�
�I��1r;�T.m�\�ټ�c��ӥ�9���uaF^ao�7�y��!���.Q���C�z�{�p����yt8�����<����J$�~/!��FE����|���!{%���C(�����wh��<?*���η��"Tf����8;�5�"Bz���i$/�^&�:*���4���t]�Gf}�bo�P�PHg�'[�n `!��-�d�cU���C��I��7�G�ۅՑ��n��/�����G)D��4�ꨮ>��W����F�O\�җ�����4�I?�������۷'߿I�_}����CZR�	0�J�:��=F�:�Ŀ@sTTԷD`�زe�h�ŹL��nRy��E�A8�<:-H���SHu;�۵�I��b��K�O�Y ��%�
	K%��a��ɛ�x^γk� ������5���)Y��@@x��Z̒Џt	a�}�M���J0�X��Vү(��P+5��j�i���� �i����X���OY�\�I7��>�F�y�d�$=ҁ��&d��Z����kL���J���4���9ΌiT@��p���"NA?U�Sk)jPWw��w��6ò�	P����ND��P��b�ֆ���uP�"�YP)@��"�w��q�T��rNkBRA]!Z�\���6��H-2�q�(
Ei&�Sͥ��g� rM�4S�	��"����T���%|�Y���L1�(�U[�o[a�U[�і��h.!�������s��_r���N�[W�|�lC�%��9���>6���"�w�JBu
fh�l�(�'�	Q�Iq�����#ya������`�kc��;�1ԁ��Z]PS���S�d�ۛ���P���t�h���.1��!�Js��_��s�$����bEG�倻�KЎ���w�X&=�~-��
�g	��O�8�h*:m �V��mދi��v�4�k|�F�������vm4\�Q�HLN!3����_�|����ԅ���ws��r(��v/#B�A}� A��z�j�4�ix�zѰ�Ѭ̎�̿��
�ԅ��yF��M&��u�^�Y�zD�3Y �,�cY3t���2�� G���b��'����$S��n�C5;�����n�"
�"�2�F���Q���ti˻�h�X���]C%�&��@���<B��w�/}trR�����`�zS�5����zQ���{�k�b�����W�]�*�|.�@�f�DhwlҲV����k���N.%#5�D/�́<F����#<��*�������>��NK�K�j�:�_X�������V�\]�o��!����:ע�A!�@�
��[��]B_w�;��c�q��HO�Wm��G�N���Rxl�Z��V��to.o)���V�O��k�I����8�P&��|��Pc�4�e�Lk�D0�"HA/s�,�QAp� Ki�y�9fV�C� ���w���;$[�)'u]�|p��l�K��|ҭ��HB�������ߊ�Z�U�k+��j��!�m�u��Y��s��r_�;\�tS5v�j��gqdz����!m"ʶ��,O����RR�D��1��454w��www�M6���l}�F6��l<���|����8ӳ�p���C�8���ܹ3r���"I+�^���׿��������BFH¯�i6Mא�>��Y�'�Gd�MOO��~r`q���X/�7���zQ���m酧8���=�2z�dk�=�IƜ[H���`|�ȶ��c��B5��r*F\��%�J�#-!V�Ɍ[۰��H!Sd�x��*���7\�J�l�=�����W�v����%��0�Z�%I���rksV̫���HdY���T�AD� ��
a�"�麍�Y��q� �*���E��##���{��
*�3V�����bŎ��O��V�&��}�K���{� ˎ�L,3�~�V{uUwWW�X	pEє%�93!�&b�����?���1��Ќ����j$���I�XH��@H M���]]۫���5o��9y߭��"d�|�ƫ����{�<�����N��ݽ{��z����[7on̬�B��Q������R������q~����Uӿ����nZH;K�0�j	m�Џ��9�y=;?�<�p˼$E~cof�-S�8h5�v��[�D���4j͹��O�E��u{G|X��ݯ��t�`0�w_z�%hZ���3����^@C|w+� �Vs�?�~�:S����/�;S��k�.Co���N صE>ߌ�� ��z�%9 ��O�z�A{P_�,R����LG珝���\���[��3�0m�K�Έ8���ҝ�i���: �ܒ;��\�ą����_^^.� ��֠c���d�fz$F
�e���� p ���@�e	�X��T������Fy�<f�i��Q�p�=�����Pv��Z�2��ė���u9:@��3�S��B:"*̫GT1LZ�Rw�<3(�	�
қ�^���y�) �N�K����Q���,v���R�>�茌c���pRA�=�Pe)`U�E�p+�+,��,�;��"�H�?JJV.�j��D>�ȡ������Zb,Aa�g�m��^��-+��l#�~��2
��3P	f�����������ʂf��Ic�vL8n���E3N(\B����ck�N��;Wp�Dx0>"+jr�cD����f��Y�Z(>J	�L^Ex~-����dHI5���B��.�R�el�r�Rᑊ��4;���0ɛ**�4�M�n*4-�2-�_�XkZ���2���̋�*�J��T��T�Җ�U�yġ��=O�LD���;��^&�U�� mxU��mC��hJ��8s� �`����޽{��;P��O���	y��lV���j.�d�Z-�Q;u��^Z��;9�)f���Hy4�CI�1Ɉ�3�%��1�W�B��l�]��1�&D��ac���wo��Yo���+C>[&%���}�˸qG���QG�e�4�a�3��F�mjB<����Ǐ�NC��i��wT�e*KȾ�H��&*���)r�:�*�X��I(*�-�h�dw�,��YI�(�yE9�Cfj������Y��+_�@�n��Hu��	h�Çc�\�p�之`s��<^}��W^y:h�#]���p|$�o����f�Zh6���a����f���~{���^�s����LMۤD�0�J�mx��뫄���#�,��O�:p�No�����<������y�&\ ��@� �p���-8 "|5d�b-��ţ�� �>ד��C����_Ce���6LBS��P� ���2 �;{�����_���g��ܹ������z���[��'o��|�����?�777�B�?��OCW?x�G[[[��<q��bn�XŎ�����g�CW�v�b�o��'f��Y!�p�?q�"�<Z�6�q��]�rfa�n����57�I��Z���ew�:��0��Q�n>j-�զ(�����1��w	�\����Ж3��B��v�0f[3xG�����P6z��{� Y��cce���b⟕9�<�8mT��Vf�Y�H���QJ�U�"6`�Q������d���06�����U�i��I���3W.(�ױ�/e��!����g��P�%�v�|�D1�3�<�t#̥a�s	߻�Seoo~2�CS��cK�,��z���&[=	>鳘��U�M�ON���'ƫ����K����i���{�b�i�����ǆ�W/`��e������X�pz��M1N��6r�J�k�:�~�HG�S\�7�y��{��V����o�ە 0T_!-C0m����4�	+�}{�|�����M����k�2�\.��$Kkyq�b:�nG&��0�j8JS����G�fC%��r�9��a0j��I�`b�J՚�29�����<4��<�F�Z�{�dI��&�BaX�3��I��9��0����#�p�0W�g���c4%W.�<n7�� n��Q_�8�l	F���w�ڏ]���lv��`=Zk6}A���j�ȸ1��U\e`�r���z �[YY<ڜQ����Ʋ�He��H�]����"
��in����Hd1*�s#��x���c�KsAp�E%w�wj�	�V/=����|��[?��跗�}�]�c��sَ�u�A�^#��ֶw���o��\�)iOsat��_Ì�5��Շg� a���~�C�f梂�e��f�<SD�3
 �p�$��=0;�Qw��-b5����dufQ!	t�v���l��Ŭ�'�#�9��<rM-�8��:Z�L�`<�@�9����ל��Y�mS8���i+�a%
�Ш�����rм�s�Xn=��/����?{�7;���+o�ໟ��s�g�:؅�y�6�wq}�޵�K�Y���>܀��>y>��M���9O3���]s�^W�^}뭷���pn�� �X����ak�K��W����h��L��V�w?y|F���؋��{�d4�Ԣ�4kԃ&�]#�="��hWl��Cy:�ү��K��y���vg�� ��^��\
u�5��N�b�����ɨ?L�����N�2=|��C(�O�+�^e�W�Ǣ�Uf"--����@e}ÛR�5�n�
:�&Ђ���^�)�|�K�POd0!��S�&LN����L�<��P�f���_����I��K���޻w/lgΜ����y�����կ~5��#�k��9����~��YL;F[r,���+�'HzoމC|X5���U�'�c�7�O
6�ƻW�:��Z����O�%�d�05i�r:��p���� h�����i���2�Z�2-�Ln%NnOƱ��p�X�� �G��`���-fw�ry-i>�����:�`��3#&�1z�޽vXf�g/� ��	g,5��`G `���333`B�����؆Rh���$�����)�T��v`�bd�0�&�y	Q�I�@����J�5s"� Q��I��1��^1�Ɂ�^A����A��s�)���f)mlة����������
��%��6��8RZq�ф�����߼�܇��x��dEY��:
�(Z�UH�%��|���mxh,@&���j��C敃�o���| fF���3�v��� WN�
Y��	Ά��ʯ�
�jp���v�z�N� ��w�ƻְ&��@)�$��y8�#T�#y桧��h~ƙ�Ag�l�f�	=���zLH �
�k�u��@���w���p�>��^"�틟�ٟ��0� �@5r��F�Ã]�=�斖�>D�R��VG��qL�{�ȑs��֚[X����Mk���+b���k��[����Q��O5��#w�F�[;��y���0���۸�رc3ssׯ^����vQ|�s���monn���o�o}����"5N�jBb>��#��}�>4�V��c+�Z"tI_$���9��uϟ?�ĉ���*L���]88����7�Ũ����dZ�����|@;��t�[\O䣫nk~2�(%-~�L�BC�7�YM~���w��}�I��@�,-���s��x���&�"iJ��YyH*�db���Z�����>���T2BGz"?���6	�&��{,�l"��dWOb��_�Yϫ�q���ٞ�?q-�,�P��� y�0(�o��O s���s�[�'�0*���y��rуA�|*-\�����Y��J|�&G���d{�Q�}T;�=�N߳T��o=�ʠ�i��i�Ie���eZ>X��n�1�χ�L�s�Ǳ%��������V� �&�.���O��~*#J�"�����̴w;q��8Ƞ@S Cň+�P�$�1�;1*e��63aoa	�^��6���`��,����z�Aw�Vs�J#��s���H�YlaJW0�u�	Ux� e&r��I�eJ*�9b!I�QK}�0� 'T7w� �,����5X��y�f��R? >=E���"�r�M~-�<�%��&�C���I�lkп6�n@�q[l��C�bq���;2���b��K�����7ި��Z-�aI3�M6L�mw,��|�LЅ�*.x�jk�D��MO�����f0R����'A�<f��|�#ᴇ�ջ�q�i3?##�G:�Y����ko�>}�ҧ>��y2���]w{�y饗޾{�խͧ�?y{˅�h�( �y{� <P���Z��u6BIt���{C��Z5���"B2I膍���x4������g���vW!��I��G�\�>X�Y�p������ݾ��+����=�Z�	H��`��6޹���K��T��C6��~V������AO�|o����^;��o<��T��ܽna���p���0����� _h�G����?�?��G>��|���}��W"�(���Y���^����}����3�{�ݹ�Vj���޿��x䣟��1�x��ƛ��x܅��0g�T�2X�i7�^��Jv��
�ܜ9
�ۗb�h�`�xpq�u c9�Ad�%a��K����'�o��a�������v�?���mm���q+�<ʤ[��.m�SfG�1N$���}	��O��M�r��� �[*KcZ(L~P����Vo��Ͽy�*`�v/���'O�8~��V�� ��ܹ-\� 2-?x#��8�*6/�R��G���""�Uy,C�*�XK�Y^lb+ʬ�?	<��6��K���I���%v5��r�1�7���Ч�߅��T3AM��F��?��~v���x�Eqo?Z\Z�7`�lm<����d���"��5Sa���&F^@g`.ub�V�7V�9ı��1ӲǾ�|z�v��SLW0�-RiR$��l�I�~-�l`/���Sk�@8-��S�)֚�i���w[ ��r^��&�U���#���d�̕*���C�����Kng{���x�+C����E�ENٍ�2�w0�/]����3��6�OG�������Mvƨ��'x��k=��>�e��'�Q�!���~�o��n���-�V
�j�����K�1^�]��{J(Ѧ�"
����QZd��Āj���naTX�jq�����y��nook8�&J4��\:�p-,Q�ME9�HEmee��KE`��E�8L�7Bဩo�rj�4ba��쓟����<�j��p���"�+�[�b� F\�a��na�u$)j�U�mq�C����k_����U���,z���-�@�}@��!qT.�MrV�"�&LkD�[�戽� c;�zKvvQ�Ц�N�?�l6p�=�	����'\g}y=Z}�z�Gk\���:j8�|��zPy��Y��7�!P�ކN�\\^6S.�կ~��O<��sn͇Y�W��c4)�`��ov|�+_�a���@R��<���w��2��D(�r��u̠u��3�<���H��K�d�y���~�&���գp�'>�׾�ݯ��C�^x�9�K%p;/%t癃zqQ:�i�رc�{��Ǿ��/�Bmmm�"͕{ɧ�G�p~��b��X�.����Ce�]��{����4h5����7~�7�s��|�;�@�D�C�Iqgb*�Eqs/�}I�c]6�#v����Dm?|���#G�34'#Nb����1��Q/�%%�\�f���h/���D��:�fU�t<,0.���BW�+k�����$��_M���9��~��ա^�ĕk��+�Ak�U�q8UQ*���:�aR}��_��ن��m�xTQ�hw�����Ʀ��cc`�ɕM;Peב�ܞx��'�|��Q�5&����c[yϮ>�Ȼ�Z�rkZ�eZޫL�ִL�/�-V�jy/��z�&t��7E��vOu�XL��6�WC��w��5����������>=V�9je��q���8��Z��BB^�΍F��=�
� �����U,�{{�^_����̳D������4��S��s�w%�0��!��J-&��)4ǥD���,.��/�gQ�M�U�����LwjXr��*� �� [��
y$�A�	�q��ai����YB�0��X���8��l8�5׆��=�<M�?���u̶�9F*�v��qi�x9@xY�`U��_}��3�&s�#y���.Y?��8:�(+��r8�)[曷oI+�[,�`zQ�ߗ;����bѨ�Ǯ��V:W�~c��8sU ����4��u��"s����C��vM}勵ҔL�0��?��[N�݂��ް`�ӎ���cFj
gb�)���际y��ey9��!b35B����%��v��v���yT��E�����9
���W80��f&�8��}sss3�w�Z��%L* �lOɚB�����h���
��>C��jr�7�Y�8�s�!���:��p���Yg������=��@"���x����lj��w� T0��Z+oot������ �4Wffgg���7��7��`��8.\���?��luq��>�s��ٟ���������ksY3'�Z<��-,*���F�J�8z ��Z���f�r]�,x�B�n&3�>G��FJ�$K��0K6�v�{P[����v�Kc���Lcޮ�z�(F˳�ňc�(G��Cv��n�2� e�V���d�[�rIcD1�E��:�X2괡�����Ξ:=?3;s�췰�������5G+W�x��Z����Z�av1`���Z�`��b���PX�H�sd�ԋ0?5���?Z�x#����eL�#����J�a�걪>�R�V��-�P�ǂ��.Xc�R�;J�It1��B����C����k̮�2:�$N�s���md�	+��b��֜��j�&²5�[��/U5�^UK'_2���M�^F��m;:fB�)��)Rd�e��Jb�<.Kf��u	�֦��i����L�ִL�߱�q�(?[�-�&� ٻ":��f#�e"U$�)VLOҸM�STi����v��
�'�6�# l��2�#D���2�w�e��-0ՑR00�� ��9��g�`0H Z̤�-r��ۊ�z�43[�զ��|3�x6��3�`"IJ��3�",_d7��qN>�<��a��s�|3;31>��2�=� �':� [&\��B�u���R-҃�~n���"�~i���&r�U,[E� �I�Ĉ[\D���F9;)}K�{�f6�H����������gB,v���}��
s��:��U+%�:Iy���!L� ��c#�>.��#G:�W]>L���=��ܩ�7n� �-Lv]��(����H�J���p�J;(�Uh�
M�q��%�܂�~�6�].�b���Ωa�!ł�2�-�X3�W3;���C�P0�j6��^ߡ�0���!�bQ� 5N�֧̰�z�L!�!������&���� �φsU�ݡ+`LG=�E��``��F��Ȥ�>T��q�(h#��x3�:zղ����O��W:juuuyy��5C�2s�$Ӎc����0��I1�e��.i��L���XQ.����%�۔r��k�fA��i�Hy�8����&G�&�<̕�1n�	?��ZdK�CO��[��9�?igǠ���d163��X���K
#c3j��F�s����L��a�)j�M�1&�[�i��E_ynM��s'��
>U�d���ۙS�<�D�����'$1*�[���2�>Ο��
�Є/�`ܧƭGp�5¡�����Eql�d�a�2T�i�,!����<M�8"�Ԝ�e��
kM�p2p`rSﱽ�wo��ջ���=�.�c)H�Xo��O�㚖i���2�Z�2-�T�049��ㅲ7bU�])m��h�L��JB2�0��6V�����a3T\�dY��8�ÕI&��b!9*T�2�˄�02hL��}%Ql���0�U7�G�;`̈́ud��ű��g/.������f��G/*�sM���p��<� �B���T�,��J�F��@�?�$��<7���e� ��9[8ho�ڧ�G.ҍ"��W
I���H��"2��,ǞFΌL2'���*G5�����~ �N;��?��-]so3��wO̶�f�^|���哀a����Hb�b�������;�ԓ"�� ���.#�zwd10������%�2E�¼C�%�����1j̵���/`0�Y����fE{{{��{ΝF����\C�p�@�1az 6��N_{�c�y���\}����/�ϟy�c'���F���/�E[�XɎ`KKG ̷�Ѳ̙�}���k����w�"�\�g�
lW؎�k�$)	9r�-P�"�C׃����i�T,,�0���,V�r��Q��:I�3�
�ӧ�]8���v]��k���m��4�]���=y��3k'���[es�Q>��}��0ʅ�Q�+˩c]�r��Fo߽q}����`�"C|5܇~;�Zt=+�Y2H<�&���F�H6���Z�Cg>$����w��ᾀ��5�wn<��7�7R����+O����@����z����� �~��_B��o��9%�3��SAG9b���[5�Ɏ��l�GC�>s���B�7_,JuM�K"���'���׮�������������_mt:8"�ҫ?|�ʊ�;|�ֵ��Q]8�vh�fvɑ�&z�g56��f�q�(bO�lk6�
0��'i����Y/��=��֣-xfff��Me�j�,;%�B�(P�C$Y���8�������1n�l<?��J����`���m���EҬ�� ͤ"N�8	��8ٮxD�V�	��*���w�&х�䍟�}e������LQF0\����3��0EQ-��3��
���T���<���9�a���I,	C|YF{�n�	�"��V~\iW�q�R����p&�{�W x3�mr7��L�{)��(z�@�J�Y�b!���h��
�0lZ��'�)֚�i� erK�L�fW҈�+v����+���l�>̤I��q�27�rI�T�I��8����W2gH5�'DU�,e���r��K	ˡ�����Pv�4������P�9Gκ��U�M���Í�n��Id����I����Z�F��4�X�V"�>Cp���^8�s�� ��.mS
N[T�i�9U�1;�`2�MG�A���^��a�3����_h΂�m���<�<Ϸ9���{m�w��!8���=]�����a��Z`�����V�iV9�<�31��e٘~�ۨ
h~%�N��3�(-`㉞�r�Fh�Zf,��������_"4�pu�Wh�h�)��Y�R�2��l�3��,��&mF��)���{Z��eܦ��f��n԰����HŤ_3;�$�y77��I��G���0!�e��޽{�W�Vp/ |�ӊ�xQ��I=F9	ׁ�:u�f[YƜE��9����[�p�����uLT���<�� �=�Ё}��fH�1��2Ճ;­�Ļw�����ht���j���Fs��B��/�y���$Td�#�JH�Y3]�.���+߯E�r���6����K����7�	�<y�$\|kk��^�re�ކ�{5�ڵ����?�:��mZ��LUX�>��U��Bw�5�߅��r���rm�fH�A|�	Z��pV��1� i�5�J�Ҭ0��)9j%���1>��`�n�aPq�<�(�U�K�5b�z��Ϫ�ZfP���	Cs�b"'�)k,,]���D<�ةūՉ)"J���q(b<6��b3a��5Z��q:�ڥ�@�����J��&>*K#�3��ȧM�w8s̞��u,��*JUc�*M�����Q�Y��K��\�)*��e2@�~yM˴L�߭L�ִL�#����9[8����8a�s��M���o(n�Q�?YT���z>b��R�e7�p�� ��u�z�d�"0�mD�� [�\��ݑ�h��i�����$�e�yb��w	G���{�#��`�<�k~�"\�k8�Pd`'!hс ��	hXJI{��Ư��/����5���)��'U�#�h����z��RAQ4\"g�5�i�����t�T=��j�����ޒ�����f��m��������J>���VF��)X�n� �t>��o�Sw��y��YPk��a���ض�����h���`f,g����;w\���<&15��,+���Z��SWh6Y��"�V�92�"��g<c�xXN1)�p僡���;w �i� �Yz,7 C��][x�"���Ymg�������~�׿�O��;�<��׎-c<RZ�{�A��e;9�a����)Ss*�m0u�0�"Y =��.�س0�9Ɔ��B��J���J��+!3G�`�)=0��WO�|�`��d�-�є�N Ə�먠�l,.y�*�E��ܦ� �X�ͷ��l_��#�!�>����ǝ��]��.���:.w�V-`��'�z���?~��O~�田��|�ʕ�?��O~���_�����Ç��t% $xJ���z���s��ٹ��!����>t�I	�4q�������	�u�u�n�z��s%ښ�2�7B�Gm��V���L%ܡ�|�u�r/�3nS5�h@)��/��Jv03��m�Qg��d�(���49st������?�������h����_loo˃�?����+Ԁ�d�>WH�

���2�{E!*���>�p.FVF�q�CÃEX����Zk@��\�]��9��y,3�`s���F�>���&�w�7̹����B/��{�#���3���^��ŕ坝���v=���^����e��*��ˡ;\�s,��q)0� ?�Y��Ӆ����b,���
AMFL���0���b�E(e�ZX���@5�+KD�{Lx�k�8j `�T�}���W(���܎uK���<˅,��C]��V��"E�!�A�¥3�;^����TI���21�>����4�}\9:�2N��p`0�1 �����H[��)�=�\�y�_f^�u.,ǵ��L��x����t�l�^�1�_�aS�ִL�{�)֚�i� �z�F�������#�U||U��#퉪jg����3e0��"e��WU�
V�qY�7��K�7{��j���7�@�=���`"���G6�DUC�g�®6�͗�ZjMh�3���J�Q~��C�1��I�,'C��
{��(ª�q�0Ŕ�� F�COT��0$����dvӫ�'R)�W�n�C�.l3j��̀�gc�l�4)��AG��K�|U�� ���)�RM�H����&O�$WA��䎗�/6V�0K`r��$�!3�]f�y?��ΨB+��}���ѣG�?n�m��C(���Ɔ	�
Ð"?Ӂ4��� �i�@A����l�W[���J�!t͹8jT1ӥ&m�����R��+�l�+%�i����⽊|ff&M���D\���:��EZd�3t���P�Ch�����\���4=`��*Tz��<y��'���(�f�\���K�L���@��������l���3��Z=t���ꚣ!����Cen��2�J�����5���ƈ}g�M���{�((�N>Yhvє�&�Bn����x�>� ����C�u&Gm�Yyz2�PC���r���3�0�6����-��D��lT+�4�sz��Tu��?@��h�7�y���p;��fQX��\݃33��	���#G��/^����w��#������={�s�a�`�Еmr����aSJ�)���2Z�S�q
�I@U�'{�z��]\��ѓc�3t�
��X:�P���&�Me����15#K�<�ee�Y���rzT���/`��t�Ie�u�"5KZ�g�RFO;����(R�J�>�l�x���b�8~��U�Y��i��R�XkZ��=����Ox\9ü����c���0�0Ga�20'�Bk�oKM���mL�iX8y�ȕ�$En�!��v����,P=��j�: 0�]�X6�
eg�o�x��+mg��%
�9�bX�(R��0V�6��g�`R���(���G�)�J?��ǵ�?����J�s��-
s�X2����c#��+�*��\��2Z������(��Ҏ�{QqTZˋAÊ�pT��f0{dv��l�V F򠗵��\}_u�>yb�G`�+�/�7=Ƌ�+�^A ��Ŵ�UE�3i�XF��Ȟ�%Q�Q�N�F���T	 �nCN�����IJ��K�~���LTD��̳$�< ����ga{�.�������wG[�Eo�Yk֚u��H5,]���iA�� �8~(�Ϡ��9"�F��%6��+,���e�3JP(s�Z�����
�
��3\>&�0T��[�����1z�[�_P0��4J-`�����
j��ť���PI�9|�@�^�
�)�40�XER�}�F^���c�_:��^�_{��<�̳瞸����?&V�+&p���D��yA6�����ٌ����h3�?-���+-�,�a�ڍ@.�w�}]��1�E�Rv;�Y!$�)�,���0��\湘?�w(�5��f�)�x�LI�P�F�=��a$^*4�(�I����(KXԂ�҇~�����zy)*˷r��5����$�`)0ڞ8���0��%1�v�X!Ɨ&6F�FB ~���b��5�sݟ����� �&,A�(E��Svc?H��8G�YX����3�,�i}ii����/� �O�Xo��^ϝX���'>�a���G)��(B�7���,���SƲ�ZO
Z����a�������6��8f��G�}\F�|��=��E5��V�:L1���L+R~��iʸ*qad��`P�7�
f��r
G'W:�e��x�5��I
�Aq�ı�(���e=�ulG����u������$��� 7~?��-5gR6�a(AȴD~�vL�4�L��t�Ox�M)[�2-�S�XkZ��*dc�9�?1�Lz��o�F�� p����$�t5��J��eRdפ�g%� ��=�u;;;k��h4贸���xiS�U��r!m:�����~��	��,̡z���H�6q��X�=]n޸�4��6�[��`K��S"J���!b|nc�F�hacM,�������.�wy����ֽ1wq��֘���j����ʺ��ZFad�k)�F�[l�����l�á"�;([���۷�s�MHv�Q��l�:]�;�Cφ��@ �2N����8�e�*x_���F�ob�W���?�>�U���|��Jۅ$��/���o}�����i6�S`��j�D�������각
�.2[q��4����R"�A%�=���uA��Ȩ�-c�\ѫ&^��%���*���S�f<�	t�����޽{w�<�������בupP��׫�?���y�/l�ҥK������yrP4��`��}�,�m�R��W�z���o��o��O��Ç ���Na4�|�j�fF�9 �O�N�s�'�z�cǎ���ѣo���믿��?���Qn:x(0�Y����C�iw�9j���{�2]I�U�q�Ʌ��n�DB��3�Vt~N0�D���P��hR�?n�O�{��?��O|�(*%O�v��Żw����w���Gv٢�DIFzR�g�=��Z��!��/��l���~��?�Go����\�o�'O��y���S��^���M	䋶JW��uX;w�s���������˗��=w��p����~���o�0}�������0�����p"&M���4Y�/=Ó�Vu�{z���U��j��:��yՑ��������rc�����6���{�Z�-��V�pH)���ã$�ƥ�ncVq�n�Z����ry��@X8�|wK'oZ�b�q�QL4��̆a�X���8��:������hM˴��b�i��P�����ċFq#��(����↦�h�6GYv�%#S&,n;RIG�=D�h�ÈLj�@R<��x��(דP���vP��d��H��H��7�b�ō�zh��� qdV�R��Lz�Ej�-KTN�H�7�b��lb���(Gc6V�gN��_��[>ud��hMP>)�ӸЎ�)����rY�:��-�3U�Z��w:�{���vl8 m2�o��eC'���$CW���W���OP �z��IΚ~Z�XI�p�ܾs#Ht�fn+YZZ�Q��3�z�+��~+�&���ٌ�֤���3s-�QHL�쵑c�&�ʅy��횼p���jQ�h��4:����q�n�;��-lf�h=�c&HIb3k��a���B0�wz��{;n���l����H)香S�,�"��gyf�'/$����"�"=w��e����(<�qm3�sW��P��H�eu˪	�[s�!}�8�=�R:Z;��0�{A���N��N�`�������t�4_ZX��(�╕e�3sP����_½�6L���E�{'>�]��L �Kٽ�75�B�7�G������=��_���U�YXX�o\�􊣋Q�::uk���+<Ň�8�0+X���e=sY�uГ�]�Ղf���L�a6+29��,�<��'hF86��;*��ܨ��Cg!f#B�J�(O��l��S�:>��.`'o�+�h)H-�um#~@�/sz���Ks�������G?�O �J��}��T��V�~l���]�Ӛ�<���� 8kAx��
���	�،A�K�@�(A����f��ґ��S�uF�+q��汣3��F�lm�\�C������^��}�����?�x�?v a�Y[���݃��|�{��9���\�7�������]<�r����"�	�4͕�@֜�DG����X�j�FO��w9�~0���&u�̟���g�	�qNd=5��v�p�F�Y�2J��K�*�2*���J*�(�g���Ɨf6ΐ�#�GL��"�	(
�L�T�LPs�ky����P�پ����+ɽ&J�0�u�T�׼��崃���̇e�@0�V��L��^jˬ�Yl�^����a�]M˴��e���eZ>@�|ͳ��b�G�8�SJ��q�?m�k��ƻ�`��j5��#`$#z���~��?��q�R���HF���&3fB���o�6��
i�V�� ����̙3���ݻ7k����5�2k�0�O	���C�q�O>��Ҥk��ŵ��:u�I{�O�Umd$}Vd��,(�S�J�� �R#T��K������g��/}}��v�i�R��0)(b��n���A����� �JE�5(�+�f�!G���z�M��`����t;��%�����`� !���|�4NQ7���d���/+� ��ݡ���ʲ�|���%cϸ�ߧ)��՛u��� "�3́6(��)s�(����P�R��<f������0��n}�0���o��`-R7�(Ǘ�c������ge����J2 x�[�ф������e�S����5�\<�Ν;�;|�~���o�箯�c��9�J)R�����g3�0�h'�-�� :yr�w~�w��g߀��5��_~��K���w�4%�1�����ܹ���3H��e=8`��x"nQ h`��*��i-i�ܘ�D����<oƹm��L�v�G��ּz�&��6/�c�x���7$@��8VWWwvv���/A�,��[�pA۞�8�f�k΅>�)�7�����!z������ǜ7�ut��ݻ��!'T�G��\����G?�����+���ĉ'6`��^{��[P�p}�B��J��ψ�� }�[߁~ޠ��/|����n����L����U��͛Ы���_|�A��v���9:�MT@��Y9��'h�ծ��+U+�������גl8&5	�[�e&�:�t��7ٱ��Hձ��Z�3��;)�&��@�RMb�Vl�-u����~��@#>$�E��Ns蜽�\�ަ�`U7�=�R��l"���^7�����0LhC���ґNK���0��r�/�cB�yE?~����=����i��i�b�i��R���)��M��DH�#�K���n-m�w��sV� x֥�^��x�>�8�"G_|�ۦ���V`�Ό����m�3�ZU�v6Z��6<�<BUC��|ᅋGD:�;^�Y�9�'��A~8W�RqA�!]2��� J{G�p�+	��q�B��9
PL�E1K�D�P��uP�//
���l$�h�R��$����ґ�v�8GY7�\+V�����KIE =ZF��谣��.����!�B0�$�ky�ڪYv��Ʈ�X?����삝������n���A�?�%��]H�,���\�u���P�!�/TĢ��=��t�f-p�uH��Eae���C깘Ք{�"V��4����{PMM�xT��UA��~`�"���������������"�$+hB5,k�q���3�U���u�1���ÙVu�� �RE6tp����r8�DcZ*0�m�˼&$W�Y�d��2i�rle�y�VI�"GCb�2g�����~��i� l�.z�,@nI̸�u�\$(:�N/��s�揌�#���.�-���]��xp ���&�����p/���'Z3����wr���(�����wSd*IV���x",6w�Ȟ����(?x�%�)�sݳ��\ZY�^z�����Ml���|���A��kt�� ����� MMD��(q�l�VC�����p���]��x�s+�IA*xd5:+���Q��+�v�e�"ooo�����g��G>~���׾��=K8�u����ׄ-���$)�0w�ܯ[*1�\�]�s�\X}D��~���2��_;~�13#�`��L @o��s3a����s�����\xL�Z��|]kFa��z#E��;�H������!��d�:sac �W鎊U��p�>��;{�l#���mB���DӨ��=U�]�WWF]����O�Z`�ۚԵE����O�)8����]F������kHiե��Sz|k�L�%:�a�q2���ĵ�b0�7E}ցT�,�y�Hk�6�kkz��&�1�,�}�ŀ�"���m7��`Ǌq�ȉcY�G�E���|����)�:���E���"{P�Z�2z�4]�<U�v��L˴��e���eZ>@�%ע()I�ǉL�\O��'���[
��b���$Z4��m"X��Q��%�ʂJ�z��&���Q��rR�K�lZt5R{3����j�> �H;�����1wSrssӝ�����Wo$����-y$x��bBGz�r���;�ta!;�6�M�T�˭e�ñ�c��4alRdr����Nenqi0�ۻ�``��q��$���nD��Rjx�Eh=[6���ݏ������P ���zi���k�ز��or�)ׯ_���[$�n$7'���ʌK
}h1:�X#������Q�O׎/���͏��W�r=��O�F�v�����>�J������0Q<bL��\���A ۠���t H��I%�3��睝�����Gr�'O�F�9��{�Mߺ��p��y8�j��N��:C���N�B� P�C��ݻ��d����\�]��Хy4h6չs�`ntff�8�#������CoDH'��.�ɉ��l��#G���q�QІ�666l�����ݡ-4�8󷶶�V���r9����l��0���n�բw��* ?qָv��U�y��֎~��@�r�{0n�囃����3g���1��+��!�W�;&�.��.Կ���4�خ4�m����Fc����y��6� �b�$V���6=�eǦq���S���8(C������k�+�`\��g�:s�a�N[�k_�Z��)�����G��~���J�*
�� 9TC#����pss�͘��#	�	���k����u�f��sO_�꭮���ñcJdL^��������.\8�lqZv ���g���|o�zu�O"��ҥK�?���VF��_����Pr;{��趭��D��JY������8\]+g���W���;,� �x&�u�T��z��Sm��;�bd]����S@!�cQD#�_99Kf}(�hđ3�ܽYy9�.QR�Erp���/b�7A�+8W��6ԡi�cǎA�AOfI�5Y�L܄�=a�lF��Q֍�Ǩ�盚�eL�M�E���5��ǜ���	�eZ���)֚�i�`żx2�����gc�5g��v
�=O����,��F������$�[�D h������DkG�)T�����D� S�匧 1ʃ��P��]I;Xj�����i��v����Z���p\ÍqkN����s�4r˷U�
u�Q��C�ٱ0�2�օ7:���g�I"��<4�`^�P?�q���ʅ�_r��&�́�Q&�1��Jr?�\��i��2�LF��!�>F�9k�w��v�ù�^g�P�-U�J{*�`��Y�w<�m�gZ� �rɴ��s�i<�MJ�),�~����tF����҅�/� ޺ݽgy����}�,ظ���������/��#-N.�����������Pҵ\�Z9y�s�f:1ˉ�XZB�33�D1�sh�o4
�=�}X�������ך͆�ǂ:�d^�Y�9�Q^�L�]Z�ݙ�6?;�I��ln��f���ż����y5;W�����&����LP�u&��k,$E��(G�ݡ���r);�.�{�)n��ȴ��L��CJ�t4ư�Ⱥ<Nh�HT~g�«acF�|�$�(Y�*9�̞D�a4��	���B���d�+䘅��ģ���O��}�V������,F�� �ܺ�s�6��d)1��0��`� ri2����c�"KJm�g�!��X0|��!h��4�A�I�����[�4z��N����X�����4����a����v�CG��ѣ3��TUDq����Pk���ck�eP'ۏ(/��AK��Q�A  .��$��X�bMמkw�����)�t*��92ØUd�2'�ew�u����z�ݜm&i'ټfV��Ѱ	����f2���-�/��=z������믛���ɩ�����b�f����h���,!�J�ܶ�i�� $�`e��MX&:n�{��W�����+"V
%z�D"V�5|]��Ȉ#��0e��pMe$�#iy�h��3ɴ�;��#n+���~C�y�9�8��Nµ ���[��T�tL`1��K����� �W�N�̤�E��ce�e��iB��n���;�b2����z��̈����؄?՜�`cƖ~���i��i��kM˴��P&-�I�V��'pؘ����o�.}����}\�:���$K�-KL��eM��N��6�L:�@Q��h��+�B��
Fվ����dw�T�sHh���(W�~~�rl<�j��*������щ�n�N���Ab�LɵP�O��"٦6)�[�b��ix�)���luCKP��#!$'Εf���g�����?C�$�0lol�-N�� �s���܆+u]h���*���6�At�ĉs��]���-//��E�ٜ[[;s�̨�*vG���je@�D7�[^|��'�y��|���2�.^��˿��³���%�F#�hms���FY�l���(MVѠu�!�neo��F��G�c��w��5����a�d�I3��s�4�V�7�s�#]a�4R�,C4��F����0i����e+s���_pAh���9aR\0��is���T�I�H����5�F'�pF�q �͚�qŔ<nQI���沚f�����ld�(5��E�X��ݸ~�������
L�#��Q^�(�����z����1���r?�d�W��e����c&[~b�L �0Rno{}���a[�(��0�ڶ�85����3����������o��k����j��Նgi���̮v�K�.�%I�����o[�W��lOvO�>����%L�h���󻝣�֗�7^�^�:��:0o� �cn޼y��-϶��&�&�<�[�?�� �#t������'����������?������˗/?y�8\����PC�7�.e�-��bq��RO�x�ϻ����V�����K>Σ��%�=�A�#�<�8>��c���%��b�֌�%7�sf�QM+��1���B�P�r���$(Z��w��J�����!n|�qzO�X'L~�:���BPS5-����L�ִL�߱���|Ĭ�Z��&���Ql� P���s���`��)Of�(�a't�X��	u,�T*R��1���x�T� �akM���:���X�\i7���Gg��`q&	�Ն�{��i$��^�U��o%�~o~e�
�Y��� 2��8�ij38v�����b����41 �����t����H�E���W���ԫ���r�-\�����K�w�S��5	Cr/������;�ЀEm�9���8���ƪ$������ɠ�u�j:t�g 3�t6�ۮU����p�E? �o�o\��ɓ'?���pss��߀���K�
g���8��E����W������}�;z���Sg���u���>����_���j4j���j����G`�{s�Ն=w�������Xϝ��]Jfw��^}��pTs�s��^g/�o]���:�+MҀ���$�Ԍ�8I=�=;e�)7l�V��m��HI�~v���;���ZU��d�rp�uzۻ[?z�;з��PJ��v�� �{©��;Ȓ^O:�����g�F_0Dt�2q�#�c0'6?�g��Ck�!�BhN:�ʔg��Bɷ�=ύta{�JF��9x,W�Js�z���&)K�pӏ]�׶]/�,�ƛ;��+|m�Q�=�ē�^�����sp��ׯ¿ݷ��Q"��CmE� �q���$� c��*(q{�{���=��?L��>��M�l����D@�r��2�T3�Vk�+3�qY�����Εw��u�y�����@_�L�E��L�ب��&YX����]X���@vw�~�f��Jά�PY<,��F��Y�[�>��P��Ν'����}4ܸq�߼v�x�I�ܗ.`-[��G���~��;��c�E�������/�O|����.߻U�wN������L-�uw7����'N4} ����7��_|�������&'�@��Y�j:��ܴ"C�KrC�#1s�<�K1{/HP��<�����o�1_vRw��qT��5!�Qn��$���9JJ,�?����@c�:F�*�O�^fӥ�+�k4ݵQ$_�'����a��r�qC�6\�x Is�t""5aĘ�H|���e]��+����p|�m<c�z$�V�,�SEY}��Ե5-��e���eZ>@�tU�w������U��FA�|�=�\̍H�E�c�'Ł�����*�w��^BY��Ek��)#0eX��&�8ǉ���k�Jj�0�ZJ���`�e��0V<����G�;�N��#�A0x��p����R�:G���`L�*�M�W�n4�O��)Q��#wP�-e:#�EO�!�K��|���EI��4rKP�Y(\^`�dݿTC~�%~Nfg�F] �Ӿ�f�QYrݹ�� ]D�R
��7pp�݆�ݻ����O}j��y��m���j�.\���:���W���%�m8���P�՟y�ݝ�]� Xg�0ݼy����җ���W��T%������ǎ��>�x�ffff���/y~~�V��.no��34]��34�^�A{�9�����t���4��d+����[��u�ۅF�)Υ�04L*��l�&)��a��@�z44����A+�U��e�̓,��;�s���[��^��K��"aKB[`�fl����x�p�D&q�x��wĄ'�˸c"f�6�ƀ���a5�f�XB*I��$Ֆ������s�[��eV��h1�{�^ݼ�޳���-�#��LA�1��sp��ǂ5��BE}�:~Y`��ð���u�&��:�!�p�+�زQ[J�Z���$'�alw
�&�ucc������hp��w9r䦵�kk�Q9��y��E���K�$[��5#��]Dv�S�q��2s�.�^b,l��v�sx�q+l�j�	��A�za>R,�@�üj`BB?�8^ѕ��$�v� �E*P@�N:�Y=7�4�������#��h	.�'��C���O�����^�r�����>�t&� ^��p=�b�L�P?+���7�v;�r�=��#P��{�o>��w�u��K_�ҷ.>h*j��N�|��7����GV�忌ǰj��g�*Yf(���Q�z^��h�ݺg��5�\[ꮞݴ'|��&��4SԤ'�<�b�Od=�t�Zm�<y�����R�5ˈ�hgsK��l���i��� ��/XsGuf?j�;A�����O������7G�:P�k����m�L��JqG�B�x����}w���_^x��Z�e�|�e�痯�a,�.'�v��R�EHL�x�6�	b-�l$��-T�a!��)� �,/F��1'0z��e���h$����9�E�aH>H��CZ�VR=��x��,�%ʩ���
}�E�̷Z��|��'E��,�;��[/� I,^ZI�7�(3K�E�)tĲ���i9�E�q��q�����"$;l��1��$���+��w����=���[ɼy� ��q4ЗOYz±�]i����w���M7����߀{����e�EJ$C�@Gϳ��KpV���?l{��������*�=��X��-�R<�u�>|��ɇO=����s���m���f4X{ɉn��,����W�i}u�O@<[Z�4oŹ;��	
��N?X]��= �r����񘠔�G27�- SFE��U<:��������Ng��ŭ�O<��i6g ���D�03`�ag粛G�#<Sv|��������X�,̹���x����!�`��Y�\��x0@Y�q���'���=7X[[�k�q����B�(�Z�Se+A�2�#(�K-K�`8���ʕӏ�}Kˡ��0	�<w<��b�w�f �}�ᄚ*@��Y8T���V�Hi0�|/h�؟����_��� ��N­�%`&�dن��4+�4T�#��3P��Z�#�#Xe���2/��:P�6eY`_S���-��z5��p7�D�oT�(�S���,'��v�pmm��B��n{��{�=�tl��U�0n�i�f�Z�o�~7è�8��^���B3�,�0-W����\x�Fq��=Ғ�|۾p�)l��`Q��{��}�0�l��O#b|ű�������ɓ'��)._�Y��/��u���S�_u� ���,.=������Z�'>��Q����!�z�sc,�巘�c���S��W��PGR1ș��ۃ%v#(iv��+bFV]�]!�3��z�0�=�)�?s�"��)(@��=��4�zzf��ua7��4�L�MUuܘ��Hl)��aSW��ĳ�HӼ��z4l��n�r0���$�#��6����L?\��h��*�x�*o2�!C�E�rW��L�}����_���=����&��{��=�wGdM���Lbf��*+1�,�i>ؗfVD`����,�mJV����,�-Q`�j&kX��2���,�ñc�Pa��8����l�)*zf���峠!)s���J�r�΃�x��c���($�"�*'hB�?A��3DD[V����m�i�p z�	�֡q�x{��]���T���;�@���չ�T�n��:(��A����D�AGu\��P�K�V�!���㔶���x��ӧO���"��YxΏ}��~�� 6.^�(tz�w�u�]؜�9���\Rl��H'��l��૫�L�6�<��A؅��۠u�/���o6��o!�!<����ew܁\�k�໏�=���|�D(����{�9x�(Z����� ϟ�c�waFZ;�v���ʽ����3�`��A�A��'A���$�q�^�w�ׇ�J�T���:�NMuV��k=a5�����'��V]�)��ma�k_�Rx�^Ά&�U#�I�G� CX#+C�D�_��F6��Ė���T��c����<�t�GwB������֌�LW:�I����Q)&�[9���;�L�ʸ��j#-�&<�V4�X��^�<y���O}�S��h���*F��C3p�!@�����[�;W�;�G�}&������u^f�h�#�{^@\ ��?��?��Lw��ӗ/�,���`�v[A���e����03W�o_J�c������X/�$Z��{-ِ�f��Ls:Hz',!�g�`��� ���!���	?�nO����ө�h���Z�4���-�S��<�b�#�}g,o�;u��O�8{��`'�9��Zg�C4��P��ٙ+t�˃���4]JS(F���T���8���j��!Kkw�ֵ���z&�{N�ߦQׯ�~�/����9�%���~��Pf�p<�ʩ��6S6-8�
:�{��|��i�c~� �i�
�L���'�zp���4�'�ܖ�1O�u9� �+t%�����^�RiJ�
9bG�:x±}�t\	�a���gQ�N[;H&F�Rp�O�
��@�Xp<a���^�	���J@�x:�n���(��V���ˤ��q�I��Ӟ"����B���Ӥ�Av'nbI�>]�h�[4���,a{�2(�5��2*���7C/�eT��.3�s���kG�'N,4��a8T�*�2ĥ���"�J5"�������b�jd��� �[����k/�y�[���S��+[�'n?v�;� 9�\����\\\9:?�r0l_�HG����N/��Eg������Ҩ;�����r���h��t/���[���ˈ?/m����[#%u$WdSPQq���%f�u;s �o��p��y���+�����ܴ�\ ��h%��JY�-��tO.��t������9��x���Ɩ��V�9���n�6Q6KJ�zpe]@{(�C��d��1�p�v(�DɐT^@ӆJ�T҄�8%ཝ�@�_�m��6�Q�DE��ܦHE;�Vf4N�25HJ��Q^��Ȳ5����&���7��۶�j)�Fg���:�����l��2C��iӂ:��eʉ�^�E���- >嘉�&�
�K,���H#��rBb&|��0ׇ	�*�+�����ۘd/h�,ǣq���e�~?�\ϗ���n_��5ZY�Ǆ��`y������xA��p4j;�o��x��4��މ�Q�����<�GA3v��|����,،��8��<�r� �[{M������k]�v�㝓�N��(V��׿	s�t��|�j	Pj,��P ��:�0�����<0iZsssr�
Mx笕b�fIػ�br���*N1A5b7��zR�x�=����Z"a*%�FY5*c�����n�>c(��0�<❒¥J�C�,��h�qVH�!,�)wf��5��my��c����&}���U5`����I*E/�-��Ø�I60�u i���&�4_u_i9b+GC&��S���j�#���!���_��u��"��/��_Dم��z#Mu�׶� �ZU*V��K[�Nk�k}�v��|>�{�B^��hK>��~�L�U��L�
��� �g*M<
+I�)�0��\�(���$tab����S����1T-�h�Q`�r$��-)|�˝�����p&�ZX��i�ιqA ì2ĭ������68��A
�Y3P��1����
_c<:[�7f�"�.��s���|ۉ�gϚ���	0@\�<QCG=1���"��n�x�����n�P��_��7�����p󫏾��͇��]��A/>|P�����u(o�w����o|Ð�<�%ſ��P�_��6�z޻�F�h���@)̐f�R7���qqqm5��Hj��Roa��������7ߑ�A���iF�	P
���Fz����������o�_�w�XZ��Q�f�]Y�F0d [wV���ECq_͵���+W�@���aYFq����2�4W2�*JÜ%�,��L���Q�Z�~4l���L��B͡9�j%���L�9��!3B����B|����l
úҤ� `�W�߅'�=*�����jW��N�l�ȑ���hgY�� s�e4�`Ы��((юJˇ��Rb77����a5�5� �̕@ӥ��� y5�d)r�����l6���������O��<�hAg��e���C�Y��v�5���~�=���/������́ٍ��T❥�%7D�t��8�V� G\�HFP7��+%ٸ|�����g?��O��:h�&Id��^/�Cx@S�C���A���m7�[��=�W�e��]�^q���E�Ǹ��N�ϳPj�O{6U�ۚT]gۑ��BNh����if��g��8r��0�����>1[�Ә^����I}��i��n!�{`��4!�Mޘ��p�Z�.���z����=���e���Y��ֿ�elXK���O.S�k�����Q�`1_�/P>`�)�ԕ��

~�р�hs����������@�C�[�ʋ�!�R�r�ilH���3���'�c�zU����r�u7p�3��77�_�R���u�A�	��Tg<;3�ַQ��Q��fa�L'z04C[��Aq.T�������\�J|@�Wi��k�A��qA>5��e��z�W-�m� �U���OfY���L*:��>ͦu��s�����l�
S�YA����J�£��o�n�dY�8����)86�i��qF�d��lt!��]���ؕ�oy:.�U�.׾�%��$�%$��TsKf��E�"5b���q�F"KK��?��r.E�9�F!w��D~��Il2VT��g�TZsAv�C~�8Q{�	 �s�
��g9L/�1Y� �?E�|>ϛQ$����8H���V�l(��W./^Xv���|�b�S�Í�*MZ�9d���sv�_�9���b�Ey��#�V~�����z��g��Gs�p�ټ�J�^Q,���	���l�WjO*7�ʍ(=[d�j<�~&��R�D` ���g
����F;KCcyQ��c[��(U�f����r���Xnt@�o�b�Ն���]I�"��x������l�Ӆ�nm�I��A�y�FsA#%�L_Z�l��2%�s:�Kt ����)$�B4}o4���þ�F��P���uc���3% }Y)�>�㒩�R`�b�!2wbYZ��,a3��8����I3�l)���TG9i�ۖ[R|�������*��(���7MS�^K:Me��a��=�%�qX�;��N�4+x2�&��\�n�흍m�5MI�>y��f��hm!?'�'ж<� &Ѷ�ډ� ~z���?�|6&�BױR�x>2�d�a�Æ[kՐ�)1J1���v�Bo{�Xg��9k���~6Ff��9tG�&�a�BL�C ��e�)�H1�_i#����j8��>t����%V�j�Y�ؚ/�ė.̐�?*��(� KG7����q�ݹ��h�	þ��7��[�a�̤E�6�d'䊉Gyj��Nwl��n7�i�i��)e99�dMh��_��X��PS8��(�T5����m��t^�2ae���	J}�
��`�ca7���Q+ �'��d�9�N^H�B�?T��jQ�X ӴI�K�2t����pr~>V� ��2�ޭ�ι���re$19�`b�Pv��q�Bh5�FF���
X�^�+s<��*k �����d��(��~�/ה�9��_L��e�+�"��|eof!Ĕ�U<����ϡ��~�W�*������s�kk2�,N_}����OI|/�����^b�C(f���)�T�]`�*s��s>;9���/���&��_���J�L��Fvqa>zF��y��e��,�Awdd���J+G&4�j��c� �%E<@<������ژ�(,9V��+�l��ϙ�"����lP̌�} t����e3
9q�^�I�r�+a0�ֆ(��c�w gE�jr�Bnʤ�r���_����&�ʇzhs�ޕgϞ�6�}׫@�l��b��^���v���O�ӏ���{<σ>��#kkk?�?x���]__�2A�����!��v��j�򕯄���w!a.N=���	�H�&�[P��C{}�d�'Y������ի�箬��B���4m#�<���V�|���*b�y�k��g.��,�/b�V� u\�-d�Ær��a� PVXv�̰����ja#� I]R^8J:P�8I��H0X��'CW����C!ۈ8�G��p���%�Y������rݵ)w9��>3����	9�0�8^�؁Ym��G��?�� ��o��N��OC���c�I`�[0+2K�籅�9QQql�3�v0���hp뭷r<LFY��-�E��8ځ�p	c���g�# }�.F� ��w�-��666�F�w����|�p����w��?�O�O>�,�"h����s�=����1h�J�����`yy��?�q|��Q�����#NL
m'kv1�<ѣ(���&ن����#W�6Q<S֬B�r������3A���N�ّ��_b���M�L�Z�n���3��/[~,�oYU�g'Ƶ�6�ɺ%��R91�h	�m���'v�Q�{L芛��p�̮�M�q������Y��U�xF�E9�����I�_��1ek���Zdb���:���/,M�nK�T��l5����{��M��A��D��W�L�r���|��&$q.3���g~�kV]Y%�fo�=,+�y/X}�e���?����D�������>�$�6��
�<f���`�E����e�(9��S�r���e�����ǔ�|��+{`�$5;�u���J
֙r�K�&� ��~w��N@S5�����Rf�D�U2E?�PJ��T�!��&��m�.�	�I��43�L8�S�(��KY�Ty�5�G �����(���*.�)1m�b;[I�[c@d�psC�a�!H(R�R��E6��f-��T\I�Y.F�X�-�mǖpAX^���K=�+�r���a�sm���V��z���7@�,;�7�<u�^X\�y�������ҩ��Vo{�tm��7��?s������I�����*l��<��3�YʃV����O-8�����;N�j�����N�LZ����Z��5�F�e�e��3�4�8�I�WV>��3_J�$��'ˆ��~�l:vj�hO̢��A�����(��/]�t�g4C:�����ꄍ\Xe^�����C�����Ma�Vܕ&ו���?�=�Z!��L\���`�����r�w;�n��r
?�繖m����8�%���,Jl���	�H�8c�RDȸ E!�$jӜ�'��hN��Ke׳��ɪU#Ys/��j��kV�vپT`�oX�������q����6|�ؼ���^q�˃�K���2C?Ȋl��-/G0�=xz)��Q���L�*,7�$NN�r�9!�6��]�t�%���j[�ȶ/@wr���
S�D�����-aه��`��)��o���\v�N���xE����\v��o9�8t�X^��؇�!�L�:㻑�G��i��,p���})���ߺ�m���8��x	��8���zn6����zS�*�4��I)	��Չ�EN�&�L|����3N�b�����b�X�`�Z�ot�;Z̎x�tM��8U�|k�6m��%RJ⏥l���O8��S�ѽ�T�t�v7���G��9��o�EH�[��k�#5 =���K�r�G �efa����L��A)�"ǣ`�_��b^��LZ3�f$��$l*ž:����?�)Z��~�/�/�X��/f��
����4�����Zo��+���S��텾��c|g��NP��r�^������-*Wy�wj5��g�Zlt�����L���5�|��n�o����J�PS�/5�^���>1a�6$ q�@Idki������ɐ�[��h4���A����2��/Zց]H��$������` >�q`�<�iڴa<O��MMfPn#ͺl*-�
����1�Q�.�Jt�Z	��Z-̹L�"��'�!%�(.e#���Խ�Z{Ξ=�W�B/_���t2|fkqd_���+�/�>}��B�%�m�������\D~�W���8p`�Cz�2F��3��ҥK;�6N��&敇�%����"���훃��;.V[W�e�w���=sssn�F���L�Ud7�t���ʥ���h M�ǘ�lts�u:s�i(�
fJ_��������C�N_�8u�� E�V)��;yn26A��=)H�E�u�8F�>k)@��[�'N��40����『�c��g�XW�I���xm�џfgTm�g��"��_gQ�=+�g�,Уe��A���P.�����%�d����	_D���0�Ďx��1����B��Ӥ����E�܉��y�3�H	�8�h!I%�DKѴk�xa��Ջ����gVVV^������	*L	c�w���m��v��A��d�۾z������Ǐ���[ؔٻ��n WϞ�ًQ[�l�4s̢��^^^���}�C6�l��w�oYB���[_��c�:4��CY�k�4�ۼ_�+�'�����	A�s��:���<v�)��̆,'�0S�:R�p���=KZ�v\�b�����pz:�*�خ�W�bC���V1�H�l݂�j�[ҢphGeܘ����y���>;|ϙ�%z&��5�'��˲�~�/�+�X�E.�aֵ���"T���6��M�Y�<B�9>���P�E����j�m@�]�=-*fdQP��^ʘ��`ݳ�H�'��L��&u�G�6r�����FJ���R>W$�uJ���݅F�#�a*۵�$[�)&B����=�ZVn0��h	��Y�-M��N�>���T_Z�%5������VB_-a\;�X�_V�OX��R��K�Aݾ�8�Ja�]Kˉ�U���ȼ�H�%���W�F�Ù������Bo��a6��<�3;7%H����*���1�4��ZƑtm��U��8|>��0�.I<<�ԩ�ȢEag�%d�پ�r?hI5.��k�E�%�PI������$`���|�z�D �k�R�Z�QK��P����Ǐ���gJ�iMYZ0�QX�i���-�n�{;�0�*I���PV
}my")t2���sM>�f-��𣋘�,��H���bTF��m��D��6Me���ق^�S�)̔�E�(���"��� �l  �J�� ���1 �ߖ�-��V_z�x��Y��,6�\,��d:��LZ�L(�*�)�ڭ�p�����g���ͤ $��ܶ`�EY��&e��
�yU�������@r.���ʗEE��E���)���ŹC0�*�pf�YSg��
K�K
���D{��h"FvD��47��
 lѲ�҅k�w5�8@~A,��F4�L<~���.sGI���V�_�`V.悷]���v��~��R��h�
[��ci_g����X�����5:��D�>�0Z%Ӄ��/}�)7�D�)d�L�Ұ\��Ғ5�� �B`K��A� �E��*��l5Zaqa��̀��7�Ճ=�[__���y��'.o����^9��$e�	q')E�� ,��X�۽t�ӹ�mUi-lx�u� C�������bi	�CC�D=��:��m,����w}'�h�!&>2�����XKL2IhAjq=�;��e}@�P��jd��vi����6�oC��K���<yHa��F틊�	a�ax��RW�>o��ec ���jS��5�" �#�iz��ʖ�횜���`3,]������`g+����041g�U��"�6C�ZVhL�alXM����l��u�&{��cZc�^���~�/��zek}���������,ρ���k1���mS�v�=�3�95_$|�^/f�~Ѵ�3��X~&��Y�;'Z�=����h��z��-5|������:x��*�\������T�O���גvBy�_���	+���f�#�S
h��82�S�:�V.����0���f�^�9�1:�?!+�9�n�s 6繪��bFҝX�߄�X�%L��ז�$3dok�/ �Icx��V�9�.]����a�~1.���fl�am7���,6�ŗ��;�&|�7Dm���<<���<H�����K ��N�$�&g@:�ܾQn�1?h �bC����;݁D?=�������$�=l=����ٞ'p�>	
� -r0����������$������m��/) >����u~ի^u�m�=𵯂���^���&���U'/��l`��b�da|�����z�=f��؞�k�dDT���0�/��4{%ڣ2]Q��y�m�d��)�7���<�-�u��"g݅��'a���b���M�$��Y���@�{E��=�p�ǚ	c��tL�EZ��ZQ�j���[n�%+r�7nb��7�����S�@{��>�/t,F���-//?9������իW��)dt[�4��?^�~�:c�"<��{��t:A�<�Ņg�}����ݲ����<��;^��W�|ӽ�~�g?���������30�ݭ+��"=� �p$O��Ok61�l�����ťv����n����~����
�G}�tZHC9��0�Ν;O8�|��ɓ�{�[[[�$Ʋ"�1�,|�Nj��5�#s9Z�"v�ԛ�1����nV�|֓��wg��:���7zj�63���Sv�	��U���G�_��5++�ǫ�^0�{e>-3���F�<�5Y�]z �G����ƸVdh����0��u�rT��,)k���<�'k�/��Z���w���[̬��
�A��O,:8�f�A�Gg�p�hZ��G"71=�5���h� A��-EhJ-�������5̙h�Vӻ�@3�;�?���bY$v�ʝ��"B�F�E �K�vM��1�����N�=�Ue)b�ٌ��vM�=<:F�~�ߵ�%�V//RZjb��&���lY�2�L�+��43E_FT��tf�, ���XLcdl�߲���xVJx���4i�A�#g:�����`�]�m��u��m�ZTiZ,�`X�i̠�/L�^=¥X���i���7��X�W�L���x'����К_Y�K��yL�Z�5�8�2�z��GL�$�L\{��VY8F�4V4,WH���Tq)T3�	x��0=)'��6*��|f{Me����������ʳ����UVi#Q��X%Ɖm����r4t=��ކ̆�I��(˵���M�;��Ҝy���mxT��vז�L��K����0JK^���d"u�\�
mo������\�r%ϡ��֑eF�廘A�hXq�U��Em��v��9�z ��e��)��;E�B��_�������KQ��h�p��qM'�I���/��H�ʳ�&�2�
/��̇�M�������J�B�L�iDl�A*K�w��i��R+(�g���Az�0�JF ��R�$�����7�Z��r`��B��������]J?�y�6)!�rG��@�eZ�^��C�?l[��SLJe�iB{i��(%oO�Lլ���.�e�W�e��!�r=�9�?�:��Ƒ��q#���E����a����[G�[v�h4 
ò�{�D��d8�ʷ�TSyʨ��մ����̆�ny��8��_Xo?Y\l&	`-�����6�*�y��p\lw7���j�#���p{��m���x8�;�X��sK��!]5���;��][=��Y���%_��6��Ћz%�w����^X�.�� h��K���Μ9�ʠ�itng�ܼZZ&<v 5�0��qʟ �[�4�9&��+/��*��[D;��tP����J/EѲ�v܊���UI	���*��d��e�ND'�,G��d{���	��d݀mPb��+��*�o��C+|BK���2�HhM�Ȇ�+læ�����"�FӤ��7	���A���"��8��6�p���Z�}'�I��&`� � t�����,J�A�+,�kibE���p���_^�����?*��S�`�;Kr��Y˕�~k��Ym�w����}72��lI�l@����}�Qfa	�ZT���.M���L�e]�4E���JCi���Y�5{e-��	o����e��b
K&כּbVKzݮ�z֢R��M�x���/&*ҩw�Gb�g���T��Η���n}?�RQⰠhu��,a|@�ח���`a.�Fsyy9��(���	�fE)*��$�]P�����owĞ�V����(�d���o�Wû�,��Q�Y�fi*��@��z����@�8qO��`�ϒ��1�����<��lr�^��� �@淢İB�/�u�"�!G|1���"Y����Ŗ=�]3�As�:f*��PF&�>��C6E�~�v���J2h�A���*v�gea�G��F3�"/�1'/%�j ��>��om���CK��\ԟK���$Q�1�51Rr0Rg�RQ�N�-��ƒi�
��
J��Xnuu{ ���!&Ȍ�eĚ�픧�E�ճ|��_k�27�m�_� ��?q�8.FUA��
m��.l����v�{��4��b��K9��!00�]
Ѵ�Ɠ"6��8�ˌo����ڲ�EƴҸ���=w�\�0vq��j�`����W���<{��Kp1J$�i��W7��?��X��=|��7�����Ύg����фK+�����O���C`&��:u�ѥ�ứF+٣�>
�|�cge���NY���h�f�SO�5ɫ�у�ֽ簘��0iv92�����ß��fb�~+��7��B�ؠ�Ι=Ʈ�֙	�P}����6ML�v�+_j���֙�W4���<�ے�b�G�w"�|\����~�/ߍ���^�b(�$����-D)�-���CQ���e��b�k9e�d�s�����đ%�T������I҅ʹq�c�e�X�r��&�b�~�_�mJ%;�+<�;<\(��;��0��(�����z�|�(ׇ,@J�<LjpC�ș�@�$1�����>���s��4��(��ˡ� �R�)<-0
)��P�,ҡ;�+hܱQ�d�Լ�L*�G�0AM��y&!" �a'Xćk;�Ʋ���2.L ;!��=n�`V��Yjϲ���i��LV���Lc~*:��"c��" ���^1t�A+����R�c90`���ؔ�EnH�H=�P!��)Hj�5��ȉ�����-{R��ҧS�\{A�4O�E9f\�D[̤ȡ��cߢ	�ly�o%�U��Nw�Ew�K��C�C�e�fw�7�z�����=r&u�9��z+�]h4���K6{�x|��^���X��"�)h�9��c]:��1.?��Px�� ��]�G���ᫍ��t���~��3���H���o!�F��㎝�n�}�A�i��g6zW}%3��5�*-�qp�����zν8΋�@(�#AXi[օ!�\m��K-�^,LsyiQ�E.X�]a��i������YYY����u��`�cec!��tہe��E�Kk~�(����,oy�hxemm��j[2l�}۳�n�?���Dc��|  ��IDAT�a�� 𧽰�����+˘�8t�,à�i���}��G�V�/,p�̙5LG�|��ܻ`yk��p�(�wa=��6_�@��p�7��g�FgEY�Ш�-$,T��D����B�A[�tF�E4}�U��m�9K�8B5�k���kQ�:�8����9�����0Q����LH�P9��(M`㠜Y�a��K� f���˶�ϊ�WQTb?.s����vP��J-�𞉮���t��%f���׷&WZ~�Д}���UE�0��|�c�,������ �.���Wa���:Iz�2MC�ͣ��v9.L����"o��͝������W:��݄�^!�|���12�:�O(��g77��K��̉�|ٳ��3�9�hx~�ܳ���}�S�h���EI��+�"4�"��y%���#/?�Xj'���\����?��?�,�>���]~�ٻ_��n�1��O�X�뮻^v��A-�*ɋ���q$����d�=Y%	�:g,���=�kB��b����c��U���X���M~~��`ܟ�p:,҆����Jz�26&�6%@��v�i��"�����0�K���x:ȉ����*4JQ`� u�rm�g�Y�4�c*�N'�?�1�12�a�g%6O��IF�������V��s�u�",�VF�+q��� VB=	g�*N��}��~�//��c���Q�Dc������I����u(M3ʒAb7ai[�]� 
䘗���PIsD�[�LRT��I�R�����*�Z��!�DQ��>|V�w|�p`�:UK��v|�b�����B����@x�-��� ^��8��A�F8�Ɂ"X7r� ��5*Xt�)�N��� � �E�+�8Q��B�	΄	�R�
>��:���z\���%�6�7�9 t��T0&�P�G����6�1�Ol@x�6���u�B�9T�l�ڣg�X�F�?b�>5q����_Q3�Lf��Շ��gf3����G(^b�t�ɪ�nquY2�1��i
֡B��xT��h����0T��(�ۣ���MQ�$!�Jr������5ɈQ�2� �QG�&��v�N� Y	������p�>:��z �<��cs����(�x#W��'����-��1�����S� ��V���aZw6!@�L��pr&9�aC4��C�b%�,&��X^��s��`�y���SbRh���c-��ASn0����0͂@Y�Oa? �'�;1y.��xD��1B�f�4/�XD�A�Y�� x�!���d؃��` ��?�ޑ��2��F�A}��1�'��A��Ա1��x��z�7�&3�,;�7��"����W\��z6g^�bF8�xʁ�SW����d{>e� R�����݆�O6[`���2St�F���C\6X!kKn ��Dl�ہA����&o�U�=��6F�6�7��;�� ;�8Ί�Z��q��:��(�'�|z1C�a�9|n.�w��<l[�6Ix����AB�����z'X�������dh�vm�Es�6�U)/_�|�w��� Ii�_��b�-����k�\kD�}�j��@;3����w����I `5�r����;�d�NMj�u��0g,�T�!�#���[~�{���y��d�2�gAI1��F�ѧxO��[��
i!E:c��~׉��֭��_��ek��D8�`#�m�DFv/@��4��|�
2Z�lH�E��.�h֐y��pQ�y��j3���#��%d�26��5kd�}m����{+\���~��Ίh��j&ނY�� �*�lk��"��$ �b�ځ����}��2���)��J�xNC��4�Z�cI4}��#{1q�HY�f�\T����N8��2���*�A��4����DnX�GaN�1Q��<�7�u��*%ɚ��c;cR�,p~�3�_;+��'K���
��q��L��-Np�jI�Z��l��}�-c�U]�fa�H�=�'�8�$�<��D�X���%��b 4�K���{reZgv�z�L_5Ud����B�D��T�0��q�v�*��{n���4U���5��ps�aBx��䷆!O��E0'q�z�p$6��|?Ї�^�sS�ԌzY0���u{W1GA_�R�SiNN`!՟,T�4M��$;Sde2R�݀����������K���n���Ð�lgF�,}7%�Y
��ʹzK��4�'=�����\�
��)�%��l��-�X��2doDm��ruۨ �K�M���l�N^��˛���D/�oa�8�`}�N�Д��a�'�t�7�֎���EoL��p4܁���Q�����o��C��:�����~�7~�u��+ܠ���ɓ-�`�� ��~�M'�^���?��D�H{W���Tߔ�B��ʢ5b���iĊg��q�,6�;��J�F �f��|I�
�9�`���$�<�`�6ѻ��:C6=˖eS��I��iB#`{1���<�0P�.q�*��f%��Sb#�$<�.c�f:�J����d��"*�b���J�Tq�j{����:EꙠ\� �+��ϲ
��G�{lR�홥��� En>|�t�) Z;;]���W�]�W������~�u�C�I�� �~q9**�P�	�	\�v�.a\�b_ǖ�=�؈�S� �a��J�ɬ�d�pg�����{@JW6/"6�b��3��"xn��~�}Q<ē&�]�\�8Yb)m��x��ٸ�{�>�=�zz��o=1.�w��5��[�s`���Z=|�ĉe�j�H.\��?��[o�����o=y�S;"o��~�x�GEjibtD�
�#2�i��RGzͩ��5LU����W"�ބd�Ph��	����=��_M/'� {W����h�Q����i�K�)Ez�2�gYd��|Uj��R�騺�sNab5�(A�5�l�"��tʯU$�h�z�+�L�"�� nr�ݰ,~�y��3��g 1%rC����D���vrS;32�&�B�%�U���~�//R��Z/rq]8M3�PAd���k_��=��W����|!
�����ȗgd��������yn��D�dH7��o����0E���qC��nNO���СC��{�����Ϛ�)li�&�\�G��ԩS?�#?r���Օ�?��?��_���-p�)���?��?�����j0 ��+�a���������������_}�o}�b�:R��_������Bo�K�]A�o������o%IL	���`�J�M0�����=�����[��6�<�V�	��=��_�����c�<@e�#�	+����<O�~����~�F�����0@��oy�[����#W\ۂ;���?���/�ڡPc�󐙄s�X�,f\Y�[G^���wu��y½�I-j���hI�W�4Y�-ˈ~��r��Z�)&�Ұ�D@q�c`*LW�zZm)j��mI�6�fCkmA%oI�B �wm�I��k�1E�"��aV�>Ae�$��1`�D��^��pN�̿����f��� ��dMB�j�d ��5�� ����rss3̎F���-S�s�Z9�&4=-��4hO��ƾ=�@��KP�IIR�	��U�,+������J��p8����a�e�X�t8p`}�R��@E��׻�Ė�1�S���A�� X]]E�=m�z���&|k��t���"}�G([z�aK��P�f�+�T�lR&�.�ٸ�`��{�K�8��"Y��#�������������F�԰����F���B�"ں)Y�4җy���C����~E����K(�F�q�Y��]{�\@��]���ó�iBS1�}���ϭ���7���z�ГTo��Ŋ-��O�� �,,,,--^�\g�: .x}�߇I�����Zm�j���u�:�$��L�e�3��(v��!l�4�7��E���V��{޲� Y>X�FS[�<''��6�z�Ǳ8z���K�NZ	�7!��8FDW0'��kkkG��:;y�رc�7��KN[YY<P��Ehnd��Q���v�{���jSҵ=��0���w�,K�9��;�FVb�&)*�6M�U��o���<6�W*F�M�mEB�7���:8bb$pg���~\[��X����ߢ�w��v�|�;�n�&���?S�Ć���_�{ek��vK�ͳD�²��D�2$�=����N�l��C�����,7��s4d���V�O��������;Ｓ4��Z.�q��������_@�_t�b����$�8����w������t�&��i�%/;��U�w�wo��|�#�^j+G�z���}�ڂHٴ0���iz�oTy��V�XXkt�['��2�
Y����9�У��A�Jr<�9Ɨ�Q�go`���g��|��E�1��8�A���*�K���N)
�$/��% F
����aÅƂ����>� i���g_������]��o?������o��o�LɑZ�"��������ݦ(e�Ui0���PX��$ծ`g�.���"|J�1{�Q���Xy��5a�WD�N������H��,^��WS���g�]��lZ��J%�^���.?��0E����/�|V�[�����i�x��y(� 0����Z��X *�=ԇ�c���h�Ei�	[ƅ8��#��
���D�g�#�f�­�m�2ygq�Y�*�vi�-LG���l�H�"I`ƶZ�bgG��Zkc����,��E���Cj���`!yr/�J�\��/3�[��?��P��%�%�B��w�>��r�wȐ�1^]�.ooô}o�=��C����hs[��Y�V��~Y��б�!-��)����h�}���Ϟ{���&l���h�}�����x�]��KWw�:���[�_=��q��,���l��oK����Ս�����x<B�.�N�5�X����i�#�~�W��N�����A�F�8\t^�_>�|��,+�����F;�"+�q�C_���U��;#���t��e��m�J
�V�y���#lQ%�q��_�Kj8A�-m����/�:
��W
��4���-��箦( 5�Z�j����&�+f�-��
}㸔��]���T�$1�E<��L��X�
}�~������@)7��u��3e��80ߴ�g�� ��^��Wz����`��Z,��Cc%3І�9���(I���Pb�P��@����uU�Eqe�zݟ~����D��Ky�ܹ͍�����O=�ؙ�A#<�����[N�6��i>|���1M�j�YΦiw{ki�}n{=~���5Z�=?r�p�������H�߿�WO;~��cЊ���?9s�̉�U��'���k��5gķcznxp-~�Hb)Y�eo���O��jN���TԬ�ht#�E��
U�*/d�x	Y
Q�h2�z%r�XEZdv!l�^TV&f��k�ϕS��E�&�x\H�Z(��B�\����x��%�!�T���&�����L�DW�k�si�wwe�Bp:g�z��'��N*���_��wT��֋\��X��(�2�a���84�R�s�=8i���A�s�������w�k�!����O���>�����=_���fЋkW2�����O���U5������}~������_��_e�C�_����w�[��;�=s��k^� $_��W_�����>��O��M�L�i�/B�^x��W��]�|~�G�K_���E���>��w��(3�UK�@���?���������{=��.���-u�����<�f�f)������]�"d��p�D���)6&Eo%��������ͻPwk9��3?�3��'����AU៮���k��ko|����7����e"T�3fް��`�_̬�������Z�*g��kAS�����Xr� j9��:���v1�;]W1L���s���tl��1m��o��ϱhw*J�y�����'�i��jN����<0ha�B�
���X��%�*��0?O#�8 �m������P��4��Ć4Oh�d�T)Q���S�]�4�IX}x��Q��`#���Ŗf��{�7$e�����f1�{�K�^��jmmmւ��8Y]]=��3P�x8$��7ƺ2��$���
��Q�w������7Z�K�@�.̌�6��prZP!M�aW�"L��l�f��3�"&풼1���°B{¹�[z:�޾��[�������СC2n9rDb���F��,�F�zF.�'e�%����h�:@QN�#]c@�,�ɚc����eq���ŵGz�3���n��_��d���A����:�;
s.&�����Rhq=~���`-�5�Q�.e�777��\s�.Yh��.5�(�R��c���E��:��r��Y��>��ʸ����i�߿|i��U�`�"�s��e�������ɨE��[�[\\�晇������.]�;�򕯼�������<�@��Kz�!��1׀Ʈ��scѼF�Kz��r�<��q2ʻ�4�N�1�ș�Z�B�:���OH���Ȫ��+r&�H=�{�f9@QO�T�dV�QS.2O�h���J�>�g#Y����QxeQ�\V���$/�Vk��n�� %��[J񫜃KQ�jY������+�$fx�&���� ���_^Ĳ��^��MI$/�p*�1K������@�]�� ���B;�+ͨԈ�>�ѿ~�;��7��'?�ɟ��]p48"��׾�_��O����W��ԩS|0��;8����g>������灠r�C|�6��6t�ؑ������~������W݅G�2���?�������8z~ӵ]��G��|y��o}���?����z�M�BV;����� �QR$�����^��ן~ꉷ{�!wL��z��('Or��h��ek}�Qgp=/��4��l�I��h��P �f#hB������s���_�{�;?��|ꓟy���:�h��s�=ozӛ~�w~&;����PoZ���3�`F*���o@�N��r���{W �,�!K�yա���M݃
}h�I��uU��sU����&�b�p�
T���]��J�I�`&Y�lDM�8K
Y
׆��gi�����Es*�p��`����f9ǀΗ$�`|	j���p�5�K=�eL���9�/e��7�G�Lg����������� <��3���o=� �Sy��O˹�;-/�9s����R������Y�2x|4����m�������iR��1 ���t���)H��ضp[�d��%�k�r��bd�.��`t�'s���WmO �w��+�NK����܁y�Y���t�<)�=������;��n��뎯�áq�ޒo�.?��v1O�;N�72��\^Z&g[*� 6��ŕ���n�#�Y�/@9��ׯ��R�]4$�斂~D~�����1��[�#�]S@;��~.���Ww�SB�Ǟ~�O---!q��D����wkkClN9����N,��U$��  _�P���n�Ѣ�`Ji�!��@N?#3��K�ܲ�jS vGX�A�0$.:+`��@;�XH�X��)H��KO��;��9��4:�̋*F�y+�1��2y ������%����qL���9y�2�Y�#���>��^�ïyͣ��1��==�����G�B+������4i�ª[�M3$&N�4�LӅʦ�3�"�TD�h��f/*���3��g7��	a{�0<�6����F�����;�L�}�U�s��`<�[�V�96֟=>7j�o_ʆ_���Ʃ������� �Zi�v��Ï<4�76`^-�X^^�.n̅�n�ZR1n�-Ru�i�V]f��3s���,�y/����X	eM0��$+j�<��3�yX(�c�L
�&.e��_M�Du��s�S�v�+��	P'EԺ�D/L�%�^�"%EɄG��%���o��-Ez��:v��~�����nK�󰒥p2�%V��~Og�Χ��!`������S�
�!��%�熁��e��R��֋\ h�<�(�OH�K֎g��ab��yDE�^)e��O�{/l���{���|�������O��h� ����>uO?��'>����=�4}�>Z�+p��}����+G�gνJ#Hi�@x�붓��_��_�={��w����_�G�F+�
�|��Is�w�~�~�����7q4��y{2/��F��h�=B��Z7N4��!Ƌ������	�tY��A0ĚE�^��X�K��(�(�4�7K�D� ���஻���>𶷽-�M��=�Z�{������C�L����1&����?J_�`'�RV�s��X�Y�V](�Am#�����@�:��+�!⹧���qʟB>*�cNf�`k��v��D��pe&���_�����zA�b��YM+����H�7PҮ�Qr݈3�fiʥ�Q1�MO���`��w�[o���~��SO=%r��s��'n�����͒��.e�)����w����7���*�D眫�{�}�{��r��=In �Q�)!�IBH�_�g�
:�b�+�����V��=�|
�h���!	Q H @Br�Mw�ӟݭ~���f���9��0
�d���Zs����7�����E�^�-��Sk״2BK�cЧ�b'��!�
�2�H�=--�2���[(�ܢ�U���n ��.Ez*(�X��sȕ��Bk�E���l�i���-��	\N���"�ý���Ԃ���ѣGo��
C���ĉ��S�����D�N�m۶MsZ����?�5�/��r$�_��wH{.��cRE�V�3�:��A��fe�H}{�֭{�_��?�&�&�`%Ct��S��a�s��@m�ױX|��g=�䇾FI��T%L�\��|Z�"G!�\�g]�N\�:�ј�b�x��r���mr�,�*���E�),����\X�jlYc�J̕:t��O<1\���` ���Y����!Q�g��$Y���H�����3H����Y�'�!�ݻwcvVw��rH��M���#�HD��k�<�"Z��m�N��5�D���+��۵�_��l������ǁN��S��h��c���
˶�O���{aS�Vm�k��9h��lS�����n%s��j��Пو�D3|c�8@@� }�A@��^�`n
�Pb�-J���J�J�YX�Y��@��?�Ҩ�"C~�k��^?m�ӧOO3)�T�5�b��� ��m.���>��D�Gc�A�A���v���l�֋�0P���1�V�X�8�6����e��] h�m���63X�Ʋ���R� ���nm������O��-���k����w_�	<_�~�D�N����9 �"f����"8?��O��÷N��H8*t��df%�@�)�ɋ<H�������O���L����������}��锸����D�g�@��� �D1!n�G/=x��R��T�);��v��h��z�?�����}CQ��-�m�B��N Z@<��8R0|BN鄄>\�P�@	���>F!��1�+�n�s���b&��Y��T���P�5@��Fu��}�x�k�����'�X�S�����V0}�'?{�u=����(C�~��JV@�Daʠ�A���bi�� B=���H06(;�� U#F�lCea���r�)&l���� M{A)���Z���<�M A���=k����w�����BgJY�����X�9I,�iɈ^SW�yY�@�@���b�YE�2JA(�D�J�CՊ��J5��3�u�8*�
��:�E�[�n��ġm�%ybW�B�0��R���?�ġc�C����(m/��S3S���g/�t�-�yMgF�:�0m�2i8rl+�$���9l�L���/�jD;2:x)&���9���?�I�íll�)\���
[�T�@"���P�i�+��U���"�e���<�h��ȳ<�cd��D9��׎���&@�Pݒ +:�F�pM�:[�N٭G�>����䃊��;���o�}�T?|"M�r�a�\���'�?�o���@G�b�V�(w���8zSS�IKĸ�@ޠ	#����L��EuO?��+��5^�c7<��>�c�޿}���{�ǃD���Vx��K�Q���]�#'&&���}����*�W��b�nS�"p-���6�C�
C�pF����� ��ڥ(J3z��Ӊ�y�Hd5I��%�$M� �61=J� �����E|6�ޣ\��_Yϐj͕*;q�2M��eM!����Ca[:Ç�#W	�b�T ��lS?R��D�iR�Iu�G1L��Jfa�r��� v���c������Q�Itf�� �h;��-8F�A�6x��1(�҃�ƒ����!��"��W��(��D�MA��^z>��tL4@�,F���0���RܘY	{�%������^� �T��L�8l�Zf��`p39���r���m9����Qy�v�쏻��=��hU�&>���m�Fӗ�b
�6ŗ�!�܄ӢBY�*�-ȦcY��x,x���@�d�U 4��O0~��eD�[�EH�L������IY9����4Wx�OtO-,t��-[��cof�C����:�%�//{�A?Z__O3a�ذ��}����Dh�z=8!���,�}��@X_t�E _�4��3�w��{� ��~�$GL���/�v��I\c�9z}m Wsr���CB<:<S	\��c�E���������ZM0��H�ld���6p|�Z�JMo� �M=���y��������O�*k+ȕQ{�*�^[VEnkH&�B3�� ��J��D�#շ����h���#�?~��;�;'�pU�N-�������'R ��r�TQ��W���/�A#��h ���
���x��Ǐɣ���Z�Ef#Š�x4�[HN:�=�����\��2O2�Z���ɟ\s�5�����5C�}�IԌ	!�_��&�e4z�w���;���9)@��H����~��k�q�8V����0r8D��Dg�)�b���/����ޟ���OӼ��e��3�h������Ꮂ9��X��)��6WIvق����������tR29����q{�((�Aϓ�e.�QW5{��	����
bD�reL��Ζ�>60�f.VFK
fj�+�1$rwKWj݆����u�ĉ��4���N���g�.��ݻwW+݁/t�]�|��� �e�̮�M�m�5�(����zfKg�)#x���h�%��b�F�����N��yT9Q�W�C��l-�KɐK���kee�.��:Y������T���VY.�vmFoqa��%�ބ+�xbbb�.R�6���V�M������>}����\��g�}�.�4N�U3��!Bt*Z�0)\M���
�Z��e� ax��(��囆�o�F���A�#kNR��0��v	�13$����y�T�dU7ޤF��1g�>sF~�l<����1��5p:�ـ���N�X�4b8\ݹ�PaY*M�oa[�YѠ��ݡzz�K���X:q�$ʐ�^rxz�M�gHFB����4�S�TUُ��Ec|6�2��]4��DCZ�r��ͧ�U]�MRь�Y�_�U�hnF3n��+���#r�_�� ��N�x�V���J���a�SX�Lf/&'1>s�~a�h���neeu��s�{��-�Hۘ?��W����O<+|Ϟ}�� _��î̊q�I�Ʀ�]�~�a/h!���� WzO<�D�[K�Զ
����$<х.��⋟��s�۹�9�4b�ď@k`���������Yl��[b?)�O�w���Z/zc�9�>����G�z�,��:g�k��Q(&cEu�2���,���1r�dw4m���>:��d��駎��o<x0��p��<����4D]�� zɥ�������wFh���"y�k�߶c��z�1�z�i}�#y��+m�79s�M7}�/�{��bt{enw&�b��"%�X�������������F��6�Vf�grL�F�/��ȕ�)��B�"��D���G��T1�0���b���e�a\�*�`6��$*V/�8��4ׅ��RQa�-F�u�[��3kK���g�:����,Q:��@G�<a1#jx��J�A�U���yAr�5�q)e��0TU�5i0�-�2mKYS-�l%(VD�1(�6����Ya�M5�<i�BO��0�Q;�H�yc;�#2&6�U�ږ�xq�`����0)6ư��yhb#���4`W ��DRxl���9����{kC�N���ss3��[��VV{���N��~��=��n~���\%%�y�;r?@?�j^�����h*m%����qq��	׽��х5�?s{q.������=��	�E$ڠ[f1,:4���%�V�?�-Q)8Cӣ��D_g\t�JGQM�!�UfQfkfj���y��:�S3��u��m���d{�#���v�:�넰��̖�#l�6�ւ�:��T�ۦ�� w|'��j�=�3�Q2�����|���Q)r������۞x��"�ɓ_~�駎///��0+���ڰ�@��:��q��mپmN��3ۗC�8 =:!c`km.�"4AE��v9�N���!��e[�6�(���^����&a�먤��\A��*R�wu=]��+Պ?��f�)��v�.��Z��6kQ�i��ez&��&x�3�9�H��;��8�82#Zӓ���(��M�,˫k���;�8��txS2$�HE	f��by�`�1�Mq�S۩B��K{?�af�������z.>�ҊW�1	s�B@{�\�"��Q�,��J��`�Y����a)@�[�9B���N��v�E�!�� �T�\Μ����j�㮍��X�����>�����1w|Ә���Ry����,WR�h�Ȓ<�i��N����-s۶E>
�'�z
�H?�aݶ����G?�W�0�2��i�l�� c;�Y����z��?jO�v�dF/..qD��SQ��B�G��ܶ�?�zX��zma�_������ }����`{���� H3�7k�Ф~��KW�L�F|�AF)#=��2��D�o�j�k���LԦ7�Ǻ����c��Ѳ�lT��i8�7��9IV�vP �AU{>�h���R1�2M���&p����&�۶m�v;�(W##+������;o���~��o��������u�]Մ}.~�7����I8B\w2p8�����ӌ�)t�
I�(UW��������/�<��_�������گ�ڇ>��.�6̸+�\?ۉ���J�E$��}�����)Vu%�f�Zba%�T���>>��y�!"D��)��H�9N�#��_'O�ܺu��ڠ�s�S�oX�G�5�,!�-q,�~Œ���/Y���)���(�`3ZL�"�ୢ���R��8��/)���Y�Fv��}ZT''[����4��(�ĨF��f6�[����P�2Om$�~C�F��vj����0PJ q�쀶�AVJ���k���������ٿ��_�jX�I9�;^@5���!ۧ�Km~��������<���P����t>�~C ����HT#�75������+�\�F`nn�.@�𕡧������!�����!�C0aIF���"O�nP���4l�BM>-�G-��!�� ozzzvv�:otǩ��cǎ����� L�jI��~�-/��8ڲe�m,@_I^v�e#�$����3��<�}W��ظ^KBΣc�ʜV'aI ���𼚞���8�0>��xF�����f�ظ=e5���'�����j���IDg�#
�L3�Q�x�5�8p�O��j=�t)��y�I)bS�e���*})�Y�|����ï=?�G��A�2��dk� ������<��t����uu�HK®�@�$��V��'����)v��O��U�(/��mJ�;[*�h���3���hb��I�e�?����<��rMᤀ����`*ak,���Z��q4�o�UW]��s�z�llت��z�#��Ԗ�<�=2�ා~�񹹉���)|���?��0�r��!q��i��C	{���G/�����vb�Ν��{�=�>r�ȑ#�����+.�>>|v܎���.e���1�v�o���#�W���c�#����}��c����-NsA�Je�&����Ȉ�,W"W���DY���v���m�5�~���\~��[�gE��tTYd|g�p�,#�V�f5�B���X�~j�FC����ϥr��I\ u��۟��ط�=������n�[m�m���o����{���u@�����=?=l���cǮ|�k;�Fȸ�+1"�ԈI4�CE�������=��������;�p[�&_E�	* i���M�M�w��-�n�W`�S���:�Y*M�ZYq��~ ��u1MN��7�	����WH��|��^|`zv�HT� �Z.)(@��/���=_��h���PI�ˊМ�[
k��BU���e�4�,mx�Њ��8�GK!��g��EG��#�yԇa��Nt�~��$Uin�W���H�q<ϔ�e_[���R��C�DK"lK�+���V�v��J�)1�{b>�2�g��?Go�h��?�4�*�P����d��RLk����tH0�x�o
8n��a�vo��=x�K@�(��u��]��J�k������@w������&II����2�.ٌ$$@�gO�)�Хƌ
�ٵ�Ru#�%�u0�5.Z;�[cq��A�u#`!����SZXƃ�
�k)g|�":���́�gy!@1w,�ow"+�hq}����˫KA[Ca��8f(�5�&�H%�B��;��](ۨ���r�<�Nnr4�{�sSX�5�µI�a��=���YB��.��6�c�@J��'���?��}��xu 0Y L���ݶ����mۻw��L�nu����/.���1�)�y�����C,��`�v����=<q���5Ƈ�ٱ[i!l�&�Y�(va�X�d˙���5�T��!e.�r�$�۰�x�F�Ui�s�N/�u�׫ܧ%d�P9�70I�k឵otE��YEv��!��fm0\\_���l�uzaap����:�-�d�� � ��(��I�:΍y�P
)�Y�I��ih�r<N�}b�(<��( ���T^^}�H|J,H�a!Wfgb��	--�L	 �-3<����Dr���tI��uA�pTĂ����B;����Ey�*nS]���Q�5�]�M�K�E�;��
+�*���5ِ�g�	�-&�
��^�c��)�h�rw2�Z]]�'�E�6�"�<}2�� �Z_Xk��S�3��믟��YZ>y��ӋkX3AN`�=�|�/�������ݻ/�����(�[�h �<���':ޏ�z�m�����ͽ�aL�(�����a:�^���^|��o��m ���0(&J��oYX�|����od�w5��)�8������\T!�'󜥝���D,�-��4lz�L�L��\�o/b;��^�f��| �;��n����h�Ґ�����~0<x��v��V[�9M�*t���
� ��`�����=T����H�g�H�G?��W���?�3?�=H�x�����H���/}�����q��Da'����0� �|8��Xx�g]$7���]vٽ�EI������Ji�M�[V.Qe,��HWP|�flB&�,�'-ΐJ���Ƽ�^И2��؏�x���0h{��,�B�>�ģ�]�N�橫�9j�_�QU�4�t�u�֦���׌�#�6��1J���?�"�E��S�i�ի�"'c-6�s|�e1o;6�ja)��V���&�jmf�ߨ���u�B��J6�/j�H��uoʄ�Ô6�:͝��JFBk4�����w�ރ�<Ъgf���� Y�o~~>�W\q�[�=��S'A��j�4�m⼹�ئ^/�=���ihx��)��ު��O@T�r��`�8Sez4�Cy���"��X���w�ڥ�r�prr�kLOO--���B[�\h�tsQ�=��&�ڙ��zm �msf�
6�*0�SQ=(�s���;������'�s�S�N�\9s�
��K�qi&�~"�<}_X ��]��@�2��/�P�5�����;��,��p�B���L%�GƉ+�c_ǆ��q�6V�xޫ� ^xk��zmȊ�g�>�BU�᠏��1z�F���Z��I���}x��2@�1�)ͫn�}�uU}[��^М�ƪ3j�̚+��U�>��A6���jlǫ�h��_$+��� �}(����Qu�7F�!
b�a��B�̱�:SO���3U�z0E��餰tU�E� O,�\^� �zKȾ�sz
��;d6
���Y �[�l��_�O.�4�Oa���T1	3�ז����+���s�����~�t�~o4��5La�q�fgjޣ�^�Z���}VVV@�L���-_gh��-ηs�z�m:��]��_x�~~�/�o�Y;��^�&�Z�ˊ�\���r�`B�BL�1�Faț�gF�&Q
���9;�RS���������;���6�Z�e�)�LS�M���[��%�i�.����0<q���n��A�L&�H|�J��*ɢ��������[��[�����/~��J� ���m�ۯ~��?�o�����o�K92�3��Z~P�y�l��g;����èX��2NR[� Lf{�	d��N
���$�9ť֮`p(���#E���$&{�A�������C+u�)��L���FL�t��&�B&+P\K��������;�m˱���ш*]S��}{wei
k�mI�yJM��f(�H�5QT:4)!������V4�h�ʩh$F��Z�I&+3r`���r]X��4�V��}٦�)����$%�Xl9�I �[��"�^ �:�Y0Q,�ĥ ��؀8�9����X����̕��+\���K����aU�20l}G�iS��WM�+����ʵ�-�MK��Z-Pz=�i�0M0��^�k���Y<~�����w�s�Wqjl��C���G�>OM���'�{��T�2���M�L��W~;U�BtA��СPV�E� �Q�|���4Z�		C 7���i�K6|zf��r�eBc	YY���Hbn,��
�"�(L0�B��fAW�r���1 ���N2?w�^�7�	b������T�d�Y�׹�{����v��dW�)FS�X�q-Z
_hX���Z����Ed��3V��0
�ʚźjfÝRm�ߞ{�a�e+��G�Ny:Ib9���p�o)�F��k�#_��-�?Oc�#_XE�Ӭ��R7������*vJBWn�Y��
��w|�B\��$�y6==����A̩2�Bw-�Q,U&%�Q#0Q���zU+��!X>�[�V�e�Ɋa�)�_�R��R���+pӤ���M�F^����Z���h0=s�Y��s݉�Ą�5�u��0a�x�� ȢrFJWt�zAY�$g*D��S��C.=�+�EtĠoF�4����G�)��8aB3å��G�����/F�@p�0R�率���8K�ˑ8'�J��"묑ܤ���cT�	k��x��h��c�5XA��DC�k9�x���ae�Y���ea|/���7�9r���㽡��yfi	�i11���`MN��n�����K.\�t�4�o�>��_<�k���.����.��}�+_�Nu��ȧ��*��ڵ9���(�{K�̯�h��t�ʢ����0����O<����d��}�����~�W^{�֭���=z�����I?�mO'q"ű�(t#e/"9s
�@Qo�W��EۄI�%��n�z�Q߭vk��5����KY$m���uei$ݔ��o������ڗ��[n��k���αf���tT�sc��۟�饗^
Z�׿��7��m([��|8�#л�`IG���{��>�|�W~��o~�W�ΪL�я~�U?�{��7~�7?���uZn�L�� \q�K�p�l�h�^�'eIFX�GڨP�C�z���z���$aw
��e�+5nM����Ku��(B�z��'�>����<f]��	��5)�0�I���|�3W^y孷�J�M�x-�$��'>��~P��1����uV���M��dr��К}��p.X��Qڇ�9�8�)<ʶ�]��liQ��"��˚���ȅ�|-2p�Z8"怼�}�if4w���ƽ�ՎzT���l����,���fm��t��U�pF&���yl�_XXx���k�.�@�br�ă�[! ~�O�r��!f|XW�rQ�6�,3r�*�|�Sp�J�F����Úv�,�}MD�J���+Oi�"�N��\���F���СC�m���ba�<���jg\t+UD��Ӎ��N���.9ut��R�3gs��]���
� UF3-�a�z�����y�@��gڒ�c|d�w0Ol4��W�(�$}M0�dcx/���\i���Աҽ�A��?-2�+sUE��W�5#i�tL�I�S0]�6k݊�#�y�5�r~�c۾c}��v��X��	k1��g�����~e���Ż���B�GIT?����>�����\T���Cm����4��اM�R��*�g�39��H#|�_��#�,}��R�]�&7��L���0>�����mN�f'���b�k�@�~>[y��;��:����yw�ر�{n��3��9L6rї��;HS�ѫk�|Y�5�4�hG�V	X	�JN���l�T�$V��I}ʢ�O����e�I��?u��z8���8��V�˽s�����o<s�����vQ�Ge�l=��p2�}�B��v�S����εΛ��-N������X�En����AY��a)�]��]wkQ�/�����G������K��'�񎷽�X�!���Wuo���&���9p|�h�m�	��=�fk�f:�� U�P����k�\p��'��X�J[n��!zq�i����L�^$�*r���m����ͻ~��~����������%o��g�}��_��#_��k�\Sp���4�_����_��,���L;����� 	6����i���i����/`-�,�yf�x2%Y���\����m^��H)�)x)Cʻ���zӛ��b�x�O���K_Y*���$����Ç�θBbQ���[뷡�Ap�U>]���?e��tdA�F��N�8�����R�"��H,9�Q�l�$]���%�u}��P��\�r@�(,��YRƔ����(K�0++�%P]<�uHe��B�2|b�G�mEUw]��lM�[���ypK9���h��]Ob�������֙��I�b!)�O���<��a�|�5���r���k�k�T�-l�f荥��f���RI���%�fYT���&O0�l� ��vmL4��Ųd�ɋ� IF�����Z_|�NM���_����c~����-Z�0�^t����:�u��+�vƃ��#�s#.ٿk~n�^��-��6E�4~���2!��!"��,�"�	�PY�j1�DS�#�wk�"!�/d>�1Ą,����g���m���t��#}77Y��D�����R2����Uw͆��0�� E�l�۶e�T���{쳟o�L������^{�Lwzmi�nK�!��8Y8}*��\�!L��{a�HAT�D�v;
C���]>�BU9lc'�;iŠ�,3�{E��O��''�v{���׹��;�La�W^8gvf�0�#<�#�z�x�۹��d?	��³\'p�_ ,p����FCV�K�l	V8�����*}7�5���;���SS]{&��4κʲsL;t$bF���,!�fQ�� ���
%�>}�r~l�-뉣��<��-�t��/w��("֌�(�T���'*@�)2�(;�h])��sʙ$q�e�S��C�>Z(q�|; w� K42�1��Ucؕ��~+@�OAL?X�>��󵈲P���� h�`�N�B� !Úh
B��	xe�1U�vF�Z��q�0<5�a�SQ��������:c�� ��U�T���n*��0������	<&���]*۔��h?�0%�~�ٚ 5̨��~6`1�e�,X�5�%�X��5����N�<��6�y�C�[A�l��^�Ã��v��o��v���г+++�㬭��3$���:�[9� H�w���G}��Sk/{��~�����^њ��-�ή�p�閰M����;{���Ǐ���s�]?6�#8}��,,�k��?��W_�ҫ���ә,N�~|~���۬��+p<Mt��ƕ��FY�{�2�H���vЦ�>'�`%Gv�rDe�j�ϣ5X/���jr�$9�3~��Ig��#Lq�隵��wi�g� �h�%�SQ�J!�9 ��6����Ͷ����/x����U��C���?�w�D��+���[kD�R�>o���_;��^�FJێ"t��p����`IY16�B�0U����!M5 )��f���)W��/�2`AzBF�@���gIilÛ�Y�8��۾ڴ�+ ���o�6����Y#� X�����.� ez�c?�c����O~�O��O��.��Ö��o����{��4��	�2U>����/��r��(j��=46�F�r-��#��$�ߺ袋��~/hs�ms} ZY��<�^	�ؤ�c��c{X-Ķ� �	���	� �`�uܲ~q������erL,�3���|�W�ݿ�
���#�1��<� ���F�ު"� ��F���U΁j��f�Z
Ÿz����]M�J�(=<$�T�?M"�G�D1g�kIQd[��Fr�)
� �e)<����
��v5�Z8R��i0c���S=����>�H�c�~��
\C�F#&�cZ*J|R}DU���򭑧���a6!���~ি��4+F��=�x�/J�tX��|�	�Y��=�IhP��]ֶ�z�5GF#�Dn�x���T����y6�o%e(���� ��ۆ�ڵ�"�?%H�733+�!���u^��lJ�u�̉�<* 5]�Rx	bi˖--��Zl�WF�Y��vVU�BT�9ֶm�{��Ǟ�lo�֎;��n�����5��#�@����ʝ��.��R=AoWO-��G��j��/U���Re����;��D���Oy.Xnn���ȖU��I?kk����G��Va_�zEO��,��Z�CH�����%�`{�Y�P}�zC�6`�ҫ
�������^�Bs�7y�e�<ϻid6i��n��;���d��R�8�M�Wդ��s�noz�,%�s�qI�kY�H����+�`�?��c���iq�J{A���s�x�n@$�L���U�NWk����ݗ��sqq~�1��<;<e0B�꺱�a[�(��hT�b@tm����:ֲ�m�$��m��F�X��c{����?|�v�q��d0g8��+�:��,s�֠��A�2�\诌��X�!�K�D?����#�O�z��:��ý�����>d�ņ&]�)�v���i;��^��Fð=��Q<�H
���� ��r������!�pE?�w���o���da�&]���Z�>�I �ƼQ6@���w����~�z�y�滋Z>�>�=�z����я~��~��~��^����mo{�;�5c�6�+E���Cm%:Ap���|Ϗ���p��� �x�Ѡg�����!V�/�(����,J�����F���l9�!D\c0�;ej�x!���d$@h��˯��$�~� �D�B��:G?M�{��=�yOoH���	�"wl'�,�aK��W��z�;����� �����=7�G��d	��<��?����r�_u�X�+	e�)!6]p%�ҹS)�Vt�x]�����N�XJDT��~�N�W�f�R�b�0D_X�+�XD� ���ʵ=�"�ł��ӆ������L4����ٮ���o~�k�����>��O�����b��m���(���Vz*/NK+�g\T����]t�oa���"KL	'��õ�����e����9r��ɓЇ8�4�Ҍ�m04<F�0j��>5-sa���D�CO@�甝x��L�N�2�'Iη� W�О���f9�
u�3b3 ٌ֥��yj���2�Qg�^�g�X�U���Em8?����נ�� Z��N��T��*��p;1(^.�f��>�[[�В�h���p�%�335	2��"N�0(�f���gAs�t���^������K�������%�+wlݢ�n	c��#�&��dy��0d���n.
�٭�nz����9t�S�뮼r�ĩ��:j�]a{���W������O�ś_���n&}���v�~��S�7�h��1l=�Ns_�/1B����A�D�s�$��C���8�q�n��,΁�]�YaǻK 'E�XY� \������7�eN)c��ő��s�!gƙ�0T�k9��KBpK�l��8G�%�m`ж�zw�N�-��fr��iNő^�8X]�M1Ѥus^0u�ͨr���(������Eլ,�#�A��sLu'*��۾�2Z�w���6�Ʀ�p�h	�-�V���]\U	rw����1�+���+�`4�*���m�u�%�u�rC��\4Ԫ�����|��Vev�i�ȓiP�x(�.Ȥ`8�b�}F�E$=0��(|�<�����	d\GTO���tT$��B��[t�6 ������u�x�%LH��Ĝ�d塇w��}���%���+A�=}�ߚ%��*�L�<�]���P�xj�٣�"����� �r_R>����x���m�.������r3�0�\����K(X���8^�D�ğ|�}[�;6.��t�<c�V��Nm�9�T�_�f2]��[�� e�\J���Ù+<���W:��[0�3!��%I�j�i����+&�4E� ����*r���H�S nӾӴ[}���X�En����V�~��?i���"�G�����		����P�����,�/����Jpͮ/���'V�A��z�A+���l��p�o۶�-oy�'>�	�Z�����R�V�,�p�r�IpP"F��j#[;��DM���Yܶ<,m�J��n��j+�54�%���= S�xA����6���w�k�h�[��vTE�ȵ�9������N���)*%�L8�)�h ᇮۍ���/"h��o9g�鹞�4�x�f	G��,% g�(��7���>��O���!�;�)ķll�s�M�1�|�BW�z�z �^G��Hc�b���V4L���Z/�
?��h�[��O�^�� � �2���H����Ř�>���x㍠,=}��	���9��JjǱ���4�l�%�Ph>CH���d���)X��<��h4���YCؙ�Y�b�Ph�%��`�	���30��K#\9��jk���<??/��#�l:Mo�o�pPy�,k���]�M��鵨��l�#�AF�JWx���b�9��F^�eH�M���ٙhF��NR����gj��M����~�N�2q���M�v����v����+k\�luuuyy.Ȯ¢0����x�h�;��.�|<��C������p�Ç���Nx�k^�]�a�� ka�.��+�E��~���j�a��4�o�2��4{  ԡ_܇�4x�i�+-���p�虡���ƥ �V?�yZ�h4J�m깫ӄ��79]6X����#W+��Pe��\s|�,�_U�y��uZ��lǁyɓ�]�\b��F���S|�E��4�����7�n
�?ȷ��� �VK��n���2���*]湍-)͟�?��)��=Ŭ��\��sr���#G���V��2�IH�u�2�ꑇ0._G�@[���^Og��5a�8�,۷o��ںu��J�+++�	�Q��Zq)6Pj3Z-�O��)e�زe�IA j�9l=+��z������Y�e�w8����w�8,�]L��<݈p�5�o�6|�;�ҭ�{�𿦈������ �9g���%
B�����9�8>�dͩ� ��Sܵ1�+�5�2���qr�)T�/i��,M]�8�W�|���ɹ�,d�/W�y��"7C�=������CNQY�z���_��O�Ex+ƥ�"=���i&�@�A��~�8��k��#�Lbz��ہ72A�zQ�B�Ā�"߫����+W]q�����y�^@��ч�o9����f'1�L�d��Ҝj�$"��_i����5<�	<��Y����D|Y�ň�-OZӤa�@P�(Rd������n�MFUe�,J;�N��Iش��4�(���G6K����T�<I1!���� .-LX.Pׁ��{���0Щn���>|˭��馛�i|�L7�f&��s��uȎ<.�)*��R��$�,�����)]�mBE�H�ᝲ��o�I\畄E gY��m��MMK�)�}4�.��0^����$OG:Gӓ�-�������%�����s��hM��W��'�9 ±�_-������\[�	��T��k��S#�諃^{R��|�v[F��F#P ����& ��x���!�]��[��� -�F0c�M�Gp>�"B�ZIfe�9$��1�P���Y�B�? �.WRSc�/
�lF75,���+��.A�
�QcSUf|��Q& ��)�R���D�qq��I������آ��Ũ���/��Xv7�B�Q<fY�5��n�efr��Ro-���[]��ޚ�F�h ��\�ff���C��];w�����W���'����wb��Jo�����dGy�:����ű��3)�z_3m2C�fv� ��55��^9��s�ζ����������嵷�Wzao��}&���[���կ9�:�p��Q�Ïbw�T�����J��XS�pr��E�����;� �k�w�0�`X��J}�[��F�}t�p�NB�x����#y䘹�����)g�oBX	�!k��@!�*�!� ��5��@B��h���M�~�@��פ�5���镕)Daf �L��B&��Hi�U+�Pk�NC�G�����e��@ 5����`չ��]�gܪ�X]}")9��MK���U�2��O�s��lg�D��&ˉ�c���/��VCeR�*�w��D��r8z](�˥ z�G=uIz�MDJ����?͸30/�|��Gdb��j<97����"�Y�<ey�_T��s�@1: �V�M���0'fSľ��랤�W�p�L�)��7�禅s��P�h���LK��cE�<�½�{E$�:)�ȳЧ�H��U�N�{^�H�R[Jd���fp�j�16�G�W�j�!��H<�=��Tm�:�-�R�@��R|��o�m��G;����,��,��0�˾�a��C������)�Xt�8���Β�[��8�Ps#���gS뽌��rE� ��g�|ߴ�X�En�J�	��r�
�hȯ��y�J�c9��=�쑓㕯����,e�I������y���x��mgi�xtK:�������Is����>��׽���{���l~�{=)Q��=�� �w��'1���`�Ad.�@O�4ڎ�!�f?51�C���@�II@O�����%�!?��(z.�zax�
�wC�O�G�<+�(Rrp����.��THyq0ҚXD��6|y-��9��Q$�i�e�0ټ��.�_~��N�8�/|���^��\;��%kʗe8Ym+j��<��
?˹�W�Aul�+��ï�w�y2E��у�*H���K0���p�z��=���I�=��㧞:������B�t�}����ǎ�K���]}���"=??�0���|�E�t����Ҧ<�J�&�V����l��T�@1w�Ŝ1Ї�������+A�ĥ��Z���#�8bAT�](�S4壘|��2���Udř�<
1����R~�
��x��8٥t/0�u�aϡ��1OFU�x��Q����XԚ��v�y����?�f�I�����y����Z&'�xS�u����f8�חa/+���aN�C��ģKKG��tt���OOcy�h -�y�����
&f��Ӭ"c�%�~>Jqכ�	rK�
�郋?����� v`�9�1�F��m�ݶu�֏��G�ݺ�837{��wo���5F�>�j��p8����|�BV\���0ƕbK�*�65Ӆ�O�6R��1�d'	�(�Ŕ{J�	-�UX�к��n�<e%.M�]�I٪�N��ƚ�k�cA4�Y#��(3�3=Zuc۰�H&9g��0�-+Йh�&F	&QTiZ��>y�]v�m���g|�4�L�}���n̋���jv��}��XZ$+�
˫��{M�/a����r��;t�,�'�x"79�;z-���U�'��z�Îa�y��R��L����_���/>@��
�	�o��
~�ܽ{7\>����?���`��ĐG��D1A����رcrr�/[��1V��6K����x5�`Bؤu�Φ��z �Q�C[)���&����狼R��Aq.y"H�0Ъ�N��W��=�Ri�9?�4z�.h�ˮ0v[1�,g0Z�.��C c�E�#����e7D)>7���&�2��n�f��]��tm��Z/v�h��Lb� ]8yH3
[�\d��1+2�iRPLE!����D `����vg�(�w��e'i���EIX%�H�D�i���2��K�·1C馛���u#\An&S]����P�[i�	
�#�6 �,����.�efDn�4C��0��*F
��9L鸄 �������(�0�HY&1x^�@��S"�n&L��0�|��E^�m�)�-$u�Dl�$o�-��D��WH��� -;NR������H5N�g!�U=�-����ɷ��]���0��²�d��������Rk��#6�MU�E�Z�0s5%FUKTIY�=l��0�q�K�?��f!�b�#.S`P�ﶶL�Q���tTx��x�Keu��0F�H�ht���_��(�2�f¹`߮������2���-i�{/p���o<�>��������0^Y\b-�I���jz��˔ToǶ*zP��-��΃��h5�ĎB��k�%�=��EV|M�pNL��K�%��k����80e� �[�K��eC']R���8�]D�ke�o��Y7j`�a^h�Y�+����k�G�ekV��M��%^:S��`h8� 6%��O�(�څe{��l҆�b;�iLꝶ��EY��	��Ջ�ՕޓO=�:S]hā�#+�Ó��Y�L2����Tw��^\8����l=��!��� ,�3=����k��fg�"��g11 j����|�!l���%��=щ�@���Lt��%#V��ն<����������8N��gQ�O����y��-X8a*���L"��0��?���ay8�-_i�h/�q�he,o�巕7m�l��0v3Ӳ�ǋ��E�A�Ջ-����q�����m[��YHt<g�2Xs%�pmS�4C뵂3N)���G�UV��.��B����v�DYb�6��O)�,�Q���S�5�hO�V�c����:q	�Z��w8�?R��d��D�[���ht�K?U��hQ���ǨrK�m���c�|��nX��O�[��tX~����Z�E�J����+lx���b�k*�\G{�����am$��1DE��թ�����s�= �ca���mn��j=s�Y�٭�Hda�E
��M&�?�o������:;�(X���0N�yR�;�q�,�V�n�[���yά�jgJ�� ��
벤�1߆��'w?J
e�0Һ�H�)����l���?�Z 	���a���^��1���3u�f��k��'9��K�@�\!]#��U�?�^�VgX��Eo�]QíMƅM�&O�KQ�VV�j�D5y�A��F�б; ����eX�̠C6Č��������9�.��
hZ��b|H4�Ӵ�hp`a�o�Q��,q	4s��A�C���7��{���Z/v��k�!I��3TS�L��.]j�lG��,�-ZmY��V_���&�#��D�A��{��e�n��%}�(+�%+�x
.II�b1"�y�����c������Ж\�%��/������m x&��Zfy�3���ƀj(P�X��T:&�hUE�
�i�_��O�����^/���s8�<U�C��k��&2b(���o- Z�(6����5�t��/ ��h���5a�d�q�Z�����Ҵ�?�{���ł���:|Ɗ�Sߌ�iL/�kQEB'��-Ś�+l�f���E�?��d���6$�+Gf��ĕ:Y�E��عs�-[���	O��Ϯ����<ug����C
xI�.�Ny����v�K.�d$�ѣG��͕*�z���믿�s����В7F>��#��kE�U���ߜ��܃��KQ��ZU���7�<����橮+|�i�qV	�u����kG�4�%XCA{����4�"�S�4��F�mc�2$��-(ˮ5�b�y��ڻP�_�*|��u,b#��\gF�_w���!�U-2�Ȣ��8%7ڟ���CB��g��x�|��lꙞ�����9x��+`�Lat���/Y��~��a��#V��7Ng�>�XPR���7�Y��	Ð/�g��H��{�8p�_��_/,,��I����zpSX`p��a�7~�7�n���7���>�����mO�t#7����\phs��(����n�y/���u��h���`ev��h����k!^��@&�!e������0�Ȏ�G��Ce~Eb��]-��\!J|C�3F6t,b�?���t������+�Ȃ0A'�MMua:`a.���_���~��k�:^Sl$�h��Y3g���8�l샭:6ΏU�l�)/D��E5ʝK�YB�Q�Jr�ye9^����~�-�Xr[�n-z�a��O`�j����s�ZH@F�J���O--.--]������W���>��ţ�TK}mղľ}������~+�2k`�aR`vVS�w�6����we�����/���;�|�/?��L�Y�����j�\��^�w�����/�ҌV�jH���o~�t���[��Q� �J���6�e��V�D�;�z����ٔ�I۴�(_����ƃ�B]�\U���9��/�`&-�"n��&X��9e�����?Mh�d��җ�t��7�����w�qo؊�]�3��r_�����?��;��0��v�N��~l�֋ܴ�$Z�� �N��� 	Ji�.�L�e<Cl�2� 2������HC���[��X�IbRM�1$�m�pz2�J;h+��-�B�F�[b����)B�R�;T�o
�j3��F#���vМ��w�,�ob��o���=���	*�+@/� r���hl��)|�/¥��w�q�:��	���d�ÆC���d��'[a4��,�ɇ�ĤY�"|BǠ�Z��i��P��G˹�Ȍ��X��&8VQ�Y[p8&q���A�c'��y��/E�J䦩��Uz]$�ї����z[�B"�� �g¡Jr�*k,��\��*=��yV�����
�#Wҁvd�C�@��"T�y4�)�2��eZdE'�[��\�
���{�+Gc����3XX��x��������t܉����ڱ�m���ݶ
��Gnnϵ/���L��n��k{l�6���
�Uf�#f�:BynS�������<L%tl�|ۏs@�"Y��\��ҔM5�
�0�O-��{p8�UA��Fnr�2B
��ӧt�Q
�eeL(B��$�3�Ѝ5�m��� ��qz���s��VĔ�%l	��F��ub�D�����6B+1Q��Md��FQ�&c�}�P��N��r"�Q(K9q݂:�ڙ$mo�8�-1�)ɐ3ݿ`^�f��-�ɆY�1k��z}�v|��[hҞ��lQj"M}#�������"G6�x���t2������3a�8�#upB4	0T��I��[a���������tt��E��߳{�����N��I��-�?��`]~�%�w�~�����_r�4��sځ��`���������R"��X.�HG|:�M��=��X
�ڢ ���Lőg�W�'0��jGR9*\��5�4��
�Z�'õ�J�S�i��q�+�0v�9�+��9ig�;�N�;)��*�B�oA�~oPS(�J�d,����� ��rQ:� .���-(�fPĬ��oY�Kh��/e�UŎQ+"�Z����F� ���agyf��3���=��8���v0b-�4� �)�q�ThT(6��ǃ�9�a�%U�*�L��@W�Ќ�,/J���*�腂��6�|�&�b6ճ��K*��e�C�iJȱ͂.^`���ʒ��R�x�.8.�T��`bk�w.�v L-�*�DHGQ�1�i���2ۙ�x9�3$h-
mEI���$��ن��Ȓ<-wJz8��J��}�o��ٵgW��뽕��:<�J��DLNں������؃��{lu�ζX��ֻ3vǟ��e��8�I����}���9���f}A�S7���6;9?מ�ھk���BS�e���>f&�ݞ���'�U�R�G�sBF�D�U��T҂b�H����[%暿G��?�&7J|��i����VU�)���4�a���rU@n��1}��+�y�L���p@�����o��΂���Z�uϒ�H_������Ї~�e��Wm�$~���s��\d���,����������W���J;�(w2�T�X�؁�X����)�LaB8@7�	����ᣧO�JDRP��"I��Ժ�>��uk��-I�b;t3�R1��x�h���Tv�X���?�Wi��]��󻘌+�3Єj�4SE�(*W����p�J���
�8A���l��i�v�tt�k����J��ˎ���!�ci�AoE�n���~i�4��n�4IZ�l�0�X^��d&�hc;t��Vc�;�NV`��D�2����0 ��=Ԇ��d��Fp��_�"z�
RD����8��@�Ѧ�;��d�d���N^�*��@�n�yA|*�UG�f����B:��4CFT8W�?��%�Q^U�l
\]�ˡ�#��?�C?t�Kn��Z^[g�>D�ah���׾��œ�N�>�Tؾ���?}�i�G=L�A5GH��=��SSS��Ӡ�H"=��0h�/yپ[n�E�{��O?�t'ˎ;��x:I�8qbۖ�pM�p?�,��*Q���rTDUXLU�@VU��K�t[H0������F����̲��.K�%�0����Z�\6
g�q��{�D-�'h6�!3;;:
��Ă��;DA�_e3�� �Z۫��T)9��PW�ڤ��6W�ơ�<���᫪��9��BZ]���+��i��2��M0bp�Nx=��������?�/_\\\:zV<��(ܿ���Ҷm�zq���㹋��"${�Fʒ'�|r�PG�ݻwo�׋c��n�a1%@N��v��I).n�?��?�����k�������}�eU����ƪꪮ���MGZ�&0���!�2b@d@�qTD�cB���錱����π>��IM�P�+�prx�_��S����1�{�����Tݺ��s��{��_�_��;66V�������ʕ+��*ͥ���$ٵv�Z�;B�_�җ�nݺu�K��z"�M��K�U4�^.dUEh�`�E��~���$�T)U�lN��Y���p[�M�2�?;8{a��X�H�ز��M:�Z4���'��}M[#��~[4��k�Sc�k���C�Q�D����?�ec��󈟋\�Ü�1{�lZ�d8,��H�U3��͡�
�z�kIm%j�(�?�=0(=V(�y!M���8͇�n����ԉZ��R��s�~7���_�b����-����E��x��e�mI��6!3Ŝ�,2��+��)�m6�lCl�iV'�%�elbe�����;���㏿��o>��K�,9���ךP{+���z{{�͛�q�F��[o�	�u�p$���e�^@&6qmb��{�ݵ����:�s���w�ܲy�fY��O�>s���˗w���m������{�9��Eۤ�O�6M$�I�T��q�����R
iKh�����v��O�v[�����VK.�[���p���yD��P�����������P��~������t�Gz�7s�מx�G>W��?��O��/�߱sF�8v	q]��+������>���^�3��i4�V'�:�X_כ�~br�<���S�?���7��DQ�0(hK�Ԇ��걏k�ʇ �1kh�ALLB8'
U�����<#!?5� &�CeI��	�;�D�#)Pt�14COU��
e"��&aRP�4&[*� �3ȫ'F�#�@KA��ح"�<¨���lÔ�4��Z$�e@�#�h��N�*x^ �7E�S�	B��V5�H��:-$z���jr��h�l�J!A�0PܥiVq[����#�Y��,+�HV{U"��F��s,��YB�ĸA�����],'��LL�*N}\64۲��GMu��~�O�U�|/�zKSu�@&�bӲ"�D\�yzm�M	
]�'���*�7:�`<��Lu-�r���s��ӑ���
����tY��jl��Ḳ��Hn���R���a��7(�3h�B������N]M	s�b�E��L6�F$G�^��=a�o�`*J��U��K��&��5�<�͘�h�����@ʹY-�����\¬	�i "?1T��u��Tv;h�۴:��}�0�Ϗh�pF8=)C�i��o�8�t��
�ߖ����ω�;f����`�zc�ņn�<�|p� d���Bp��*�61�	�D���=rK�=��*Œ�ދ������3ì&mKr��I�&D$w�.��w�3�+]0+Y�S0%<��.ۡe����W`�M%M�PWF�4�Ԉ'���Y͆F�1�Lq�j�~===Ƭnw�ذ�Biɒe��^PWw��(�%b_�ƣǋ�����|�š�z�׉�yI�hI)��E'"�11>:4�0�a�o4�TP�J��z
�lH���R�V�v�۩�����[�*ֳ[�l߲=��PU5Y7�xצ���\��ؼy^__ٲp@�k�|b{�v7p�υ�4k�ұU�9G�A�zJa
%�*TM�{K�b��FnB�:T�@�@���&A�-��c��j!n�W:qme�uZ`G�km��f�J�bK�*���U�>C��~բ��fä�M��@uV�l2`���%hI"<L�ł�b��*���$�[ 7�N�)1�w�m���@e9����R����M�ҍ�J�XU�T.Xvs��@�3����F�H�@��e]��l�x��*�j��@��w�˭n����C&DƁl��ճߡMD?{L�I��N��x�Po���L��GA�GD�?ZV3f�(,�`�� KE�;�Yn!g�
���T%��[
������J���j�k��G�dcҀ%ӍB�.k�^kx�͜9�oFς�s�z͝;.�F�u�Zcrx�6n�N_�,2d�S�	"K�z��q��T��C#��z��٭��~K�wt���w�O��j�=��/�t�m��@ғ����K͠]ex�`R��4���&��A���"�����X(�ܣn���BCBx
</X�m.W)T[-��n���U�ȾrLez���?O/�[�Z�d��%\d?�����?��{q�q��(٣|�k����������Z��l(Q�|�+_"3���߸����P�Eڡa��9�NW��Rp;YP�'��o~��ȇz�o�|J�$YͫѤ�걏k��`(g����6�d��B�3�g�:A�EAn����	pNG�X��ьz�^�m8�<_F��վ �
�R�
zp��,@`���q ����A;�uo�
�vὓ����\OC�в(qV�"g]��R޹��q�%/� ���J��Sc���X��x[�羀z�M %s�y�p� �Թ�Ka�E1�h���9�|⬅r���{��HQ»u���Ϛ�	M����/uE��a��zS��!n�V6Z��Lp��I�s����-0�oI��Ș�1=+���?'�p>:H)�4F�=IBf 
�����l��U��1��pUl��8N`�,�'�x��ٳ	�u�7o�����j�&�o����]t����w�,Y���S�]Z�h�H=��������?ޜY��z{{''���	��d<�e����2�X����C��i:���_E��j#�"�N�Bh8�"��}�@������e���E�a�2D��t��c����Ǘ�.�d(J��*gU��Q�[9ZR��ۑ���ٿ�i��p^����
��^1L�0��.�.Pu�'�Y>��G�L+���F�G8�9�j�	=�Y���͛�[���֭��w�q�?�'�[�n���{ۂ����?Q۾}�-���z�;�ժ�&��\U2��%����6�'p#:��
i"�-�xZ�������ڵk˝����^ӣ'��3�<�f͚���[etxa�zt1��Y�x�4�B��+�(�&jF�j��O�x���ԃxP�(r���-2��NjE0�ߘ�N��Ƚ�c�4�z���W�&�rK�D��Z˩ ?4�|�G���8N��_e|o�)���=���/���!�����V�~#Y�'L3�A�K�.�IBF���m���ĸk�0тr�}%{��>��/���N��x2,S�Hѧ.?�(9E(KN��ߩ'���"1O���Z�%軨��o�[޾}����}��Gka֬Y�V��ɉW>��?���gi��yP��y�"E�G(T��%BӲ��8
+��045D�E���lZs���'�G�2ܸq#=v��lٲ���>hmvU���M��4Q�(z[r�=WH����O8�MozӢ�s鄮�1+���q��/~�'sm��fM���[����l/~knYz9C������:�6	�U�"�*�5��2���{{:�-��d�U9b_(�¼���5-@��w�����n	r���ӟ����UW]E�(��#�5M�����o��~��6�B.Ub�BCt���4'���/�5���q�w>����CG���Y���ﱏk��Ӓ�0V^����ޯ}�I'�N�t��n�#�����[�����|9%���w��G>��8��;���λ@B,֌h��3Y�y�-daS��z�%@V�,=��#&��4$��1eC��w�����.=�|'!�3�8��n����㢩I	��3�X���}�t��������DI�4�%g�y�]?����o��淝���K���b`
�[a��ʴ"
˖�ؼy��h��:`�c�=F��� ��j4˗/ڱ+Vx�<��q�*w˕D�aʁWS,+��ޙ}���F�Q�z�A�����
6{f��*I���-���y�o}�7�����z��&�"��[���|��"Bg�=�� �
$�r�ƈ-�W��p�@c26�����V]1�G���+ F������4	�]��j���E����.���	�gww7|�)LU$��b�V�Zit�z���;.�cq��6j���,�j�]�:�r(M3�^P(�u�%�e�=��Vz:��;g/_<{��R G����]OoX��ڶ	B�s�f:�����P� +M��� �֯�S����D���T\���F�zq0ٜ
슩�ܬ��r�f~�T�fI���!ZhYĮ�g�F״��2F���с*��[~Lȼ���4�UB$���Y<�l��w\�d�j����k�Pֵ`txH�.���|�]�wC�b��E� �d��}��U���� �Vq���[|K�;�0ˤaw5x.�� ���S��w���I���SZ��+���A7N������Vw�tvWKr��;�a���NZ�/����|�
������ K���ܨ����ڬ��OۨnZ�m�|����E�ߨ��_"�Y��h4���MmbBC;V�fY��7���]�Ν�^��Ǝ?>)є���z����S��@ȵѐ��`~�b��s��U-S	����@_�J�P�t�z�h�o�`eǐ�d��J{P�=�-z)�� �kV�f�x�2x�w�h'�%��ɑ��XL�r�*���D�ډ�<S�oA�u)91M�щP�\�Ҙ:%���q�*�m�*q�qvE�U�݉���p���ٻ�r~Ә��729D�˭!���q�Y�f�d����i�s�F���+Nｐ��
�I�;)�WF���@lj�LӖDM�W�%��\����/�:��S��ml�T��"&mͲ����A�i�4�ġ���T�4Eh�*8�5���c.�lP[�rE����SY�*��7]7;EZ~�k�}א�6�wZ]C��S�PT]�n������]�`��R�Bkjttr׮]I�ڴ;�uΜ91Ye�Y+Ul�ݦ�}D�ØyZ�O/Լ������0�wڱ��Q)ӕ7΋/�X�9`�.�܉���3z�tԆ�@&岥G��Fa�oںukĳN(@�Iʫ%���h��k�?r���uҪ��A���ۜwIY�T�1ۉ�g�M�M�8�.]�x�����-Fǩg�F��`U=DDwZ��I(�A��ƭj�k��vi/H㕴�m����,p���L����x����2QM-J���}��><k2���Xd�q_
�{��Z��Ad��1���f��%�}�|�ӟ��k[���~����ÚA�4��Y�i�y�w�G��Z�E���-j�0A�]8BlΜ9<����W[�.�¯V��sC�%�|��|�#��!�^���m�w�y�-��%�_~����"��68r�GO��4��'�|���op`4f�Q�׈�m�:�+j�t�]�z�eW_r饗6z�Q$~����aÆ�>�^C������3�L�>}�����%s�͇tp��0u�|�N�֭#�=��i�Ǡ,��<2��-[�:��	�@<�d��:���I�(f*=j�y����j��R:����:��o��뮸�L�K��N��n#����0�MmW���2�5
1����
�e�rG09��@�7m�$����@�x8��t+J�0�r�f�~"##�'����6l���ۏ'ʴ��%�J� ��O���e$���+
~��[z��=�X�3�Ð&+�iv�ܹ��]�>�����h6����=��n��=i�$�"�r/�X�Il�Q�E9�ɻ����0�@c�3��R�{D�W�\I���(��-�:�jn�uc�w��Z���|v�DG���_�U�7c&=��#�����Pj���Uv�R����A�+L�����)JK�n��?ڣ���Gp�<�B�)MS��9���7���2}��<PC���J�&�222�g�Xt�4���͛7�[�q�&͟?W�t��u��47j��Z-��	Z�Lw �YE4E���ɻ��t�7F�dLظ�����>k�4\�uے;v�%D�`7	Q��^�u��ͦ�ۚ��z��g��mC �'��x&NM�ӄwt�W��浕%�E0AV�����#�2�vS?�*�ڇ:�-��WZ����J��8c\t����v�����^��7ii�9��yy�Ȯ���3S��E����0�2	��\�?�h6�g�~�eKܵ��{��O-��/;�I�ݶ���q-^YQ�w�ן�7ptH�ީ��/jw��ۥ�.��"ZN�P��{zz���7�|�D�H������9�̵��:E�'N��OXlV�������ɆGk�ib����aF	v�00���իW��1��S�����E�Y�hޕ�w)�)�N��ӧ��Q�h��a�|Q/8�c���)⁴����Y2�k�t��{gs�A��~�v�a���y��x���嫣������{G�:lJjMB@J�
��+g
�ڪ���Y2�Aw� �IG}�?��?~��מy֙�a5#���/�{���WG�臘ي�v�ڹs�V�EN���D63�~j�IyGC-|71��K4��݈`C9EMY�Vp���e�ѥm�.���~���֫|��j�T�����ӗ^~E���C��Kr���ں��}䱒��r��7�|��������<���������>����P�Q���5s�����5�̽�(}�c�^���}�����"B �E�Z2�q�ݬ>|�����hZ��o��ۊh?E�#��⋿z�7��͝q��gӮ��'.�����՟��h��6hy�~�yw�}��g����ݑ��m���?0xƙo��m�Hbi��m�r������~��=1Ti}�F�e�9���?�l�]v��>�yQ�x�I'�{��}�~v���F�O\V���\r�箸�m�r�����~w�~��[m�,BJ2��Y����6�O_q��W]��X���v�������;�C.Wb��W	�+.�����X�8����������<��_�q�u$x %{�C�M�Ч$Mt B����14��V�((�噥�dڴa���i�Hj�a�N֌T%V}� ��L�G��7W$�>��m{~�z��
� g���Hk$�ê�J�#�P3K��Uz�8c��<��	$�\0;-��=����.�n�Bݞ;i�v��oE��66���է�X��E��z��A��vvT�b\���Jwg'���F]\���[�S�rq���.@1�[4�0&�K.��F��CU4P�v� �%S���
e���=?��JJ󊆩Q������ݖ�<� 
$1�bQ�ø{ڴr�D\1�GFc1Vt���j��y	\�
�M(�����a���[ܗ�A9��GnK �Z�\���?d���؋�i�a2EL^���Fc�ϊS�l��J7r>C��I7NvL����W)�ǟr�y�=�}9���,���gB��T�Β5��B|���=�.���f��)M����X-h�5�d�����w���k�j૖��{��҂j�R�������좙Y�ࡘd�ԇ��h���7�?0m�4b���J�w+J¦*����j�`?F �X�8�7�*zB�	¬^}O,B�K��fVQ��5E����Řdy��έ��D����|�'
@��-��C\:Mq�*e�$����"�o�0�o�Di��1�h��H���լ_<5�2B��,�)��C�=BK�[�S9F���(u���E��;v
'��(��vq�j ��9�p�h�=��������u�M _�k)��i�e��i�寴Þ�,���{�C>?�v��8�q8I]p�TIi�̸�;H�Mh2�24�Q��5�a�R��&�~A��2бb"�1�s� ��lnݲ����q�^��х��2�-�����%���(��?�q�k�;w�TT�,�\��G��?X&���Ih�V:�[��Ga�U�sk�Xta��݈�Dv��s9�����AL�F�.w�7��>�1t�F>4��(�շ}���;1���%�5�����ޱ��6��>��0P����!�eӉi&�Xy�,�c/�%ND�O�YA'���k�%ڳ�]_��/����<��!�f����"�z�e�}���H�LԜ�l�EZ���{I�X)�a��'��0���.�k'A��Z����D���u�Ή�1:dǱƾQ�0b�1\7$4�H��k��ǵ^��fO�*5!Kz�M7]w�u�![‏~�)������o|�;ߩ�J����0 �466v�;κ���y�C=�s��@�WΒ�St|S��m~�s�{i�����O��n�J�nOAՆ
{�t>��к���~��#��z �a|�+_���t�A���N;�4�����'W�Z���vx�;Vѕ�^���GnvMO~��t�7Xp]o޼������ƍ�_�R4�Cї���ڵk>�@�v\�e����bŊ�{lxd�X,�������+�h�����o_���x����B�9�L���J����,���Kױ$4�#�E�7���j]�
!B���[����G���v�r�!��t�ҿ����W�z���(}{�q�L֫L�р��h�lHSq����(�	�D��A�� J^(�)o�I��a֬Y�F����p������뽱����"W.E:�:K�����9�зp.v�ƸȖ��g��Y�7vu�"�T�uß^�[��n5%�6}�t�UC�M�>11AS���S?g\��KD�hK}Ƅw<a��L�*W�{EIKb^ӈ\A?˳+4�����py9}jѢE�;Itʣ˖�A��wǳm���X4eIJ0��!:�F��B�"NY� ݣ�V�b��v���v����SJt�2�3�S�-=� �E��%+�kA����1��������i�:Z�����������*K&Xz��p��t���/����%iUm�̙�����-[�mt*�?ĵ�=�C��X����
|��j*jY����u _q��X�"NV�S����K@��f�XA����om2p������'a��֐�M��LMTQ������݌�:7a}�诂��\N��$�Ե$�v�G�%�M,e>��hsۛ���l��gK���bbUo��6B޾^v�eJ�.4K�i���#���x��
e3�G�'��0�v��(��A������6�N�0�5�����k���
��`�����޷)�<Sb�f����SiOd�����<�(�4BD��lM��=��V��th���*�����O j}�*��&B[m�����N���0� �9�HZM>gv���N�^t �J6?�`�l�͛G^�Ҿ08:`���O>ĖE�`��ү%JwD�9�+Ґ�!���Z����\���&�v�u��dd���]�!.�o�7o޼}��L�Xj5��}��6�m3\�o�_��x�C����\uPl����t��s#;�Zc����i��~�ι�{ǏL/�9�������j��
A�����p- �	�VȽU���Sn����P͈��(0Z�Ś���{��9�}9����� �+	�����6��7�5ܚr���7�<6<r��W�~�;��Z���F�}��K.ۺ}�ʕ��˰�T�� zq)YmYOt�ؽ6k�෿�4�pJڌlݰeC��!R��o�qÎ�}��G{u�+�EZ���v��k>���~�K_��'?}�Y�X��s�i�	���;�G��l��0�R�[n�-���*,�A�K�D�m\�UtHz����7�`�w�}Ҿ�:+V.~��'��U�֦���L�ԗPO�z�h�"⇪b��dk�*�Rj{�k����w�.�(�̅�q�-[�t��@!����9�������S�����أ���!�>�<D���3�?�������h�Q�C H�2Z�ə�[�҈���G)�\�v�����Q S�Ԫи4�֤�Fj��Jh�#S��tR(�<��~O_�robB�;���^�k{���p�p�+(Zm$A�R��E���I��^���\1F�v �`�v���b�������h���v���_����߾�d�d�U4��gљJ�x���H�.̙��L^ae�������*�?I�?5��M����pMa�e�@�a̸VWT}eME�,����OK -|Ё�<�f;���d��`TK�FG���ס�a��Fy��&�:4� 	H�v�a4'���y��j([�*Xn���r��R��T�^b�γ�,�hvL��&�[�^d�AF�MA�ۆ�T��S��$�*w��f��"- X�;x,�L�2|����ڭ��3[h8���S>1kf�쎎MNNڍ��X�n��FZ�XQ�WGQY:���vw�m'�)�m�Ӧ�����{ʉ6n�h�U��q�0�f��-%p�n�ZP���M `�."!ǝ��](����b�ʥ��'w��>C����{f��M�A}2Q��B�oT���e�S�=��:M1Q�%�����2V�,A�-���F���cEUhX�q!�U�L�q�<�#��,�Ȁ;��$b9��)���;~)�ْ���T�|\���NX'�t4�F�S�>�t��Hh�s͸��"���J�n�)J��l�H-11KM�l�s�~�cd���h����B��d����k�n�Ӳ��HZQu�AH��b���x��YnْoL�`F�-����*�Z����m��,,�RK?MHS�Ύ|Ew�խ��Wi�h���+9�mu�N��R�8�O���R�T�����Q��)����I�Mj)��-]SD�@��ʺR��t��ND�`�!�I)W:�x6�Д4ϫ��Ac$͞;����N�^@�?ኯF��,�ju�7�
J�<�c��t����"twg[h2eIcu%x(ƚ���8-n�Ԕʈ���E�5ϛ3w������/~qW$��x�A�L�%k�Mg�.�;/K����PFZZ"�F<�T�N��x�)�������Km>�4k(��1��J0�v�C�J!U��~p*����+�Y"Q���,Dt��5;Un�e����]���#���_���tB��x��p|�`�B�:�Y➏�a�!�Qx�X���tMgâ�f�R"��!sEb`)�rk�]�1����i/��k��ǵ^�[��8Qd��뮷��-���R�F�`��O�yꩧ
�IӉe�.udX?��'�xB�va�D�	!�&�~U����q��)�I�Z�TL/������鯧�v�G�ƲSΓ�3L8&���7���ԋ/�����6-��%^�Z���nݺ�?�T2Ð�l��Y����<��sW��n��4�����ī"�<�*B$��cEˢ��4����o|�Y3\'6M�d�}�H|ڙ�vmb� ��'���U��C�R��.W*R�]0�F�<�	<@�W}ꩧ�==�$J��f������׿��{�}LP��t���!`r�G
��/yЁ鱤j,���a��E	ז�_�ٌF�8�Ν;����G^�6-ͮ�vN����䤄�f�xbt�B�	M�P���o��qӌ3D�+A�N8aVw/!��Б�@_��"�MIwww=�j�F�M!{Hd42 =.�+s��U��F(v�n�7�ٳgϙ3g۶mCc������B�ԡ"B=�)%ܺ��-K��.?�I�K�D��w��g��'k"�Ĳ/���	q9�7 ������ر����7tf��b2�A~�n!�L<=��������O�F�,�$`�lD90���-Q��P_l��,��
��J�_k9�v�59�fk���,bs#[G��iм��5+D,1�8�)�^�&i뱋�Yod'�ך�C��@;,�s\p��T#�6m޼�'�QxǇ�ڳ�>[j�w\��AL;U0��n߾}�<hl���y"
�(H�P(7k�*�!��@(���+7K�� ���J6%�d,�c��s}IƋZp-�˂ke�NdpN]^��b�m����e�&�X��U؞��
%PwA������Yxm%��c�c��k��I���4�Q�f�:��װ9����Ԅ<��l�D�k����W��i!�ǩ��f�H�lV�<��0Ey��-�������@*"�+�Ă�B�RbCWK�!S?ʻ��_Y�V$5���yDVH��\�y
�ޱ�Wx�T��Z��#%5���;��5lS_̿1�1�	��ƴ��^h����eV �W&�/�6�V�`����NuUR4�CCC�C(�������ҬDfo�N�W��/��Ak�R�´6=q��D(V� ��L��Cƺ��4�67S|;]�9��%>1>B'�M�H�^�{��53�7� ]AG��K�ƵV�����J͘�GOH�˖����������+-��'�X�"j��+��!eu�YoR���_��.�����C��pl�N%�K�,��o~��e��`��Z����o�[�~4o�ן���?�0�U��8��H��[��۱�&���L]J��24PY!JQ��Ś�5�:څ�R�o�3�m�r�ז�`���k��G��X)�����&[�b�*h�%�]����έ�h�͜1qʄ� �Y�0
}MOЉ�H�7����G�2�VEZ���K.�į���:��4��B�R��V��X��'7��ƭ�e=���%����D(����O45��頩O�a�D�������yM�^d��5k���暯!_F5�8��탷�v�y睧������� >(	-�k���(,i��SS|�\�xen�����;?s�ۓ0.�*�9RC�#�Ջ��?���۶n���88[W��=�� �5��,��F�a٪eZA����k6�o��׮�c4�������?���fΙ'%��,<���j�A���͛���c�������إj�˖�&_ަ5��C�*���s�Ǎ��I�D�H]��<>M�I3*6�"�oY�K���^/$0��������܅9�U���Z:��"��qjO� �3�lNԜTBׂ�Y�GD�R]Ö�����[��A��w�����e�nx�0�mEi�S�,���d���uU���e�Z��� .$�I�ȓ!���8�(r7�0$ԯ��[ ��u���:��@�a��x��UK�M!�A#���%�$�k�o���?w)���Pip48�yoW��࣫����̪bR,#$���!��>��bWt0y�Kf�t�-]�G�f�(��s-�Ya�E5���#��=2aA���>{��!m�bH5�uIQ��D���3)SL�"�V���6j�C�UQm�	N��X�$�`�Q"0D�U88�q�P�iZ���R(��L/�嗀�6$Mv�5�Ї?i�?���Q%�m��'�kr�X����;��q�1�=�Z��F^!�I�����;f'��Wh��K���u��P;G�0�Q�c�AH�_U�J��F�P�"M�����	h����I��<W�H��%���F%�:"���@{<�̯褒$"^��IH����Tt�^��,eX�z:�8�e���,k��p���x�i6�X��D�j��&�B���*���id/N-Y-�@MUn�.�:OM@W�R��#�"+�W6N�7g�7��a%D��`*v��rV��j��+V��C3
��d��-�� C@(U�	g�-��-1J(��:�i5�.B��x"�L�)�|�jɐ3()�����v0zSXbG�Z����������f��DD(
@�C�|P8���ď�%�~�;�r3�L�P� �����&Z�D����h��eY˰�cj��� bZ7���̬�T7lAz��V�-����]�P�C���V%�@̒�1-�f�H�� JO�%J"WN��O9��#h�6��� �R�D�f��;�<��ܻ��͙]. �{v��͎��!I��I��ѷ�	����DV�k��?�&�'���H��{"V�x�P��WP�#�k�!���P8@�O'��P;��~�㟼�����<aB��JƏ�a���W��h~��w���o\�O����c����u.��˯ں���+>].U�lЌ#reL7�*h�k�.�j��s6haE�L�\ �Z ��͎�_Iy�Ψ}\�U>������ƍ�.\�P�h�Ԛn� IO=�ԪU� ��+Di,^Ew�����;?�r��C�oz�wܡ��7�yֻ"�4�K\��(g,v���G>"��E��E�\��f���Or�!P-����W�Ր�����C���D����hl�H0֮]{�\}�է�zBJȩ ��D"� qi��G��C��h��Ih�6\[���]�K/�t���������2 f|�=H����?������g�I��4$�F@;� ��?�b\R 0}D�<�r�I���H���/^|�駻����(軠�����g͚����9���b�`���t�W�>4��w��?7��Xs�T� cTM0
3j��[�S���{���"`hpJY����P��5�@EV�g�qƸ�@��٬V�s�/��Y����;0@4.��% ����vvv�JD�}bbb||�M<7o�H_�h�~,!>3{"~Z	�]��j�4�(V��\&D�8Q�Ћ#@6::��9�%#�g�y�RF�fO��y �Q�k�(�c|۶m4�El4�X�"*�E���3yeN�P��`5���'醁 �x[��G�":��	`��9�H)�0��P�\��UQ��@m�'c��+�֎J�VQ~�D��,�C���I�}�)X�#0C��p�B�K&N�H)�xZ� �b�����g����N���ʽ��;<2B��T*��_��M��b�Bs���̙3�=2�^�d���!��E����M4s����1␒������kK%��G\U���DyV��PD�b~���:=>���>$�"�KtRV�;�k��$�1.XF�`/f�T1�����S�J�o)��=��m�SC�����m&���TЕs�#�ڮ]� :G���ji��a2{��l"��C�d&Y��"�Q2�b}	�!�;o��>�ڹ��Tb�z�J�<R�݉��B�ˠ�.��М��������bA!X�Ĥ���/8�y$8dľ�<d�M^Ii��r)yd+����y��� SS�����"���IY��\75���X�	+�)�\��dcwMQF��8lIt�W����0@��V
HE�n��!��nHV�>bWJ{�U	�!�S��Cz���P�HIg���BtkbBec\y,�.F�H�#�><H/�=��������ig�}�t�D�~��������������X���X��T4�큿
������B������SNϓ[U[bD���<�V����B��7��`q"�F������瞻����'�$���Q�lٲf39�,ˬ��EK�J���|�6�~�衇��^r�u�]g�bϕX�&��f+��o�%@~�F�A�T�(�ldT��Mؕ;�-K�>������j��֭���t�
/�,-.�E5�>h�/~� �'�lC�B�5!�B�}��zه�o�aJ�N��T)1iuE͐��o������'�e�^�t�u�M�`QS�����~��1��5��@�#�%�c��f�ȋ�-�����~VN�5?��C��	'�pŕ��[5#�X�L�>k��>�����$ro��������s�|�;�b����YR�Q�rR#�(ZsiD���9����z�IW|��f�D�RH�l��6/Nn�����#'�|��W^q�4H�iI	/�f��d���j��s�mw|����7'^��KU9Bф��~�����7�<�;�.���~ܒe���sj����-�z���Q��2�� ���j2���u>�
��bLFR��b�3�Q��cr�9��(���hO�˓Z��%�D&i��)!H$'qmdl�����]P���3�"�L�v�m˦f}�J�nFM7��`���RW�XT�M��ʥ$���ޙ.������;z�}K���dp��;�WC&���jA4o�2��`sR��i�. ��,"���Bq�g��*�N-�H2m�TJ���4B��m*��I�Ϛ�hdv�6N������`rddg�A&���'B=�r��g0��F������X��CNִSY+P�@}b����3P�"X�
()���7D�8�KN������Q��*��S.���>��D������&hN_��*t,%ݴt#!�~�MxA���#"����4�D��"��4򋘽kJ��M�i�T�괒*=�%�Z��Db���X�G���^����h��	�u��z�z�Bqh�.��Bxk~o��B6���ز��9Rh{EMg�E����/I^H��RT�(QȀе�)g����	�?�Ɣ�`M�k��8��7��C%�Z�H�[�G�1Ex!�Q��XT�e?��*kd�Ϻ=��w�"�´�_M��3��ik��:D܈�P��kV�rc��#9�t�q��euX�<���vĜA��L|����@Ӛ��6J����`�ɤ	��jc}�4�Z�,$��G[@�d��J��7u��Y��)f��^���h��Z��� �EO�9{/�C�KJT:F�`Ed�2�����^!��G;5<��|�)�R�-n����H�*�F\�Ʉů"� *�I��~��˕.�i�KG�K#"c (�m[�Ǹ�)�H�#C�h��ju�"8��G�0}��r'n�:x!��-��}3D+Z��Z4�؁��� KA��U�x:��
F���NL5��z�R���G�Eߎ�d�-���h�t�jj�qU;�L^�^�8�{�F�5	J���.dS?��3f̰U<�m��-�lڲ-�;4���[w���,(-	�6]V��O����o;�LY�uW�`_>�K��I��M#8yK�E�=[(-</����W` ͛�EbPO?��W���g�q2�ɆP���?�,�� �~��,��������9���}��fC�<VȮ���<Z*v鴎<���s�w���

Ԙu+��;n���3O$hZ*V$��Q�'8I�X$���^�t�z���y�#� ��/�C��aY^�|�����DÖu�%���@��v���wԡ�����G���	;E�������~:Mǂ�x�d#:����C��s�\�R,�,d���[6lذj�*Z�����G�������ŋ��t*���{����;�3W]I�G�A�4�<"���IB+��~AhQ�#���s��z���M7�t��䒋����t�Q֜�P�VԊ���o����.���/�\��[Ґ�evC�P���������7�Y��?��O]���'�m"z�я~���.9����5Qj��XD�9?^-�R����p�(���X���x�D�<o�¥$��%�zVE�d��\�5��0iAʬf�Φ)D�U~���'�`ӦM��N�*�:FFF���~щ�=eFG�ꍾ���-�_骖�XJ'�����SOu͟�kP�]�v���ҕL֛CCC�c`����m�M�(�t��V�X��:��zNz؂�Ջ/n5uiŊ�4s��M9�L̊��o�[1��J���%�Y.*szu]za��1WU��N�����fqVʞ�a�n��943W�+�x�
/F�pD�C�yu�)��`�=Sf�.���2t.����y+֑�L{��<�ל�6����yE���RG�c52���!��$��a�.��$�/PdU������I�:�;ߡ'3�"�L���-o�6�if� ����m�Ī$C��ٟ�]�v�ͱ	�9蠃�̝I�W���֭[���X�p^OgT��ux�h ֥p��E�}٥N�i$T���p�["ʨ�-ok%t\ʹ���uJD.�6��$��9sR��:�`L��a����{_:��S��e�|*�י��KKc��9\�U���r}l,cէ,�f��h�PPu�#Ws��m���go�E�<!@'�\�����z��S��"ӛ�L��r��U���y�<�\��I�}�b	�;������=4�/:��?�b�w�<��1�ZO[ʪMҗ�`6@��3[$g9W����"��m���K�a��f�=Za�FX�[锦��0�S�Y�;��	�8�Z"~(5��$��qR*�
��Y�h脤0*Y�8����̲e�hG��7�N�h��۹�.IM����X������FMhӐ9ͺ�%HUQ�7}z7�p���sM�_|�0�>��� t��wO�i��_��F|���$�����/���KM�/0R/·�i��v�5���,K��׫{�"�-DK�TD�Z �\^�I(L��5R ����R�<��IoJ!R��iK��_����ԱE�$�cy?Қ5�=�����U�>���|͚5���x�ۉ�;A�v��KW����$�M���Do$�'D8.�%aʀ�tH�����,)��X�)��7y�Ω}\�U>°
��l��(&"��W�l��ϟ[o�<��u�ʁ��
��JZ
�p��'4cUP�j*Z$�5��*q����h�ݚ阴j\�t�����.*�W���3����?�я[y�d�b�n�������������P�PM+���������y�?}�����>�d%?�bS�,�&����7;��/�3-Z�&Ԕ$�6	S7	�Htg��q��/���n��?��NJ��F�*�,<Z�د��������]���3�FF!
�ӂF��x�a�z��R(���\������_��M�U��-�����/}�����5Р��r�`�w�>��s7�o��@N�"tc,S�d�kJ�X����l�T�Rx����22��~�����~����UCT*'iA��$�i)T�b$��\�����Jhۭ7d��hk��5]��� NҨ�	j�5}bS�ULRW�ʴ���TL�R�Qwy�Je�E��P�N��]��p�j��f��\��C�M�Qr�T�5�P��M���`,��%�Hl#
�+�R�W#IB@�+�Y��u�y
[�V�S��zi�	(_Q��2�=��P�㬔�1KJ{�n�*�n�K'Mx��en�v�˴�(U�c3��R#A����e/v�)�q�H9cM��Y$�%-����F{"��u�Z�I�¿�2����XV�O��.ۦV�ei��;a�<?��#`��
�\��Ao]��K2�5U\
�m�qwr�9����@��}���Y}4���.3.�US�egh� x؄�hն��4�붌�qY�j���$X�Y�ltDQ��j�.wԆ�}�́a�]���H�%n����P����2@TDA�FQ�TlY	�@S��b~����,�2�����uP�s��E��T�E�� ���-�H��/�,�o�R�5pJ�N�ޱH�ҚlIN�"���]��?�9���E�^��D�7&�����ޜ�� W1RK�R�4���:;+�=�!tV��6�b� ��Zd�7�ݷ<;�)�IZV�:Ȣ+r+w��E�3��cG��֯�d�	r%�rRN7�_i��$�e�7"s�@.F'~e���n���(�in�+K��s%w�%`�s'~�e)���j�zv3#0K��ʙĪf�&�*�b�E�t2�D��y�i����fΜ�Y�W�%\��&��kY�/D!+�BbJĵ@nU�5.��Dɢ0C�\,��J��$�httxbl9�t�"ѷ����w�ٴE���#�3P�b.��A�g��(�<͂E(�!�)ӖjGAԌ�$	LCO�Ԗ���J�qG�����;�Q��_(VW/[�]頽i˦퍱�e�ܔ��qhll��Y�<�0*�����,qET��
WN�TV��q�� �)��F��p�����;��e�E��}	��s/���?%i5C�}��1��irG�Dv�l��W	�4�8�,ϙ3g`�f��"p rzӆׄy��m���D�aG��@Xl�s�2*p��P�v�!A�5RI'0�#���8Aaj,C7�V |��ڻ�9��yt8=��En+��^k��<���bx#��o?�u������
	������5�}�3W�\����N�IIH�6OQ/�Idi�!r�|�g�}چ���z!-$��6- �H8*�@�T��_t�5��˿������Î9����Yi E�[7m�袋�#�>�Ӓ����}�߿��k�|��SNI[��H��t���Ν;��G}4�P9������n�I��������t��0�S�+�����֜p�	l
����(�u�E]��}�[N?����*r��ii�]ʢg�H�W>���^w�u��x��N?����s�&����)E	�TT�����`�6̀��������͖N��.r��=l':pZ�Pٔ�M�$���O�Pg=�@-���\/a����KjIC�� �+Zr4"j�|����O��3\�������hWN׮]Q���Nh7?���Zt���mt�ɺG��T�g�y�ȝ�T��.���N�Z�
�������l�����3���ӊ���8�جt�%�^.�N�Qq_Z���p��?�(��􏎎��=k.q�F�^�����}�9��Di:kl"��f�;���`YR�7owhj�_���d���MSm'�S�M�O"hY�-8@�,�Z��� !G~-���t��D�[.�ƴ��c��	w�`�"�K7NcT�AJ�r΂���C�\)�Wt�5�йTF��'S?����ڙӺ�����:���=X�R�$.{s�x����"���s޽r��_]��M�6��$TF�����22�$�6Eg?�r�&.Qb�+��B�����i^t��x2�n�8�V�%��YS�9�bɭ��'/��M�.�IퟕZ��<?�޶:�As�YP�w�a�x~�G�v�T>��O%3z�x)7����Eՠ��ؽ!���w��UV�,��K�"+Ҁ����X HB6PGf��!!G��Lߒ㉩@����YsV�Z����¡6� �Z���	/Bj4���ͣ��}��]�C�k�I(��"��o�ka�D���!˙�g�~x*p�:�������|FeD1��8�(%�y���ع}��믻nJ��7����^���&2�����?�(ْ��ӧǑ488�G�q��r���9�äo�vw-^���(yllb��B�v�kt��6;::?l����:�C�΀�l�t��O��Y����g��L+���T�"-__��O�.��&��U�[�z����rw>��vI[۶m[񺃎:���7�n���'ODnˎ]���Z�bq���O������)��S�vi�i�%�;^�Cn�9�3�/V�؅��(���VyA��*�ղ�iYD���	�B�.#sh+�I�V��*#a*1�E��Y"T�Q�e��a��Ҳ����4?��X�<�*�ԣ5'k��gmV�Rh�H
�I��Y�A_�7�"qڢ5B�5>��q�W��b()�Z7Y���-���3�%-4�L�.���ێ:������=��_ߏ�l%
���׭޲e0e�0�6~�

�P�"��{�]cX2��ck:k����:RP�&ǝ��CW���o�����7���'�|�ު�6C�Ɵ��S7�pC7���E}���W���7}�����M7�z�g���BO歪����w޵�~�ӟ��>���?�яw����o�3k6r�B�`�o�ͤtú��[�򅯯���3O?��=L���:\�(w����{�׾�ow�q��'��X
ɤ0� ���,Y�+�LEǡ���57�x���t���t�)j=�M#Z��\�x�߾��&i�(��`͏/����|�{�x��N�1��u/��g?�շ��c=�e2���n��� �w��P�{Ў�����І|�+B扑Js��˱%�Q�:\*�Z#x�%�4�8�ݏ��mϚ3ol��ޱ�r�<81L���bvٳ�����k��ɮ�!pRTK�ɺlA÷�����n�H������z������6��'h��j�@Z� ��P�V#E��$pȆ"LdYz�<��3
��N�s���T��Tm�J�zU�Q��Bܜ�YB.������I��k�]2�Iw�ߕI#D��-��T��\�)�.3�E����&Q�j�����"K�Uhx�٢ �&)���v�j&d���#S�v=a�yJ�@	^ǲ���B�m��r:UϓJț����M����U��*s6+d�(�8Ԉ��j�0mU�L�����F��Ę�)���XTI�T�E�$Ց�(��&��;q�$	c�:��:Ni�\��z�6Ѳ&ϝ;�R�>�]ot�Xd�I�冧�VT��A��sF'��M"|�**���"�.�q*5�eY1�4����I�Ѵ��M�,w�.�ߩ ��9�h4�>����Ѱ4�yh��Y�I�	�ǔu����2Y����gD�
��pJ!{����'�|�;Ճ�)��J2_��d���~��Q8��sA!6�[�"\�T�,43-͝5 @-�J����(�N�L�腶C�1���4<S7;;܎�����r������;w�E�'&�A䗸��x��KQ�����E[�m�#���D�vJ�3�D���T j>���2}�]#�f�P��Y�4���h�S�\��)a 9Y�~�L�)���g�D���7�����E�o�{����Tթ�*
� AD�	���h�)�h��&��ǻ��ާט�zM�/1�1�IL4�T��D��
�����oV�֛�Z��sN�`PRߐr���^���o�f�pg�i�f�����B���M�V�|�$+Y^��8�����G�!:E˫@�ܻ��*�rP1g�$�0�4$d[F�&�d�Ѽ�XD��9THWʭ��؊҃�{����X2�s��U$3�s0[� K)��0H����R�-�Q���UX�s���d��S��SSSv��%F!B�^w�R@�IT+kU�Z��-�5ߋ6Ol�3�|�?��q��\x^�=y��������^ץ���D?�^|J�&|�F]R��6Z������m�[7�ח��U+��:�1������c[��F�}�q�]Q�jA�� 4�J��hI04=��T��P�6�& �V$s�ق��[$bHp��W.����%en�c諑�QJ涒9�>?NK�Ğ`�=�P�F4�{�%S�9T��d�A��U�00�16I�qVa�-��Tg06�3���4���lc�V�b"��H��j��mA�bƻ�`�D��:J�)�;b��V$�
��+���Z/sÊm�);���~��A�y���<H�_|��~��+�ٿ�����8JV�Q`\A�??��_��_B�RIV"f�s)���<$#7l�c�2/������+���W�B5�Ȱ!һ���?��w���X��~����w��]��rK��b� �u�ر���G?�ѿ��[?�?����f Dȳ�����
����3ӛ7l��{
�z�o��o���=�k��ĴB��48019�|�ěo�9�p�H��X.8������w���&�����<?<9��rq%s�.U70�V��̀#b�}�7B���"6X�z�eZ�A~~v����6�8�$����<T�&/��iHГ	i0y�Jn�e{<߅�57n�����a��v��Rqll,j��9�>1#b�H�5hգc����F�a�H<>R�t:�Dwǽ��Ϥ�u��Ĩ�j�`����Y� ���:�"]��ڝ�D�C�2�n�ŗU��CAw��L(��<��ߢ��
�vN��?~�xB	��b!'�J�U�{lF�K�4ZLd�G���@ؖ�鳥���*���pLad���z/�9i�R�,�ٓ�b�ET�'�`��9ד���R�;.�ҍ��i��iiZ��J>\�=����+�|q�i�����c�ȇ��e`����l�il-c�Q'po���j��r��Q�!L.��,��T�_drrrlǖ뮻�A��A��n�Z�KL/�Ęa���Ɵ���h�7�>�C��N�0AomD��GV��dn�ݜUE��oC����7Ɉ���?pˇ2��:�0X�2����h��7l؀����76s���<�2Q��X6���FUQ�u�REpGXt����������T)������.�cW`$k�4 	#UC{s]H�5��A�J7`|���ѣG������QI����Eƞ�^�0��y�S7`��9�9��!�$��>�3����pq�D�|�6�����òQi�*2��K��-�<lR�c��9���z��8 �����Ʊ"�>�rC���s�x>S�@�p���R�l���w|�=��/GVÊ�H
�	������'A��p��]�駟�L��׿��K/�_����cbb��;��2F�+�![=U�������wA^��h�噙�|�o������0�N�<y�E��o�Ma�O�Oa��O��gSB�Lx�d��k��k�����w�ݵx5�X�6׌N�g\�l����/���""]�,��ս*��Wh~��F����\%$V����3�6��a����Ti����ߟ�����g��V�������j��_~y8 +���:�% �X���_�������d���,I��X 8��%��PD���^8�pZZ�Qj{����[�������t������D\���ر�T!a���k&(��7P�<�����/�#���;n~�_��g;����
�b�����E�J$#�{����5�+�>����<Ro�-�T#�]�2�'^�O���G����wDּ����֘q�Q9��x�0��m5�44�1	�X�t��{��[��,z�\�"F�GL���6�ʔ��1j��"L
H�S���p�\+���uD�WE<���|�����:�|cq||��m��,���!�e��NTd�
�n��Vs��"�����$��1���=GK�R�o�wA�Vj��X:�ynވ��V:�y/vʤ:<�䓁����c�N��a
v�6��sLn��]SE�����j�Y��u�5�'O�bL�g-�s!r�(�
 h��DZ��h
'�:a�f��J��o�����uxH��e.��RP�L̢��&.X�����ݲm+�B�4�E����|��S���UוTe�������l\�*czM(�0��kb���B��z�*>)<!��Mxf��2#&�x�04arReg�1��0]�1q����(	�c��HU�����_{ru����F�~��_p�?�3o)�侻���ln��
��}�����(ٷ��
׼�����w���Zz��6���v�A;0������J�~��Z�Mѐ�jy��42aa⏆��K�~/��+�Z���
I�(طg�IZ�L�#+"w)ۣ�� �1a���`�J�Aɐf�RH����-%H#R5�'R������0J�R#1`}M�{@)��?�#3���D�r���{�KK'�֩�Y@�1t� ��m����/���X�U��*���jz����n�}�n���]�}+�4#^j6�f����Zh\wݵ�v��;��g���i�����v����3O?�j!�w�]�^�jI;ccc�n+��*�g7���
L@
{�ƽDY��!����X�Ͻ�Ɠ�d�ұx,�ߘ�>�T>�$�h�ܒPI"L����R%?rL���NC���)�>�/��y�J��W� `�B7#�F�����V<@vm�?����19��u}i�.4�#m.R�@���ƈ�*߰<�у� ��K%��#Ī���� �������<� �~�W֒Zɚ�E��;a�~�����?�_E�w����˷6o߱iӦ���݀�����4`�n=�w�L���Psؘ��6̜m[f_��k�|b������t���nvax�'w���?��O?3�odԾ�w:t뵸���b�jZ^��۽�e����;*�2�$0�?��J�+8�����҆Q�:�t%Y��̌8w�.CrZ0�k.:1a�*湬T�R�2�����Z����U��"T��[�3��̎�A**3/�ۈU���;��a���Њ8�Y�`F}�C��?�����c�%/����#���]vo���c�7�G�9^��F�-��������d��:���.�����y;e�A�~�����T������h���N���^�� ��+n�. C�u�F�)�q0X�`\������h����������Z=��{�/�������7��K0,ET�S7M|*�˥�^�{><y��
��K
k�"a�#��>��/�»�y<׽�꫙��J��\T�q�'dX�0������=����5� z>�R����7���K.��St<�h�W�R��eVy��R�+�(�?SC���2��ژ�~�ԩ����YZ�+<v�\.�6N��4��
�R0tD��v�(}�$�Q�փ�>��Cp���x��ރ�;f�=W*����
P��Π�E{P��N�9���*C\������L%L0�g����pGHLLG"��M��4�[B��P/�HB�%,���y4���t:�"H"O��Y:��4��UI.�8*E�("����W9�]]������"��cP�܌5v��2���,�l�E�Y����6�p�p8�Z,�4��O�{u�\}b��X(O�Rb:����*I�ճ�>���cq��Y��o~~ު���"�?�--..6���]wݕl���ꫧ��p�����0w��l9���>7 ���{!�p����pd�,&[ O�^����mUNOOפƅ�0��~9v�<I�w��})�G�Bb�>��[�ą�C��Y��ę�H�m�;��Br+-,,A�>��#{�왚���e
u�Z`��?�t'���f#����FL�K�
#8X!'�Q�Q�����bq���0���p��;w^��g����ӏ}K2���Q."@XvFq޼Iə�D}N��Şv\�j�?�s��<N�a�5;��(�x�'=3Y���
'E�ϔ�Z�1�'��r2 @��̇��Pe�tr*��v��:U8PB�TL������T9�i��S9O�$t��:��lj۷o�3)�ͤ,Y|�r�FyB�yj ���-�7MMMMό;v@8�d˖��Lᚰ��:���\���e7%��y�a�>|s�(-��2������w�[���)���Ʌ3g�[x�3���������,,m�Я_Y�ڏ�����^��	cVY�j�>.8�j�i==m�f�r��m蛳�Vr8rq�E�CL�sX��bLu�M���_�կ�� �FGGy��"�(��%
 hie��f���Κe@$�h�9B,�u��x��M�'*S`�	��BݼI�n�Y�	K�N�#G� Qn0�,H`ߏ5��y�D��j�
9��}υ�A'fg�Ŀ�����qI�tJ�K�� ����.�)&}�cf"�/���z�Q. 3���~����j5�"�!��v�������!�]`[�\�	B���UbZ�#��[��w��5@qַI�.�#��/�� 1Q:&�ivA���MuH5��s=�E�0�
�z�sݰ�]��߱����IT�)n��A]��P���k#J(H���4
ݫ��||Ϯ�[��>~�2SIz��k�p��ȍ�����*���Tq��K�=o�M��"�p��ν��9��{[G&�l�ҙ;�����ajdSmۊѕ��G��S�A���(r��AaN(B�$%2t����ǝ {^SR�$��M~*�A��li*F	!�\�Q"֟T�xe���O�z�a��R�.z�j����$�1t_$a� w�̙3pӚi�)<
���\�^r@�����%���U;P���� 
]5�1/RR�X�b�W*��z�B��qz=^q�0�G��U}Ǉ�@�Q����}�Lfi̀^���'�vJ�
bKŀK=��D���� ��F�ONW&K��:L�`�O�M�Ѓ���Tu"^J�c�����}�7́�m۶��*`��!�Sel�*{�%��z������ &o:�'#5�!.J�Ɔ������Y]�J7�X�ʃ884��0���1TISN3et]��bIQ�Jl&Rދd(�lh~�ݖ���5�/󯰟T�x�tr�b�)x�,M�VdG)��UG����? �:t���w�A�;>�}􉠅�6%��v"�UV��T�[�皀�|����馛�"�z[��:ڍ�Ab_s�O����:rY��^|Qi�����{��������M��fL�:�� � �L&�i�!fukj��F1��2_XX(��Lq����	����=c�QDnw���6����F�+b�ҳ�ⰶ�Ɋ��(+�Lf�bA�n�0�X�����R�m��2�W��E��9��W�U]��R���H��S�l/B�Z�2G'���������n�MG!FS�Pt�Ay'c��Q�W��g��㵪!1J�*��vy�������`�9� �Pz�,�v�g�KE/��`j��1�߾�~������ϜX8�T� 4�%i>����G����<�z�=fs��v��!�ݾK.>x�P��ݿ��<�w�0��Π����Z��_ܺy����X�n��9��L�RQf��H��Hj���B�y���h��٪������@&g�?>oͺs�n�:���"����f���dס+++��1[S��T)2�S"c��H�?9��n19��,KBd�V�s�f3���9ke��"��"��sX�en��,԰A\�|���?����O��O>�я���/I*5�()R�t��qV��AS�;E����3�-ɗ�B2��3�0}fJn�:k���:���`���*S��يŊ��|CϛJ��Tńk[�E�El�w�uן�韪�&)���k�DEX���뀦��������2b�$|+*�)��~���{eS�t�Xr�'D���쀪�x�<��j�*[@������O~�mo{��_LV=�����TZ�ϣ[x`��bt������H���<�x� 8���5�po�I23K���fW�O�I8��� ��l
r�T*.nz�^>�5+��-(g###l��V�$~299y�E����?�Q�u��<��� d�9�?�|L?gFt#�(2WN�̦e�Ї2zW��Jf]�7��3�]syPʓ�xu��c5�܊E��4ыs�ʆ&�B؇Ͷ�#+Ɉ�X9���Q���"���Y[�灡���K��N'� ޛ�(����H3ʽ�4F�/3*Y�z�����0��^�<xpr����x�6r~�8;���o6A{��}n
C<�cF���4:��
v,0n�Z�kih^��\g~~�q
�`Q�B�G�)��m��!Ď���HCm-9�/�� _�:ܱ�b�fR��F��,����#륶�W<[U4�f+�{�?+)��'*Ӗ%h�9r�t��3$�
�/j�f�Xg	$:.2� ��H
k��b�=���j�ةS�vJ��� Cs������Vi�Mx��� 0v���'�MZ��/���0"��Id@��Ȭ���i���Z��&�z�Y{���ʡ�.9�L�{~;�k�+u�x��2�O���vץ�8"�����0��"���9�\���x�3-F懄��LW��U(b�+*)��O�����H����q|�d���.X� qAr`�_ 8y�c���ߩI�_9q�E�v`���G`��X{M#��k�%C*���mKKK �A�y����Z�A1�f�;t����IxrL���u�뭌��1,~�^Mu�������l�z��J����'绹8�,�s��%�4-�!GXz�H��p։�,�r�u֜C��C_����w��z��"5�(�}�T����>��o��C�l~��17I��qFB͑]��R�
?c�:�2d���tS<�}�~'���!l�\�������7���!=��d�#����!�(*����+=�_���0r��0b

1�b�̃K�Ґ�.B <L`� ���Qʈ���|�`��Fi�'ԁ��,��ȌF,����P��F���Ja�Su?��Æ�����ܙ�o~��g��T�`fu{Z�f�BO���u0_KU͒��p+�~��QM?�W�@K�d3-�E^]8hJ�s��۰U}�V]M�S�UC.���;��*����n(�N��Wo�
��[��f�Ա�����%]wzhVta�q�+���G���H��k���>��<ߌ���f�AG�lC�y�!�T�I�<NRF�ڜK$�d��(�*�t�-t5l���8��
���XTQmtQRt�7��0$5��hE�V)��P��	�l f�T���i��ۣ�%�д̾��
�hmd��=�}��H.�P��d�.��exy$Y\;+a|�4p���*1��9Ԝ�q�+@<���X�K��Θ��t�n�W� eI{��8���15N1�����M�e�a\��:*d���z�X��g^h�B���������3����u�{{��fͨ5$�#�V�S*G�M�?�-���L
ʧ>��Z��7y�(��x\��潦�j��%�ۖ����j�4U�ŧ�~�v�6沄�����l[wY�}�R��T���<�Ϫ`��=
ZD	��p���,�u	�����$�g%����3W���{�B҈0+&��z��hϴ��K#������j���#O=6��D��S+�Z2��+dA�}Y���3f�*�9�B��<��3�Y�l޼��Tmfk�u̲9:2�Yh.9s�얥��<���}��}�Ʈ�{ێ�&&�p�Ex���"+H� �z�Ņ9Π�Ç��Q�OSW}w�"��B��z��n�e�e�:FCQV)��}E�S���,-��|���m�C����8Դ��0�T��j��*��X(d�S6���c���am;���d�ĺ ���EJ�2�fK\��C8
n�1�zr��%֧��]������]_#�f臖i�
F}�ѺG;�l����vk�@Ih$�'D�����j��hbl��g��?8t���M����7n�^l���5 �ܤ��xqI�-y��-��;�����̖�ۧ&gB�������(�m˴c���>1�K���N�?7MmYdh����{��F�VTm������fd��m�u�U N��	[��	�v��I���`w�#���8r����;�mU�g���\��2ϻlW3E��C���j:��!R�4j*��ZZ�FB?`��WS8�@��?���$9m����xG���.^)��z��I	dLJk�\q����5Ej�P����g��΃.R#e�a�{�ĺ��$��d�ZyyS�tIf͊��R*d¦ИX�9�"d;P�E�8������WZ��l�zJ�80#\
�lA@H�<�\@��Aq,dNn!D
��D�-�8�����^�X�W�̜���IbQ�iJ5�Z͊N��5�W@��r�-�~���ڰi:�O�q"˹������,��'��%<��<6�X#���A��B:鬑@�7
`�VHo�� �0(c����9�$a.MMM��G�$_*�FFF\�����p�(w5L������?�8�6m�:�	�Ih�Ŝz�h��D0�,�)���a3�EjeN�,ֲB��_�x�{��3�2�
�-�1�"�/�ƾ�J^��hm>��\p��n�ӌ��J�r�Ur����.��/D�.N6�8o��1Y���܍X+�m"ɹ�OgXf>��<iD���R};8<3a����[t��X��J����?�������P\�{���m��E�~��*�u:O=�|��f^����ڶ533S4�,��oܸ1�Jn�:�i�����ڋ�c���޽{K�����`T�m�#U�䧅��n�L��)GT��E��3^�X��j��Q�v+����x�K�%tU�j:�숈�g��I5,�^�vV%��E�'C�M,;N�
[5�B�v�B�ӈ�sXB�bʆ�r��naA����0�4�b�W2t)L�:%�ʇe�(练�:��åM�(�E�]�o*�5MIs r�q���0]$8�'gN�����1��D�m���~�JV�a�2|�5scM#���W6���a�K�.�N�Yy�
&����h�j���s�9W9SK'�I���D蹍�����*��bk{�cJ|e{���-������5cL`J�<h@�(��K�N�01�۔��m��9fų��`� ����:�bJUl����gVH��ldI�p�9���=я������1:�~\m͂��k�a�o�9�.�~pW��`VY��y��5WIV��������ڑ_�(��9���!��d %�JS�>��&G_�g��֫����Z"���da�ZjiXٺ��M�N~$ɗ�?�k��hh��2�e�\=l��+�:l���$�[����V�$Yc-5��f���@�?����^�CV�Ǡ߉� ���UI݀HK8SCp! Pm�������7�<��(�»�Q,��G�~�+!�����*,n�Q���s� %����M:�Dv�����'NX��Q���b%��\�;s��Ѹ�:�Kg:߼��={��l���ѧ5�,�ݠ���;j!9px�׿�Uгw�����ǏV���3�=����6L�H�����b匔#�����8��4(IA�`�����n�:fK�
R_ĉ�IY�eh	��0N3��+�́�B��?����Ԕ�x�$��S��m"y:�m�x�*)�Bniw��XL*��)H�6
�'NcԜ�{�kb9X����)R�#Kd��V����	3��$U	�
��A��gx��n0��uY-����:^�5���!�2ҡ!>�6h���k>��k�����9�S(��=��.�!�#��4UV��b���� u����X�.b��j�����Xf��,ݘ*ժ1ִ�C��%V�F�������#��>�l<S�b��c����So���ӧO��R���q\p9&n�ݾ���tU3h�
�Rv��m'��Y~����m��E��w��=ـa<j�T|$��"剌X�_-�df�F;Ú�KU��t�T�j@��*�b��U((&��-�+ !��E���:H�+H9*4��?���w�0��Ft}�D���(�`@������a�j��F�eRYX��1�ePo��ͥ�V?�ԙk�}@�L��p�O��cӫv�o����s����������덀�/�p���b����su$> ����E�TA;/�����!7�84u51� �j�Z"�[���T������E�V�'%Cn�j�c�v��5��nD�!Z�,ʓ�[
- ��KH��X�JS#7��H�o�Ō"u�=���uG1�dx�$z#~�v��}#*�
�$�6�^rz)�va/JH�㓇0=U���B����k�Cd;K��7�g)��<���b��_n7���Da���S=
�v;v��Y0۝�:'�g��6�F�	�JT�ra�.�H�C�n��G��'Zu�Z/�ܽ���g�ĀU_�m�u��ˢJ�2�J�t�lۼ�1Q�h��CR+:�B�m�T�-r`�����q��!��5���~B��97�ÚE��!��8�a=wM�B�욵@�P  ��IDATj�<���2�$3��&B�#p6K�(����!���*�&Wv��5��P��j��� ���D	Q頱�TX�����#L 1��)���>�I��-`�OqOw�4{��U�R�'�}���T��0�����l�֏�%��(�W���E�˾T���xt$O�?�ƞ=A�9�
jZ�G.�AfCEQf�G]�=��f�=��&���&��e�/c��`�_ZZ����ַ�ռ�N�����k_�a���?��O��'�@ǎ�w:�Mc��uŰ}����;99����O�<9f0jղ�ƌ�2-{�Vs��>�;���lg�S��
�{�P�Fi=18"5DGS�P�%έ�""VA���bV�:�H��v_�P⻇�&���Yh6&R����͆=0�K�v�M�lT�*A����@�bH���Jh짂�Q�Q�dba�;��2-��9i@)�<(�'X�U�T���a���;���'���|b<I�C�V��s�!�z��𲾂�����+{�1�Kq�3�1rɍ�����@ϊ��ژ�SV�y3�AOΟ9#[]X`Ƕm�������+%Do�[���3�s�-#�4�XS�s�T�6r��n8L	Ouz�"�����Ʊ�!�Sf2���8���'"���*^�
�W,g�t>@2�����a��ã����z=�z%"AXG�>��P|a4;���|�{�f��鵫�*�"
��8����^�T:�8�a��Cp_�z�����������;v��x��S��x�	8g�Νp�G����k�/�B�<Ƚ�i�:8W��=����j>ɇ1UN":<���KWe��[�R�Lɜ�)�[�,i�Y0��߲���4��/��d�ɡ�R^�d�#	��$����#�� P��+��.��*_�y�<�7J�^���"I$N�����㎹��M�6%4o5�����N�t1ĀJdc%Ja�4��i�̐	�C����t�9�6�fH�Z�6d0�=>>�NÅ�àְ���� �m޼F���n���c��)i:��w�	����J2�nB���Ȓ�[�9A�	���lI���<~��2[չ��h�M�_��h
�<�0��ڪ�PH>"�R�2whsG�`	�	��{�Z-��(��U�B��&-��Vu,)�H�(��f��b��(�5���)JM���k*�G����xpk��g�{e�sX�eo�ɪD�Ս��?B���M���W=�u�)���=oc�����{���eAl�IZ�%��Ww%+���uȨ#8�$�CTqG��/���r!��bt|�t�9д�U�
�&���+��xC��P�=�LI��V
�R"��P��,��ر؆i����:�ŲnD��p�9�G�ؾ4��Eo���3��WTS��0�cs'O.��6��� B�T*��B��n-�OI���,� h��]�,U�E�S~E6N4v$(AFþ�I����|GkY�\xl��K�zg�KX>N��q8��gH	�h��.�CW%�k�:�㹬��g�"5T�Ҩ�$t��������D9�;%�C���á����HfL�.Ȋ�e[�3�q�qat|��������Z����K��:N��`[OW� �Q_@��XqM�/�)�<ᵻ��h��A�����~�M��l͝�k����"u�0�=�8(g��t��C�%�ѧN��$1�m�T=o�v���/�Ԫ#H-���/4}��UA�ޤ5~��W��cJL�_|j��G�w���㏜�ҝ'N�!�����������n�J/F^�z���l]��(�.����j5�A`�B������y�#Z�!����zJ+��f�4�_�<��1��d8$��ng\G�s�Ez>�_�sOJ!�Z��$��oֈ/@�~T�ʁ�N�>�_;~�D���O������O�R�*u�F��	N`u��R{�V�b�ɮr��i������t�ǻ�[�oW/�u�^��0����q�c]u�n~�[_����7�|hia���_k�{��U����"A�@�{ku]-����F0���GA
�dZ"I%g�L�8Zә�B^�d-�
ʞ�zn+�ə�Jd��Ղ�{A �`��]X��qTv�"O��Rs0�;�F�~+�0�U��{E�9�m=x1� ��>�t�B�9���h2��D"�3��UAUU(�]�$�*�����0�A�lԛhA���[k�aa-r�S�4>*&<�[�&�b���b��*�I���{/u��h,�(����.�ٵ{�o������h�h��[�'E�j\U~⧯�e�X�^4��-�ʰ��ݞ���%m��\?]*$w���_z��O������BU-��v���1���12=3��w�5��_>|�����%a޺I���>L}�0�}b�d��Vʗe̎CG�Ld���:�^�F��� 	!7�3L�����A�Ly���uR�4[4@D�&��|>z��W^�l�z�čy�@���>X@us����_��^C�G�Rf��p��~��(�M]�`�	2����߱c�پ��/���nw�\4U(�T	#��Z1ձ�����?�{7�x�
���ށ:�4_a3���Q7��U9����6���טy���|���g}_��h�����P�f\�M�&d�BY[^]d}>��t�Oq/,LU�M���qn�3�;v����vn�t��]��[�kP
Nh�[��D�;	P���������kw�m.2�T*��E�$h�p�0&L�z�q�P�Jud��m4O=�t�߇�ڵk�E���������:u
p�i��6��i�`�}���5e)�"��
�ys��RyU�İ�c8�l��Z)g�0��Iـ���Nöy�
��0^y~eVI���]}JNoCs��ɂ�4v��5��L���W(�i����"�.F9�9�^ ��Mb/]E�:��i�°���S���}��
��az�0�-3"�3�|��,�Ԡ�A�	�5pڙ��|^X@�S��mH-��'���[��Gbr���6�yq�V}�~5sC��)�y��\�Y��թ4:;_�2��/�R��� �������Gy·e�E����SÈ85ںu�c�/�8�l6ӘҘ�a�"
�[�; AGGk"1�];�x�疎��М��냖�}�-�D����g���/��@����� ��59;�\���I�[�`�����%���y�q.��I3܈\�sk����u �W�T4���XIӥ�Ӓ�*�D��&�acOu���E�f,�5�f�X34��95�D�".�4؉�_V�;K��S)��V�H��)�Yү�'���B��dK� n��/`}�v	Ɨ�dkU��0^��1��'VC�T�)��:^���t��/����?9>+��I	PN��+.���M㳷�~{ߏ+ekl�����={�lߵVt��|�;ߙ���M,���CN��A.\����<����~���u�]���D�T2-K{ի^��5�5+�c����C�UA�6�3��G�\D�b��V���mn�sp�G҆"?���X𲉐��0�NLFE$�Eg8�S�
��~�7~�ӟ�4EX�~�߼q���o}�#C�Fg�Zp2*�oz�@|�+_�;˅��8�'���8�s�����}?��'>��:���iF4�>E�f��|L��vh/�~X���Y��+���a�J[#������o�{�^���o��d�JD��俢"Gލ���<E���u�H�?�{�^l3I6����Cn�B/LB�G��&���qQ��Dc�V،Ӹ�$/��Ș���2������(�A� R�h`����FM��D(��ɃG�F���l� *�ˣ�Q��D�CPޑ'��+:�Q5|B���-�ԥF���PdZ�&%J�W�H��DjtN���<��G��@)��	+�z�^�߬ק�'6LM�eDw����ح^�x3Qtdb �����|f�
��e֓������4I�)!�J)hxA��w8�	9�z�Y��4&*���C�tUJ��q�<��G\��A������3��؇[V\Ԛ�5�����;Q�4�x�<�Pb� pƎ:��"rw��N8h=��E��fuM�����z�m�V  ��2�9|��Z����
b@�_Z�DN�0�ʅ͓#������׷NML"�B�9sf���eq��h�7	j.u�l�\aIU�F/ٲ��� ����0�]����l�A�\5.��E5a{��y�3�F��i%�t���a��4����q6��C���U���@+yG��4\�$$�֤�u/��2��|�<1�m/��J��s�k<(#��'�t#I���7�������e�[�,И+����EO=����%���H���S�"7~,x�8������'�pf�_�>���b�O?=:?}n\�w���St��Y��4N���8Ң�ׄӛ�X`7<a��W�r'Y����@4��5G�4d�M�epu`^D5EC �l1��a�;x�؏S�B)jC��u���ʺ����^��vTѯ/鮣�9�E*ȝ�^J�2���,d�$ac��Dʀ��+��sf��$�v%�#�X0j:1@E�p���=K��̌
�|n�*�D�G�"�`�z�E݄�9
`��`u� �|K��	+.Q}�T�	����"����g�l��lx��s�����x���7���a��7o�Y\�C�n�W^y���@���{!��o|�KO<y�\�ui,,�\t$�4t�B+ ,T�t�����y�h�~�-?���:��}�Е�.�h��7���Z����c�u�V�'X~�l�� l9d4݈U�\S��X�Y$�� %N֦��_~��L����]�S�U&���'��_��SrxjˡU(_a�JM]"�M��,@;��w�g��Ӱ,��ۯ~�������5?��?��?��oٷo��#�l�������Y]ыh\�a���_��/�y�>��y��8�mU�|�RT�=����?����u;=ӰTΌW�"�1]����o���fj�v�_�Q>'1�`�ryX�a�Q�7����⥶a����$e��A.>������(#�X�J�t#:{�4��~�D���,V���dY=t�,���!_fi�����G�5Tߌ�-�=b�KI���,a	Զ;�ܫ���;sK��A���R�|$
��z�-[8	�9����~��U�z�d���N��e&�X�+�N��%���\��E���ٳ����t`ÀG����y�:f�LN�.r�y�=��3�zc||� ���%N?�\3J��H���+�IR�Y��D���:�b8)�>#�l�q��a:�0���4���;�uC�-�OB+Y����<��^6�Fq31��4\|�ATTR�Z�����W###�b8�(Sk��{���G�u��t(i��ju|S�\�@��L+��<yz~t�:�sǦM���[���1�a kA߂r?555k [�K GY��gϧ,�qj�;|�8�鑻Kui����Rӹۉɓ�=6~ӿ�Y�.r�������^�\���_]��ڰ�K������ט������*lG�Mm�ƍ-/|�O��b�V�U��Ky�ЉDL�&��Wk��%�#�/v���0�fzzz��s� �>q�i�':YI�?�|���<^���Tnyna	�j��?��"�,��f�Tpe�I�����ȳu
�����$�W�		����qB2X� 8�����z�@J����QR�}�QK����QL\)��$��Xx(�:�KObx5��c��p�2B�(�ś�b�GJq�!e�b%�L�st�H��Ϫ�¼�7��G�9s��v�P���gn+�7�mXA}J͍M�g`�Y�,��8.��60�����Ӳ	�9t� �o���׾��o��a=�>����`bb�UB��(���z� $�-�ufatÆ>�M�Cy㊲Z�@ C� ���5WC�֛�M%cd��z�h��׿�裏9tfll�Ҋ�*d1M����U{����ej+��P�5����<�s�҆#�{��B�⌞�=Wy�"ә��t%����7e��p���ǎs��o����.�,iߌ��O�������W���+.�B8~��k(F��-f0������������/��7�|3<�	˖�᳟�,��_��_������9���.>��#�]�x����������E�wT��_�3��z�ۋtj��ڰ^���b-U�p�k��÷�+G�<��S>1����1Y�q8b�,g�4�[�E�`	��,�T���$w
��d��t������8 ���͓���5�P ��&7�2�i�1m���)"!��
\ YY-��-LK�ò��ㄎP���$m��l�"���sZ�1N� T
6�\�Xl#���u�D%ū�H���w(�5�{�i4�z㓓�����~wi�O�f�8����N�5�q�A�]��	�Zb@�����lc�c��K�D͊+����a0+���1�7����H�e�1��Ұ�����2D�
?�*m����C��#"P��E��;-͊Y��p�;��읚v,��)a���B��" /h�U�'k���`��
V�חE�\�LT7��o³͎�j�6���AR�����#�Ҹ��7�+uff:��ѧ`�L˓�v `�Ges�4�S"<�$,�|!��"U��P/�P��5�U���q#�K�:�q���:�a}�F �+����V�\1�3S|i(ޕ�u�r3d�TR�(G�^�L������TA�ʪF~Bk��$E�c�p�����5��C<�i��%<�S֑��/~0C؋Q5M���w~�a��ǻ�kwm�S��Dщ���ыH�G�n��z���η�Qht����?}3�@�SԢ�^X�}��]#.oSj�la_�0����h�呂7_���i�ە��0�-���rReZ�7AiN���[��� Z^��f==k����o��&烹X��0C�1f����1KP��}�BŎR�R�%e���~$��]�D��Q���Ɨ��o��7��[T��0�g"!�}2A9
�H������! �r��
h�PУ����w-����Y��V�B�j?���X�{|����4Vȴ�h�Qg�����c���35�\!��$V� 1T�sC-��'� t�;m��]�{��u!�ѧo��/��ׯ��u7�x��{0.�4�b���_��g�}v����Bv���I��-OMM�Rc�Q*��x�E�����o���篺ꪭ�6n�j-/:��03s���{�u��Ç���Cp߱ѩN�S� kA�R.����[v]|��$`�$Ri��jJ��G�\�Q!߇�\�׷�E:<��Uf���slN��n!������T�2� .(�x���
�������i�Մ	_,���������H��{�k��P��]�������+������/��fd[�1��o��3��{>����Om����~�M?q�@�th�:�h>����w�?�s~0p��3i�:T���7��a�z��,��WX�^�ev��@�R�^2|]c29[
Ջ|��O��YS�@�{H�L�B2^����g�.��T�dk4� AW@>��-�2|X�
�h���l�j�_i���q�33w�&��j��w1>�qf]ł�;C&��+����ʊ�đ�	7��V2vo��� �;���ӷ�
�z�Tm�.U��"2;�d��u�vD���c�|2�X�:ǌ�F\Ԍ�T~`]}�8ccc�@�C�}�G�����D�%�e[���-V1���Ĝ��C �I�`�m�ai�U��ˆgA�XU��Ł�H�#5�4���}�[%���p�5*y����jc"U��|���n�8=)\�,�(�/ $��`�?���P^i��7\QPM�c��li�3###�OS��U$J�ڤ��̫(����Z�V%ِ�,�b����֢!䚓�*��?��qΌ��D�^��F4FD�j����3������B�";�"���N�ߚ� ��Гӣcн"�?�TG������
�z��r�Yr���͛[ČL��T����F��`?��7�H"��ӹ��h��tw耲~Ɉ�OŽZГc�6��cii�G��>�\��d��H��lt�('ɳ��� �(O$LGt]�e&bI&-�
��e�^͂��1�e��]%�O�P��{���%�t�ic�+f�$+8�K�OI�"�����PmzA���k�&�
:)ׂ�o8���@o���\I��p��"�t��|�����vmCv���?~�ĉ4��^��CÄ1ϳHL������x��:Fvʧ�z
`��������T�O�<yzqd)��z� *p\,#-�O���pB��ϯY&�ڏ��k�7>����]��/[fq�g�	�os�K+{"�qnٲ����}/���w���B$k��I()��i�pUf�	�I�0p�׼�5�y������q4�8������?�AX�7�t��SG�9�v�6�ȥ����oǪu�xף���ܬ�(�96����%N����q1������a��jz/|ˡy�=�/k���Y}�|���XCw�������x%
�엍0�#u�ȄJ܆z��7!�DUt%RC��˼(X
%|��"ٴ�	��$5$j�i���D�,T������]��8��|@��P-vM+)w�O�B�VW�JvE5p��AI�vw�E�YT4S�DV��������I]/���35�ؼ,�)F1�aW�Y�������(�D2.���8	5Cjj!�1(����.���I��(I8��$���֍�1|O?��m۶��Ltui����ۮؖK�1�pp $D�����>枆�3%��TR�������疊�2�( �9U+��wR�Y�RT���h��6�����J�~v��w�H�hFN��衒�)���R7��f��U-<9�Q�!���ʊ�{���*�܋C���1:���dNP&�nO��.�:�b<��D�[���Vaɲq˭�123���>	�z}�*%۞�1BL)ڑbY�*�7Z0�&�YB��m ���l �(P��^p�:�z�\Fͻ��-r���D�<G�dL$��R�@���� �k���,�a���A�,o��<"���!�3�P�a�D���� Y�Ĉ�0v�/�,�$���!.0\��P=���q���q�W�\�tJ�4��3��t&4�y���1�n�O6t�y�߈��F�s��C�}�4ǋ�F˒�e���Y�����~�a�!&7y�YZ.��\�m�q�Z�J��^�k��JuzΒ���IT���̹1�J�-���H���89�06D�> ��T����#3�п�s#���ⓔ��t�X qu���;X������G�"m�*醘E+c4d�V�r�G6���f�<�)K��_��Oa�$�~�LQ����,�Bx}/� -�X8̝��n������bzrOHM�*�����g4��Y��~�/<�P ���R7 �w�VBq�R`W�C����#	[�<��UP(h��G�e�����e����u;��g���>T���=�	ʄЏ���5]È_�Fi�T*Rp1�Jk�R,Pj5��ڴ��COz��g�kbb"P�����E3�Du�\.-�\�Н� �-7;��,�e�[��פ���2� �d�E�(H�(�х"{,f���o*��K<~�=��~pF��K�3j�B/�q(�O�����ܸ�"|�,k#¤`�
�Tvai\{͕��?������~�}�� �cj�]w�u�������+��� ��`��%��Ůe���Re��ǶY�b������������l�w������嶿���������2<O7A����{*lšh������'�텆�`�_�\;׾O[c3FG�%v&p�x"�K
V�͙�3�Ջl��(�9~�(1�:�ƌmq����	2۱�"m5��t���Y�T��=��g~��%�f�L�b2�=�\Y�?s���9�>�H�ǳ�D���6�zK�v��C�0��:l�###a������t���HsQ*�!�\��dÙ?kCHs3!�vճ�<!_����*鯂|p?���������E���6ڤ�F`��Nי�	�΀�J�y$'�*���Hn�ߺm��5g�ZT��o����I�S
��Z�}7f��W�*���gI۳�l����!��
�q���hR�0��f�"Ƴ����|8TC�:��jI��ڀȔ���\Zm3�/��w]*��k��mxN��������S��y�+(<����1!�d�Q�M���'�3�бL�I�T��Z���.��CN����c�v����a���Nsht�ך��b����P:(�dFa��ݕ�1f߯��qV�$�?�e:��,-�@��L<�̌jB��5�T��z�l6���B���sY,��,@���4})94d>'1�/˩�ii��*��3�\d���	��� ������0�1*�P LO��YI��� �US?���,��g�b?l�7͐T:g#�+����v��V��5hV�"��˰��+n!l�$B��i,(EU�D�9!�	��FL���[��Ei]{���b�RQ�A �R�yի^�9?�3p�r���NEzq�9���6�<�_T��T?�yo�a�zY�
CN��_+�"w� 4=R]G:S~����|��K/m�zXk����z/V~�7������a�J��6���F"�)i��pϪ{��R��n�~��~�Tq�%����~�S�z������d��D/|���eZ�d�ʋL�r���ֹv����10��{K7@蓌#*f�I����N��ȩ��b�R0$Srnr���#�R��v0���GGaO��n�V��Z)/���C�=��㞚��ˊ��I�d�g7�ݽ{��&8���ʝb��������E�S0��bz�$N�����L2·Lг�Ga9�}}|�rv��Ov��V�K�4�[���*��'8�):��7o�<9	�*/7�'N���8	u]@UR9���A�֑ӫ�j`ޟ���&E=�h"�dL�L ��Cc�zD�/]�bָ'`��nZ��%D�TB��6�j�5�\�/�x�������ۿx�E{�������M5Nl���f#�IA�@�����Ǻc�Q�q�-�KN��e˖���o�^�����Q�~;3��Wz�%"#f�:qT9(ala:��,E��īw���b��6l��~{���;�ˠ�YIJ^)��4m�B��b�II �B��N���)c��"t'UL���u��q8��(R�n�n��z[��܏����5���c�Nꕒ�|\�Dp���	�pę-tX_�8װ������cWlM�����ixIP-a���~����$����I,Sĺ���PA��:�<�ʁ�ׯ��Db��@�^�ݱ\�U7KJ��Wq��֎�Bt��i���`4>��"�JĨw'\�:z���H 5$+ևLU^釈C9��eN�$.���0J�S�D�P�;�hn	�)\s�|�c>�C"���� �&�����奮Ou����O� G!)���M�l���'P2(1=!��nʈ^�:�rN#F23R�W_�@,�����F,�6�������ֻ���x`nJ�F�:=e6 ��iX_��%����@�(n���'��i��0��8 �\��R�#����3-=O��Ny��'@24Z?�7l�Ň�B�#VF��i��aY6Y@d�2>Z� bp~n��*���jaJĂ��4Z;���-�wa]�N^��ӂ��D����֩�ɱ��_.251��Z��:p�4���8�Z��;+&�����;�Q�E�4JI�2�;�JV�_R�!�Ne��AW���2��E��X�)��r�V,И�PxR%������w��m_��?JM~��H���0ZӐo3ҩF��\�e�A�jV���z������.��\{�j�E��������g��n��u)�A�a�J�XsP�lY�g��Wl;��εs���X������ԝaK�XmmJ�gkɺt�a{�����J9W$�˶푑�R�Ğ�B��=�Jd�
@,;w옝��8��1QŴ����7������ګ��{46�+��$�iZ��!-�v9�L�m�{|N'Q|��%���9��xf�=��%��4�����D*I�+H�h �o����s���{]�@����%����^�_�r���廤�!G�B�J��-��P�J�7����~��
�z�j*o	���f�Pm6�Ì�6��Ue��ӕqUs����w�<�<��L�8_",�E��EmC��k��(�:�*h�۟�̜9p�pNb��3�D` s�}�!���;,�6�p�*S��a�v��7�߿�X�ҟF�Gh��V4RΟ?��%�ٴ�]���hM1����h�ͻ׍�QkaA���CZ#x��P����y)�,I�3�i�є��,��M���r��-ę�
�m�F3���cX5���f>wW�"��m�_�<$�0�A��Cen���=Ӕ��Ale
�(�m~�k��?3x�*��O��A�Z��O��e,�.�w��:��Ȼ��iL��&U��\�NE��Ei�vH�S	6e��(���E��w�DhF*�y�A�_�k�y��k�R�7�q%M�j��DZ?S�ǯ���,��3�D���<�R�Z���.qUhN�g��X��/�٠�)�B#�c��i�a}[d Rl�V-cWK��9��m"k�T)��q�P���1Z;�������f�F�Ri�7\�T**N��L�͞.%����{W�6L�l��b����ȫ�ʆ��t���T�L#���5����*%�i�6[hd�,M5�Q�lH�8���޾�-��U�������4`��z%�_�p�����7�S�u��ǩ+���Ȉ��<���Ha�뷀�s|���z?�z0�ԑ��\�e��݊�7�Y�S�!���n@(}�s�#@�Կ{�C�����_��_�F�V.S��V����D�nEɉ'n��������}޳gO�Ĩ��~�.�_��_��G]��� ��-��j��U�	�/�!ޮ�[�Z�G7~�ݶ�?���渎�r���t��d�`��&��a�Y��|y�b\��HnW�T�~P�����O5�� #�0,SXEG+HH�|�����ͽ���[<�����y`�M�}�{o��0dX��ɿK�� I7Z]�VA�U�=X�t�ق�K�,C:�u��X��뗵_��1!P�m��J^^YZY=v�=���Ӥ񌌂j%o�`�`M��K���J�S}�V�Wn������ѱ3�N�!��a�,tkM���Be��\eږ�κ����� V��ҸrI �:ett�V�p}ϴ^�/�.��0]&|�e.��j��&�ơi�5�6\�hK[�����b	�Q�N�:��#G|m���V"�%�*�C+�m_�j%.��{��j���D$��z�ՙ����x��zh�a��,�aP.»U�F�.Z�e��'ci(���E2_Kh-az^�%������*q�:��\�c��|R3u�өeD
r�7h�	]�vA����Ȕf�Ӵ�qdg��An���t�kO�(�Si�d���Y$���n��U���6���)e�������&U[p~hiv&2P��}A�Fjٛ-�3�V���ZN���i�1�:�$c3�xFZ�W�)'�
S'�r\�t� V��%d��ZK���8�CFCH�:<��Wlt[�a���b↧W��@A�#d̊Zf�A4����C۲�h;5�4���3��D�c�5�L�3TPa�	���*�\c=N?��0�#�@�tꁻ�ִHF����F�v��@�q���k���ql!���5M'	��;)�G�{jVly�bf��I�Ih����֞���?Q�!���$��++�e�R��触Q��٧�7�i{��o�i/m\� cO�k4
##�!�v�Ng���ab��P7ă"?�g�~d���Ta�a��x&b6��f��[��rQ���CC�������a,J�MX:J�Z�'ĵX`K����%8W%���F1F��$���q�Ki����AtD�+TL����Gnٿ��7^�x�♓��޽�{���-�wWy�}w�~;�Ï<�����J��ƮZ�*S�@��T�O.�C�E�L�8����]8�Xj�(ӌ�je*�W�s/s��`S��68�{w�y'��^x��E��q$���~�Ǟ��Ӵf�k^�IʧEK7*��IS��ٹ����}�+:a�����)5����9?�C?hێ��3�ν��K��.���LA�G¦o��T9�W`o����;�;Ǜy���V4��
(�U43,�����"N��8eȹ�#P�9U�BY4���A����h3-<�L�9]�8�Ht�۷��-�IS��j���uִ_�
v)i*r3�x���Q����^�g�7z�ۆ��	Y������]J⧹<~vD�$�!��` p)��D��O���ȸ����+Vgj������N�?w`)�^�su8DdM`W�j���c���v��QM��׃OCG�$��L͜���]�O-R��Q���J�I���~��'ҽ��iD
������e����)*��>�����Mruɺ]�܃��pǥ�v�*\)�����&���rQ�F$�az{�����.��SVxf��-��%)��4�TZ���bk��J�����Hp�����"3�fz���j-Ы��G��� ��Vh�"�T�1�g`�	<xA�#��R7�A�ٷ���f)KO���ą4�N1J�r.�ǱLU�V��R�C%����~�%Ɩ��)[Ti��%�60Y��j��[0����+e�r�"��9���~%G�Ć�!��#���[��#6����"�}Ⱦ�����Z��UB,$	-�c�R��C���bQ՚���aJϴ���WD�t����F&[�~*�)�z:�i�4���X�~��y `:��q$�-���_�W�L}��3���KKK"β��E����˩��X�~$	THD�҆�<.�[��$������՗_~�ԩS�z��E�IR���H ��P�B4���1~��.m!3I�l�d���J��,iJ�y���*�CgL��l�9r䩧�z�������6��J����/���w܁��$R�|*�Bm�\z�A'?��ӯ?��?�.m�_�������. ��j���������~�=w�[(؂���g8��Tf�|{���Z��W;��=�j#qj	=A�GP�Sy�܂]*I��!��z�-*o�%j��~���r>���jV��_}s��k�7LٱĞ=��>���͇Hn:��Б�*�=�%�Mڍ!ݡr�g9$@�?��Hה;��x��H}GK9��Vj-��$b�D��]H��?��ќ��-r� �.G�&��&�׹���s���{���Bq���BVe�Y���zڭ�������'G_0��8����|���� ���Q�=Q�FA���u��gԢ���i������M�1)Y���4��x�.�8s��Yqv��69����"d����Rl���f�'V�_�]���<�v��mt�b�v5�Yݵ����H�Ự���:z����k��Ў�RcQ��D�;�SD$�-$�E�����Rq(�:��7Vt_/9 r��N�4Ll��%-���]l�Z�
;����Iu�O�w�4Z�ܒ��;��H�"��d�",��ⴁ�J�]Y.r�u�5"�CxU�Y�t��p#K��-B�sj`H�DMB릲�tH��l�ԇ]87?M��^�>�u����;N�.�D�v��	���^�{�T"���1�R��W�SUa��BJ��t�	I#,��))x��s�3�[fl�ϥ�T.�S�Ӵ��d�˰�"��i���	�pdMЙ��f�*��ro��܄��m�ϑҨG4=|�Q+�nEZ���i����I}�(�����2�"V"-�$M3>����$�I��������&��TSqtI��j���&h0��&F'�˱5�J�N��o߾���/]Z����~߃�V���2�`ypi!�����V��&�526ܢ�~`\׶B�k�?=�8�ef#80�`��L��qf}(�r%��6��4ڷw/x�$��L"��\�9�e� ��D�؍6H!�l$�t�j���q�q�47i�1���GD��S8:B��0�SY�T
��Ƽ&� ���6��F�[[�K�Կ��3���I��p�Bg~�����s�5j�P�z�� C+	w]f�O���3���i�`��Cٔ������� ��������j�g!�l]Q���Kc���Qb�������o�����g?��?���~�٦a���������|�XpL��V��9n�+�~Tr]�c���G~�#_�˯���������ן=}��?��B;>M9�k��B�rJ�o��o����4u�%7)p�N��5$�*�2_�����z�x縁c��������ҾT���,{Un��+n�o\l�%%�"3� ?>>N�N��CϪMN�!U�t��{lzzzj�>�8T�����v��r�T"R2�)�$kkk$�iwg�X�vZ6���⚹�*�D7�Iر�^����h4���O-��3���ֵB�d�,��+�\�p�>S�T�U9��'O���;vlum�6��O��!��.�X��!L�ySD�[	3��!=�9�R�w'��Ç�����%F{�����Hg��r?.�����������]�	�22����V��Y%$����4|c=p��3{F��`%
��F8;;;5<A���ك�1s���kZ3��άz�\v��jwc��*�p�Kf-�%s='�Wօ�MU���ݤ^K��*�	=˺aN�$��U�1�%g�*�Ke�0۞�*T)y�s+kh�Ѓ��U|+�jۯێ�'mp�x�vt��w�_�[k���٧k� �XB��Z��ze*�E9:�����S�jW�z��H� �(�T��So�~@J�G��e�T�%p[�Ҡ�N��,�&��D�xE?:7��ĕ�R�$�۽@�_�\�`�hJ������E�=�g��YU��_�r��3�x��*
��K=)cMI?��}ۡ�G��H�c�t�/*4}`�W�wB�v�5�|���������B�4F���T�i�0z?~�z��ћ�����՗�\A��I���:M`84^w�y'�sff��D4��͉vfxȵ1�����9�4�5���t�M�q����A�M$�T�@�yZ�5��
vKND�����P�WV�U�1��*��	��,m�D��?����,�@������a}�#�t��I�&���:�[����W�����/��#i�fH����D������G����W}V�A�/i���Z#[�w��D���c��k�����'�> ���g�0�4����_��_�/�!�׵���R��YQJ�ߨVG���/*�;��;��}���lT�Je�3L���~��>��O}��_���h�ۆ|�+U�@�M�l:o�ㆱ�`����/��+>n�↚tś�>C���$x�~���7tCq����l��:���\gz��;=���zu���&
�ENR�2��)4ǀI�tt����I� ��PS(c��e���Вpܝ`M�<���e��_ݽ�B�.�_�󹛖W"%a�nuSsݵL��mʸZ!Ź6Q����P+ҢC��巰PK��OZb�P�g90�j('��V�,�+g��bYl�q����i�����R��A�������$ip�V�O���q�-RLG+�3Ξ=�|�`2TV1-M6�V!'n���� ����.:��9`��E���å-Dc=T����A�G}bπP]	�c/�R����eZ�E����b���f�o����6L�EW��GF̹^Җ����#��v5���pr9ٽ�r�=��\��Z��β��rk�q�t������H_}	�}d��]�z��\m?;w��c#�r��ꍢOl�1�bЅ�rU�H�^���f�Ы�te�-��@�?]�� [N,�̌A�'�ct�}�L����X&5�v�B�u6��(�/Lj��A���f��i�!����h!��25f�*�ΦM:4DB�k�A�����rA<:[L�Z*��K�[|�2�`���s��6qxGPg m蔍v�g��^/��0�@��?\�4Ktwȍz�T���:����Ag׮]E��{1�+��ϴ� Ew:��-����ZѲ�]'Y���b�⭶Zj����������J�Ch�f�˵���"w[�� �6��w��Dl(k�v)�k�ڱ���ҝUuA=������8ib	gu���_h�$��fD��Q]&H�04�.ϰ8��޳[�L�h9�#�),C�ȃ�]���[iF"�')��Rڡ�\�J��JĊ�#E�6#�)e.���TCB�u��N�V��z�n/�w�~:�⥋/�ط�����^;�ҋ'O-4�I��3$��n���nmt�@���*�N0�fBX��i3CF��}N�?BPn�3k	�f�6�ZK����U�/�?�4?71>N������r�B�0Oű����tY�\4�X�LҨ}�
�����'	I��������,2��������,]��>x*.i9�������1Vplݡ}��i5�w}jz��f1���TSB�GYq	��!9y����3�8RWE�O��jo��uC�N9�7��mq�^�)�ԉ��2;)�jWh� u��!}��`x�>���}_}��JEϩ�)�7ǵS��d�������?��|p��na�������G��GC�C���qDj&���텺����������J����gN?��_�~��c�4!È�s�?�=�������'>��{�R.q "�_��+1tAS��.�k��{����������ި��S��`�mk�jM����s�F[��z�Obs�[��ͯtw��}}0W��ϼiko�������9*�&ɴ����X]M,�b�' j?b�.Ϻ����&6�+��p�!9�P�"�|�7�]���Z�V*���%�U�VT<l����{+C��_�%�dX�+7�/}�K�s�[�Q��.����]�`�uk\\Q<ǚ��$�����<�(A�@/!�Iό�*߉�(:f�؏�������	�Wאo�9쓁K�.�{�F�jx����v{���~S-��$��:�>��?M�Ҩ�0L���*�Թ��52�DAǞ={�R��n4����a�E��%�$����V_A�+)i �����]�
����=�0j4������~'AZ�_F�{�)'$5�{��{�Ma^}���[o��z���tg���� bx�67���0�L�"\���0�5��Pta �=廃,��‴Q�d�������2\�80�v�Է�Y�^;Q��lԘ&8<��f���-r(�ß� i����&�*釲Ǉa���F~1�[�Z��v]�i-�om���cp�����[A@o�.{4����/>�M�gR|��#�ߊdQ�\�)f����&X1���mό��v	=#GW�pa�=??�m ��\(�����c/b�r;��e0���;�yl*�#�4N���h�U�2s���&]Q�~��f�+�=��ͅ*{��7�^�c�}�P���S+�Tw|�y%x�E��J}މ��5<=�S*!x���?!+z��Tf̣־��Ju���@�+���,*A����ȑ#C#��f����e�+�4iǪ��|�הU��`'���H���"���m	��%�..��Ţ�C�Z�hnУ-]�?y�$���{���`#��� �Bݭ~-���v��qD�s}0��>{҄:"5�${��q���0I�d����>a:La�D}�ə6�%�민�
��hќ��^[Y�[���MoG7���
W\G�tR��>��N�7��\���o��^�E)reǯhl�Z;�HТ �e��Բ���1���p��a�o۶�C���xł��Z͟����?�HLu�$%iϫ��t�pŢ���C�H`����]^
у_iw�K��P�(���g��v� ��wP��8�km���Q�:�/����	!�v�k�a�!��m�KG$��|���9d�YX�S�A��U�W9��/���׾�����M���kí�Y����l�K�a�tB5t�����b��<B�-мY1�4g�\��[\�Դ�^�k6��(�'�@כZ�t�z~ca�����~��ɻR�=�@���&Ǵ@�1d���$����?�ǧ�s�H�G*�#���u�T��攉>�l��A'cݴ�2=��\��@g�ilx�˅�"��e��p���ۯN(��S��V,=Rl|�K��c;�V�\��ss�~�����d���\��I_!E���$S�o���b7��u�)�� �F;�1R�5� )����`tXr���O�쭑&���*�����#\�R�N+�ir�D//��F�^��
��R�T�娳kt�f�AJ�L�iGO]�c���J;v+e�a�pQX�/[�!ʹc�I7ҢN��&���Wg{�x��P&4=h���W.�S(�Z����y�����)�e@dM�6���0� ���(a��3n����6�%"��kdC����&R3	F�c(�cC���1x�z��uzq���7{a��"ϰ�&���� n�d�.%�,Z)[Bd,�7���=Z�e1�y�*��d\_��W �Aۻ��帍�]F\��H��
�/��۩hző��]��G'�bx�bȄmBL�$h8�J� N���$6�0����l隍��ɯ~��N]��륎�؅b`����֒&��@^� �T�.���%G&�\��\�(/W�W!S2h�d�g�Ei�G��6��Q��1Hb�G�߈��7,Q\�2�8r̤E+?�A�Ħ%O�I8$�%�D���B9�-0��RX��LF��	�Lu�
���YER��2��`�8������e�C(�yS���v��XF`��,N|������w���}��k���$��ݗ�������]wݵ�����t��jр�`~�B���VsLyb�YS�@yS��(�f��5�4�d��U��$�`��p#�r'�9���Jl̢_����$�Li\�p���Ʃ��ScC����I=.]��Rõ�"����е$�9�1<T�7]}�}��07�o��I����.�+����_y��_�z}Fha7J�U�lY���ť��S���
E';�f�-&���f& MA�Fгr2��e�ܞY~�wx\[��!!�7.\�A�JF�z���`���\�W���_�Ri�J%�$�x���#�\eb'���o�����Z��~��&'�¦"h��"Z��P��$2,73S��${�LM�(�c��AJ2�J5���5Y�v�d���l0HW�H,� Xbs`�T��@\	1C�M�-��S�9p��������o�I�\Nyܵ����c��p�MA�6�¶�'�"�v����\f���W��gq)W4��7��S�˲��]v��n�~f�zބ���=hd��k���7�)��wಠ49��U������������ʔ`K�����mF��I�-TK�+VV�H����0"�� Q��ҥK�էI38z����]c��^;��ѣG'�M�hK���_5�M�IJ�S����I���`��U
E�U	a����O����7���6>w��p�r������畷�.��4X�*��>�|(q�#���#����^]]ݨ�I#d��R���P(:tH{�
D�p]ڈ}�*�I��UE�R��\�+�`����<����6Ѽcw����/�333��ts�vت�����{����H�A����?O7	����Ԓ��v�޽{�H�>��3�����{��Y�Cz���}����#y��ů_8���}���`2t-z�MC����y晴��v��h�Vj�7�m���c6BԔ97��"�S����w�N�۷��]Sȣ��g�n�Ma�m�:4��:��K_�+�]Z >����L�|[Ǆ�Q�,�%0��g	�k=`o�C��q~��s�[�f����r�r�7�8�>��;D���uZߟ�_�Z?��^���i��.\B�T���M�%�����&���\ M~���fl7H�Ju�>�*�o���7��zcuP����9s挡��[��m� 零~��8D"�l�q�3���%�l��l#:N$�Z8jX!��~-�הyP5���We�[ŐW�p^,#&Yc����JqQm|�]���
�@��!#����p�$��]8-KE��!r���q�2䧅q�f6�L3ٻ�����e���ǜW���{JȨ����/����K/�D�<�&XK>��O}��|�خI��(%7ZBq����r����0�_װ��:J���[��t(����B'�4v���H�8���ҙ�u��y���q��$�أ�ze���W����Ȗ!H�����_�����3(�����7��n���?L�/BZ���t�sǟ|�ɑ�ݓ��<� =������^V���.+�$�����R���ӿE3e�o��o��mJQ^I��b���-�j�#�}��R4V�W������Ҝ,���{F�c�s_w��MQYB��$����8���<��4
C˶}�=Mѥ�����F"���a�إ��;�,��pǆc�.�(�+@}�����b������_+�d�G�f�u����uk_���n��=H����m۔�mu�r((�������[�C޿�2ɞ�?cp��O7<qp�N@�[o����#�=�ߊs!��G�W�~�g����|q�sl۠�z���F���W���툭�0+�e7�ϩ�7�e��m:֠��r���Z�	s�,2�d>�P]Eڦ9��rM�P�0�3P�n�9��}�d�?�s�-�8 |HQCj�ò6Z�^��:9���[�;V)酧���7����[�#�[o4��'�x5�z7u;w�q����z��m�� $���qX��H��u�*g:�t\��A�0$4�T�W�P��e���j`��䭺\,ѴYY^���������D5�7p=HF��H��2z�n��Ē�iR��T�B�� blx���e��-����t��筯�ÛW��kt�ŵa��5I�J�~� l�VA|)�J�t�Ru����nvB�	\=��������5���o��x��9�\�;L��t���kN-.ځk4DRu�N�H����Ө+]�N9$u3��k�����
Y*[3;-4*��Ϟ�Oã�{Ğ[�]��v�����<8?:ߡZ����L�cDa��Y���AD2긊N ��i?a��"~I��hF�ơ� <S�X)�_�0{q�F�sj�����÷T�v��8y�MꜿY(��l�z�C�%����?���c�q'�̉�<~"NWV�N�xʨ0��R�f���8*N�5H� ��%�S��P�^9��$�r;�t+�0/��X�j��YWM�8��u��$�:��<H��ؒ�f7h��,���a��sgc��;��	1�!����.ߥf[��4^��/l�Ma�a�w��Ҷk�rd�6���'O�,���҈T��&���`˪�ZA�*�E����
Xr2&Q��g���Z�i�2L��s�(X+d[�*T�b�Q�t&�TT7 3I<��*w�e���;��u��^��Ai�\�Zm6�V )4�]ݭ�6`J͈<��V���n�T�m�%+�	-�ۋI<Ҽ4Qw �o��&5�D��j�~�͠/2ո�Z',�FM�
�=2�3�&F�D�e��^��
}�t;����u���&�[;�c{��Ñ�wbp���� �_���מ!�}���Ge�//q��b���$"���50�ƌ$IH�#a��W�R�M�PJ-mw��.�����0,�i(�-�ѱ���/���7q�G��]�H��Z~�����"�q��ٵ���k|t���3I�8n��m��0�CT��z�҆������ų���q���8�q��4�6o��X�:��g�W�4���M��[p4&�H-ԟ3�0R{���?fd��e�L�sz�!�ܿ=��]\����u��+��r���}W�c��[�!T)͢����m���m\Fm��w��Jh��VR®3�[����� N���2Ȋ	5�cV�_2����	��������Wh�=�q�Х;A4�CF��ao��� vZ�\�Z.� ��ve��68.�k�Ł����J�s"ݗ���>�����!�m'�^q9�ɩ�2�w�v\/wSr|������w�?���Ʊ�M��*r�S\�"�9;w�Y���,� O\��������4�r�*�6��!�5�Ď9$6��;u�������)]\ޥ��,v����>O���ef��l��/�=W2��(#����a���I��Bfմ��gi����wiQCc�t���/#k�T�+i�~ꩧ�^�k4�66���a��f��]�������X�()f�k�u�.ٻm-~u05���&jnT�������׈�%3�il���3�z�@�8
(k��Y]!$�^�
�w�~�?qY��Z��ܭ���J����HQk4�V��)U�^,�A��7j�Z���7��H��6�}3�F򏺢��lz��t�[#�
u�w���[���ȻX�ŦBm[YYy������=�U�|�djCC*?�uA��ٴD��<��QO?�tw�<�U������N��'z���환�����e��C-����|ط�\ee�N����@�,Pf~�z[����������j;P���C��<E=���*�3���{�&����XêGe3�����'N�@f�|�)�A��z�#�^��Ie�mk�诂���崜�G��w�u'n�����ΕUƣ��r5]����o��}��nm�Y���*/r�&�k�@�i�UR�ӊ�Y�i�U*䀵Z�ɐn�j�t�p1�z,�J5�d�52XYJ �1(c�����ݔ�F�l��`�v��S��͵�j|)Ѯr�T��B�qߚ��v���t�M���I.9���"E|)s�'��n_W5�P��,	T��ګ�v�k�}6E�^����5L�˜+��2�@O�,#>l+ʥ���	�^�Gq_�ص�KL-����ُ~�رc/���
��޽{���/\R]=55���A��4���;2���M�MAg�Jk3��%X��{YI"�\+�.>�$�H8|�OPcJn��_���c~������=w��ԡ!�H�\��o�Z�tř3�)$4K���C�^��̅�Ǐ�N@k��W�����͹5����y�$��WV�7��.�8P��y�&�q�������`���C-��\sU^�ɿ��j��Nm����D��d��_D�h�n=pj��fq4�I�I��vO�n(�R�K�+U��h%�,���
�I�ׄY����X��s�rmq��K�1��� ��Ǝ�¼k�mE��B�ć�N���D1C��x�����<>�����G;;�έ5�?)/'�+�W<�����|=���K�G�l�~�#���3�\�����J�U_�k�7�4�u�6�"�쁏��51@�6u[��=[�k0���7�b�ݷ;�d�kx�P�+]��U�X\#7/?7�FSUN�f�u@��ۍ狾�A2ץ�L8�}��P�o1ւ���S���n �؊��ʈ����uˑ��� ��宜�HJ��ɳH�k��N�%}��^����/u�{�G>����1��*�$zQ��H,3I�Ė�s�k��U���/W��T����E�"'� <dXVmdd�ԐW^���>|ɲ-N�R>d5�RGhD���8�͂͹�z�y��R�t�t�����ÇI�U	儻6���ɱq��g�yflllzz?�/tZ�b�F�Fߥ�ա�������|��I�UƸίII%�1	��vt�T�H�(X�vR�)��B�?�[���!�l|��V������Ȱ�԰
U�`Ţ)z�S>t�)��B6������s�A�S�ao4�ϭ���!Bs��cGQg����x�u_Y��r��n�kk��ָ�h�ic�].J9ZPE��Yi[~�JXD�	vB�r\O&��Ͱ�u �Wj6�v/-���v7�	F�SV�lP���=�H��m�l��7~���5}h!�U�Ž�Zݮ�ө��]��6�k��-�a�t�Y耯\��z}Y�h�r�fH��Fΐ���qǚ� ΙB�'|K���¼��|ٔ�,e�	��%s������8
�e���~��Qu�n�*���r>��;Ϯ�̬/P��C 烯'�7�V��7������`�`�q�!h����;��P_#ezed(�n�N'� ��-��%��Q���h���j��8�>��gb^!u�d������,�������Z0�+��W�2O��sIu��o��vL$J�ӭLǃ8��Ќ�nb�c���5 �f�$\�w�E����G�Km͠��rii���i������y�Wz~����6\�����n���؅85T��"�4FȤ�c�e>dr֔,��W�U� ;�*:{� u��X�
%��d��"�m�ĤW��77���4���N��.r�R-�5I2����ĉO=��H��������T:s�̅�K���G���'��i�={v���h7��N��Z��J���d�#A�r�kj�	����lC6�m���0W�\O�gI(^Z�%1����Ţ��F�Z�,�է�u�K���{?��K/m�w�c|���6�.]�f�k{�-��C���ji����M�/u�]���c�A�����j�������S�<��basx��;��h$���4����-$G(H�T�_�#�ST�F�V����F"�S�`��wM]���x�3����ڋ�YD�aʺ�֚���N� �ݡi����9q�#a�.������,a\���࿡yj}[Ůcʘ���$PIX����Lͽ>�4�?�ul[�		:f�ش2}�Vp��\�LZiB�]�M�����m;�Np��^��H�"����2`s�$�-o�I���`SW�W:� }��9��6��[8�w�b���A�C#;_a`�v@��^,e~S4�t̝����,����R�9���-�~�Be��O�Ar��G�4�*��rOW�շ��6�c��V��r�K7I�@�r��f���gi9��8i����ow����(��n
�J����\�M{�j�߿������}����7��q��:x�޽{�8�:2�˕�n���N�:}~�ȑ#�����].);8�M}+�'Eͥ�U�(&��<ԋT +W�d��6I*�oZ�9�Ф����]in*a�����2�^����...u;j?���
���U�+z�z��wz?=exxXr������D>�fۧ���M���DF�:�O��}��&�:�Iy�8�g��8���ī#�Ѳm��{���;�#X�����)�9��h��jf�V�����s�Q_-..~c�}}�'P�����R�ip��i����ϔŦ�y6��~e0-��/�>����ѐ��������*�{Lhih�ځ�K��P!�*y�e\�m�5�Z~����ѣ�=��tܽ8G��>��3e�TÁT�����ɓ}`)��s.[2���%sC���~�gj��h�w94���Ch4��iz}��N;�Q��61֗.�5K!��6-pV\B��@<a�եw���$�jr������{Ƈ���wU<�����������M����2����_J�28I"�q�q��X U�o,�tKmX����:�ө�U/���W�}�<�K^�6�ݎCw���5��b_
M	� �F�u�;��gs��R+I��Ǉk�pqv�VY��L6�
�D�Yj�e~6�AJh��}��kB\9lAcv%P�Tq�*"����&M��fu�,�܏��1���E��P�<��w������̥��4���/����X��}��yBe�4��K4��^(�Va�T`c���kr�j�����pvvְ�%�5C�z�ŋ��P1ְ~GGG��ٳ��O?�￠�-T����X�Ȕ3���PD7�gn��g��H��x���-J�|��_���$sP��4�'vш�,F;i��.�fJ8���S��}~c�z�7��6��ĸQ����w4�F�I�[��`a�F	��@HH@K�ARWC�pP��ʚ���>Ӑ 邠��$)����
�{ML^�Li��;L��#�"�Q$���Ny�6�6$�i�4m��=�,$�%�N!ьT6uG�������J-� lЂ�u���ٞ�IۖaŢ�2NL�W�ۑ4f�pD����&�%��ˣ�R	��S}��G5�7Gȣ0A�@٤KN�J��)�F��1�r�ً|GTi&$�D�����l�A���؎����J~at�<�I��C��e�o:}vX��)+H�
�I\���4	�( �J���J"�ɥO��T�':	g�;��t�LHi�^'� ���i���.�ܡ�d�9\*�&��Ű��'�)ཅ�E�:-N݈SW�	>w��\���FAv�:Z��[A/u]Cr#� ҝ"��8���Z��u=oH�����al�m�RnK�vx�H���Y�v��ݐz2�F�6e?�Xf�摄�u�&���v��2m"�B�z�F�x@�A��/-x&J�J���3��q��I����CL0�nD$����YJ-;!�⹴ޓX��i�4W:5F
�l���ǘ�A6P05�%"�C�2A�^���F�EDנ�Ax�+�E�7�U�h���$�}��@�:��hUv��T�E����������S/�ص��W^�X�����Ҏ�M?�u�Ѡ�=Ne����\'mlj������t��޽�Ti�LæE�2؆M6&Q( ������t�,e��ܪbKm�C$�8�N�Ek�Gc�����4��OC�%�2B�$�����M(�~�=�K�!iH�G�RT*7ۭ�g�9v�����ӧǆGH˹ta�����i�lue�4���åKs�{�!�f��׺���S�9""6���ŦcB ��IK��K�j��L��J(u5'�.uN'.Q����5��.���x����j��9%{x��n�jrl|m�ҵh�*�� =����L�8R+�9C�pK���+-��1)R$�H+ո���!i�� ��+s�jS�vӭ���>r�,�Q�m�5r���m�1�P V��|(Nm�ݠ,����nhiI����m�z&W�a�z���D���'����`Rr(�D}va�Y ���������5�vQ��I�n�����������p�[c��9�D��@Hj��Qj��ޖ!�(h�`���T�м�8�b�ͣ��Ʊ+��$,'��o�k�L��.�Hu�]S����{�K�����3�`�F��{�(�/<��K�_yχz|z
J��d���מ�uטű����6�GU����z��=��Iw;xh�9�m�_8?2���I}f�>�Ԙ�oо�Bnx�
ب2%KEԣ����7*�ʐ��4-(�*�0��Va��`�MXpҴ�QG*�e��������q��z�ծPd-u7i���2r�W6}���&G��z�������z��N����؝�
-�x�R��棏>����=Y������b=B��V-��b��<�;¤�S��4C�Ą-�pʒGd) \���RM�^�a(���T�i�:Vk�
�(��^s}ӯ��b1#ڛ�xye&�S�����޴��܁���]7<P��}���m��r�-��k���8�R}���^|�g _m[���E�uhqK�W���͔P�lS
H�r�V�o6�4^�ni���������пg�~����&�K�R�F�������]��L���O�9��rux�Q��`wp�":�Ĳ:<F���J��}\�N��vvv���ł�F�K�n�C����p�f��ӧ.]����{��^�={F�z�+A[D=Sw-�X�W�j�%\�D�PI�v4�mV����$�Dl	#V��y0�jT�>欨�g��Cd�fDPVuRi'f�XK��hL��W|��	�ɡ(*�	�tU���� >"���쑒��QXj�H@�nf��/�(4O��lѡ]��q ���ig��&]��1��,u��R���2�XG�Bå}����NV�T~!qes�J��'=W�XEܨ�~*�ˠ����;���������Y�����G{WY�M���V���p=#����#U��3��$�
Ǒ跌�7�
�r�>�t�4�^Jv<�3�)�����gl�fg�ٴ`���Zo����m=Z�*�{��߬�́��Td�	D��Q1�ųT�@�&F�ۣkhc���Hܖf�����$peL�B�*����\���*����m��h��R.5����~,��Wh��%��!�F�!#�O��8~��LH�g5�)a=t8>��u�J1"Y��<��SAy8OR��M�A��ó��;�C���#���-K@K�}��&Wχ��5.���֕�~�8 �5`�C��("�Co��G���ٶ͆=�F��3�}i9�(�����\�.�6i@���J��P�);=L�O��j���.��~ Ci¼�LJ,�r��gl�4"@���
cU���H�I?5II�R24ڤBA1Ę]�n�68J�L��r�'�-�%�`]���6ס�'1M_"`q��R9tC]x�U��zF���Hg�$փ�Fm��bz�-ٗO�U�%��r0P٩�y/g��Έ��[B���ݴw���<b>�\�?5`{�٣��?��L�"��15Rk���o=���Z��d��lll�� ��X�t�[-J|���Dp���߂�-j���|bjP9���	#g��j��}��/�G�o�Ce�>i3��M�\d��T�Ǹ�u8ǩB������ ���U��&��aR�e�Vdw��TG�%RAH���NOO���sH�5l��m�T]-b��0�NAA`��I��E>�e+o6��̙3O?�tett�ٿ��C�v��m2߀],�&�Y<���o�����5lh̢֪�2z�]�v�*5�rxx���K��d8Z���FJ���_�_��b�z����%�N/~����s�&'wQ��2n6����m����k�VQ��
Jz�n�#��e������-����W^��W�����z�����BX���F�S��R��#����V��F��ř��աv���T݃����P�o�I]�,��&Tp�> ���Sj�]�H�͚�]�R�������=�;�UI�ցf3??O]��G�v���_�n����5�k	�&w��Kp ���"mX��jآ��csTLLL(�<����<�Y����S
�E�G��T��r'`,(T�]�)�0�B��b�M:��A6R�*�#��4�h^�MT�&�	�	X�p)<�2UrJ�R��>�o�O�JwTM���>Ә�/�[�۷����4�'&h(�m�4K�v_Ѧ�T�$���7�|��ҋ���2�n��/}���B�� o!W�Ȼ��Ueª�Wx\�<ˉ⚄*Y�^��H0o�Ɍ|7#g�F��VV^{�5�|���OMM����?��@n��?���7+�XFM¡!ZSe��{(�&�l&#�<�q���'p6��cM�z�����쩽����9��o�ByS����
���V�\Ze�1�e�ٶ��a�$z�r٩��ت7��k�4f/��4K%o�LG�ƺ���nee��lG��k#��P��$ ��H��0�[�h"�P�+f���8K��A�9����n�4�rF�j<0YݓԞ^��!�ܭHx�w�Yg�\��C�&;�-�;�:F�=��	�M�6��8�YYF�KJMi�OlO	�Oo���/<)C�Zj�����+�b�T���S��U�� �ш��!�)��J���rz�O�}R�"�ٰ�Q�aB:��'�+�?�5������IF.�`����%�9r���+��S�ZP�u߼zmRvm�E�����A�L{)-WCD5�c�O۫2�M��	��nA��ri�����<�*0�H҉S�vB�.��=���m�'��ĵQl�7����+c(F�2u�C
�H��@kŖA�%P��cy]	��c&�B�f�$Q;��C� �t\ۢ��"+AUK�U��ĆpHL#��fT��)��	��fb)��	{ПԶ���CT�r�<U e#Z�	T]��hi�Ds�pNg�s���
t3LE�#�5&�><�ЋDa�+�[�K�C](m������aqN3�F}������z�Z.	E��"�g�T$��bz�%�^^�рZ�e]�.:�ѩ��<@���`�@��)$j;:E,u	��up�U��zeeN��ף��P���z��a(���	R/�Z�w"|z(�I�)�=��|�	a�X�q�	[�-���JO�F����$vBU�	���m��U�VB������-܍Mv����I0=��i���@&�^����+Ն�?�X���t�]��e��M�i���G?8t`i Kˋ�$5�Ԑ����5R�]�sKEҀ	ڃgl,\�ֲm��\��D��P}&M"�F����--��]c��G�foiz�R�Qd�gĚ�P�Y���#� �kA���T���9ph?���z�I(�ł
���M;�Dǎ�C���z��e�+��~L}E�^U_�<r�Ⱦ}{i�\���L�S�d�>2<H���4orT3�»��&�W�gFǱ��"雯�Z�n�?��>�o_u��x���܈�z}������/�����7�6����+�V��+��˧N�ҏG`��=�}��o���y�a�ڰUuC�i��q�F���}�������ݵ�1d�L����)u"�3c0�8���Q��ʧ�ƂF�d���88a�����Q]�<a�����s�M7���{�e�\�z�V�ҥK���w�}˗f	[����5�J`?��ԡ#G>��sD�٬�%��l.,=�䓋��XG���L��-X{P�-��LIl�3���a�ek335�̌gH���\��ձ�-+g�����&j�k���DjVp
)�c5�^b�/q=�����<�1��M�!�P�gYs�3/Ϝ9����g�1�L�[�l�(�f`'�W7�~�[JU(�+�i��h��n4>8:\=7s��j����Sv�%R�6�F����h����l�OT� ���-%��t)��3V�T�p5�
�� 0Z�t}�+!�z@k��N��]	�J�Z���:6�G���R*[�fv7����հn��\�DZ4{f��oR����z�kQ���.{��DhD����-�7�G�ݩ�?�CVQ'!�0����1L�H'���/$}Vz�e\���vd,�HtdN�:�i��������)`�ō�	�����V�<4D��~�U�f��ؒ�¹$=v�����/|�E���R�VA��m�N��t�N��Q�UHc]k5�?���C��ײ����kKd�U����-��[�f�H��{�s�=G�U�7h�-��n�762t����^%� ��yK�:^���4��877��E��X���%�Hn7Z�����q$�� с�Ö_��ٍ!���^*�C�\ڵ�b
�8�H7��L젅b��B����!�Fr�����qMzpv�5:[u�m�Y�3R�n���cjH��/зI�a|kؖ�����a�E��`xH\�����+�BD	�/1�"�8J,��X3Bϲ#	"�uJ4��^�NE�c?������rWyi4#�CA�*s���Z�6F�ށ�K� ����E�C�P��T����b�����3L��42r���������3;���sM�p���ݰx��^�eTj�ϝ���rv�"?\�f�5L;������U�8 �D1�]5��?���fdV�������|���я~���Z���jq����?���O��ϑ��lg���?��c�ğ��I{=,R1�Fę�r�$x�C����3�?�8�\�y�Mh'�t#��0E�K/���G~�ܹsO<��O������,�β�)�왙Z�&�������~�Q�1h�:#l�1k?����_<Aw@0�LFD:��_���Q谿H������g�x���d?x��ٳg��]m��Ç|����s�@,�2�%G��\/�U��ǃ�ï����o��s/�JZ���F�����瞇|�_�3ڜ>�����>Fk0J�]"���&z"�������c�:�~Q����{I���W��ѣG���b���?������1F�1����� ������?�y�5�Ǐ�7~��`e���R@C�xBQ�?������I���Sp�.?Pk?��?��g�t���2�0	��O������s�HH��{���t���>Bc�5�"��G��'�����DOc�y}B���~�k��{/ur�r�.��_���퓟$y
���$m���{i>G�?�}�/��{���~�����^58�H�d4,e��1ٲfmQ�l;���$�x��SBa�C�C�	h����n�磎����R�����}e�6;��W��������W�E��>H�v� ={��}}~q���kkk�ёG}tm}�O�L?u�#�M�����:'N�8�ҋt����d>�����׶J�~L<��ʁ}4s�J奄%L�'I{� �Ui0��	}������x��ZȊQ�ZNp������'�]N�<E_����6��Qo��w`?�[�.\���|䜔�p�l46���x졍XO��c�%v,���Ri�+CCC--K�P��~�";����������w����3�$�TH��( �B�J�\��U,赀��kA��> *H�*h����Bz2�L2}N�}����:�d�}|�����x�'LΜ����~�~�վ	�8s&�mdZ�TO��"�L�k^�1]f!�&U}������?��!О�"��0՛��k�iyJC��QEk��i�oaMg���J�E`�0�9��=υi���;�:3`We�X!W�-�/��2D?q�<�~�;,VA��o:�(����c�JrFg7��w��k*���7{�R�l��f��<0�㖷o����_#Ih7��sW�|*�Q��ꬿ���"��_I�=ǩ��UBx��6QNʍ���vʇ���`�{�9��Ʉ!�ټ��|ac���h�l\���QȡŖ�XPY�b�� b��`-  ��u�tK�"W�P�D�,[j��`:>��Y�S���~�_bYAب�-+7��L���.&�?Wbh�Ƕ���>�+�(��(��s�n^�=qM�d���MLec�ʪ�N�c������>��R��}�~�����-x*|�<Q�PA@E��-[���d�m|y�ڵN>���27f��&�F��M�V��t��W/��)ޓfp�T���s�͞={��MX2)����t���萐>������U�c�x�	�zr���qX?�NT�51A������(�We��u��Թ�FSJy�(Np��^ߍ�����{gRfPww����wl�)�;X�R�x�?>d����V	!b��>�Y���(�^&:QZC׍����E��-�5��1�M-�ШV6��$@aFM�U�	�#�:���� $Ϳ�ק9�O��ևE���J
�p�&b��jK��f�s�GX���'R���5+�Z�tժU���:���Jއ0�0)�x+��Ǒ�3�eHwol>������%2,Kn�L�R�N�7�)zlʠ�D%I����-%�)���t��ѭX,%���e��U��IM�jJ��/Ub3P&�%_78W�֗�����d�h�E;t)�W)W���"[M28=92��g��S�r���=&�R�H$���k+a���'O��S
���j����I;���*l֔ӷ ��8Ո�11������m�����G>�� ����~���\�wk�s���O��� ����G�ϻ�Q��KL���DSB��`��>0���t)����{�?1mZg�W�j��ǔ$� �Ai��먖J��g=�䓇t Լ���)W��U� RjY�<��#'�>����f���A��n�����I�V�G;=hr�}wC��_z�W0E��e�L�9u�>���￟��kD��Z��+�|�3xl�ʕ��(k1��7ˮ��5h�Ɔ	<��-!�S��u��4u�+�xa�1�(�m�(Rsf*�© ,�!􋦇�d6@�#-Tp~lہ]�_���_�~��:�:����VEK �"�@j6�ǯ���y�ݧ������$�0L��F�]G7ØВ�)N��܄��	Lb�j��Ф7+��DI.�P2�z�$]���>��+��v[ʶ6���h���פ
�M�&�e�F�ʫ/oS��}���zc������Y�G��L��t��T�f��=���\�w�y����߼��_��-hD��R�gp�͔:��0�ʺL�i�Ԅ@��!?0����bevL��7|Xr�N��jjc��8vj��F��]%�ɿ�Q6'
�^]ǆ*F�?6���E���.�(��0692^��w�tI�>3<2�e,��c�u�RD��{7$����Z	�|�S= Gr!�B���iϧ�^�ZP�e����;�ݖ�X'�=��ԗ$? ̲�R�8��e>�����-#���$�C�4�$�lr��iՊe�1���� ��6�	a[Q+O%�W��BC�3�p�Rbj'&���]�rq�TĦ'/&�BQɛR��/�X�~�0�z_>���ȍ�#�p�0��nʹtUK�˟d,��P��T,�AJ)(*�p�mK�
�NT\/�jV�Owkaı5�l-��Q-�C�ڼa��B�p}��Ќ\> lM������La� ��,A�(��A[�g�z/��)�qS��b�������D3��ՙj��jHЭڒ/W������`�Z(��u�x���{�q����޿���^H�R�����*��	?JG'JӦ����\"Ƒ��um�P�&�c�?_U���Ħf�V�&J9H���j�9���dR�͔-�9��dg�:���+��_bP59��7u?M�q�D��G�Fp�0��L�j+!��@��`a�e'�l9I�l�O����]fꂥRi+��ܷcp�ټ�c��k�Iꁛ�(�52>���m��T��ޗi�)�<#�J���0�(v@��&%���V�� ��A!��,*�� �z��$ ��<�՝;�j�0�p��$w��5Ȟ4ī'�qL&��5T������04���uk�[K`z���r�����4��8��0mI7�^?�{k�<R-�@��9�Ԉ�CR��6v*��T�������_z< �7�╖A�Y`+aw������i۹j�G�0�T�}s˕R�\�^B�aE=��6���&|�����T�hzqgK���Py����L�U��7�&_I`AHVSpJ��O1t�Pv�j�˓�c���B�++mK�~gG{K�\��4�j�w�f)��{A���gtϘ7k^ƱH��M���r�$j��5�Ҡ�vv)A[�b�J
�V�f�M�����L/56��I������kISp��l��AaZm��3��z���g���K���:��"@bQ�,�¹��ƞ#N�0GW�\AD!�P�0�P	��f��b��J����j6�Ja:��~�8��ׂ�TB7�d����a�g9(�G�cb���N=շ2���^�b;��J�u���2�L=$���\��ɤ!�wݧ�"���S7��Y^%/I/��y��0$��GPd`b�ɛMS~j�`��Ӵ�$Jь���ʉ��RM;'�34t�*�h�D�zF�^��nZu�|�с�T7vM�p��F*E�Җ�Vؽ�f��+�^��VѦ����a�?���z-u?C~����l�^��L�FD�by۶$��~��N\}$U��S���i�������'>��C���c�{��nE���׾�w�^I��=a�PNB�*u:\�;P� _���mmm_��p�\���tӍ��Br�i��ɗ���^������q� Al��o���3�0��fqN��x��?��3>t�Ht��瞾��a�����;�SS3u�O���/���k�������=����YC��=���� h����+���o}��c��lo�i�:fJim���SxZd#IC�|?W�'	%��wu6�@����O?�X�%D&���Q��(N����o�@
�|�n�3�wzG�e��o�V�2����3�{^�ɨq@u�5�9�7ah/��Ҋ+���
��`�d��-j�i}�'�-	��@jA�M��}<�e)҃%No������^����:�D__߽��[��=MzY�v��o~�{��U!�E �6��KŎA�;�p��w��'�j�Rsr���}��߽�ۗ�29���K^��������>)�&(&6��_v�eo?�]���l��Z�)��^��\?V�̍<����x�qk5���Rb4_�����3��'3}�a�w<���/^<::*}rJ�
E䰎��/���m�R���R ��>����^6�S첉
pGq֬Y�Z@y|�3>y��ǶuwG��=�ܓNLq����ҽ
������Z}��+�֒��)U�+���%j=��F�pH����R#W?��ʈ���`��z{0ұ�	����%�Z�֭�6mx޼y�����θ��tw�)��ڦ3z.^�r��m;��
�MYF�r���;�HX��f$y�%�*���-��4}J�+�|;fspp���Ki�mb�a]�-23���x���N�U�[@��$&��=kމ'����Pt�'�&&&�$Y�~�PB�[�Z�/*Zf���R�304D�?�
��|N�$%�A˸v&cn���0"�u
�p

�@�̔!$�s�4'��Zm'����nVO��.v�y�h#KI1�Ϩ��F��{�u�2��UGC�J����muw�ٺ��B,[PW��0 �z���:>ٞ�Tɔ�Sݷ̓:�M���}�8�;��9�isg&i����$<"1�00vmx��1c�?�+˖-�3:��L��6�[s��J����8ٺ-��]y�gF�P퍌�8-YHE��Y8�~L��CC���K��Z�,�\.�Y�ԑ	�[��H"�q�&N��5<]bJ	PÙ�p�	�I�b�nA��Ғ���&���t<66&-���@�'0.��.����G�v�ھk����M�י;w.F*�@|��f�7�:q��Y�1�����-:���c�(�kVC��HEh�.x�S���ǵ� ��ǖq��~�p��1���&����}���^���@pA�&�KbY�Oc�!'+�CӪM�e<<f�~�U��g(|m�X���y�\����&JB:�4��|�`��Z�/'a�}�e蓱�C�vG����a�@�������>������Oc3rZ)KCpYL������oܸ�mo{ێ;ƆF�� T��Ξ=����w��}�c��-�S�ٷ�j:�r)ㄶv�6���z���ԝ2u˼�K�E�O���5�	ҙL6! wjJ�c"�TeR�F�(b�Q>��?�n5�G�fd��gg�i74�t\JDe]��(	 �}:��D5a��!�!��p|��]��Z���u�bM*��J]��(A���y�>S�lZ9�L���h�ph�:���2�Am\K�YN�-�(���v��F78EE76]0Z�K#�ҏT*?�jì�uRYlC�����~����>�'����,Y'HלY3��w���T�ݎko�[q�!NS_�dٚ5k�R�`�"��<(�Ǻ�|��[��w���B0񈴠�fds8���n��1�H]?�4��Ud�~`e��~�������o�����;/�4XI1Q�O?�����㣎:�C37Hu%�3�<��LfP��BQ�m[����_\s�5�e�V�ܪn��T��I��N�jEQai�}�ӯn��?�ahd���WM*�$3��Z�M���3fw}��W~��<��o�Xu)F�ʹg} N�O>��#_�{ĳ��7�u��?�N8��?o���4s�iXO=��w���CV��Of-f��|�W\��ث\�ë~��|�k_i�4:�m�Z��GJ��Kg����ɥ�0li�qj��;��F�ϊ�Y���F���7�^�a�8uU1��fDA���}��3{��SN?��[�{��'�s�yA��VVǩ�a5�c;k��FzJW��%���|�[��ԧ>��Ï�8�p��j�jeL�����l�#:T��U��+��d)���8�*C��8�ɏedL�Z宻�<���6o~-UN3mK�f��7U$w����ێa9f��8���dk�1l�ﻷ�w�E��w�����}�٦�sk[�Z�r��'6[�&��@��� ���3���t����o]y�ͷ��j�Q"L�)\n�4�v��1]�S�+5d�N�TC��F�N��%�u�PJ+�B�*1���B/��0��tpxd㖭�jͥnet�(���J��J[���/e[s�ho	"\����Hڪ��F�1�������|f��@ի�tt���,dN���pg��e��|k�k��)f�P��r��	�(�8�D��6Y�	�F;q�Q[xJ�W��9P蜘��ѩ0s4!AE�(H�F�m=N	���J��9ͬ�ttaԄ ��1��|��BP����Y3f
���9�DB�`������@6�������Gi��ڌT���4!�j�`�ҹn�;�.x�R	1�����M'n�q�G5�@�]-��Ȭ�����h����1[3�Gs�
�hu����m8�GǢ��" EK��o�ϕc#ѧņ^�x~kPv�Y.W��J�V��1b��wP�b�&�Nŏ�D��� H\]��m�OLJwTf���(9Sa�m��X8�-����bխR�Q�{��*�dbсݢ:�{4j V�Z&FE���`6��Ď�V�={�#W�޳����RuGv��FG����N8����nL0z�b��7�h��^��-���#�b��1�J-�A_2���F�z2��n�ӥ���Q�Q�Dc<�%�b9��'���Q�$A�!%|G����=j�֦���F�e|�X,���!V����0��}cI�B�#�3k�Z#mh��ps2 �ez�����o�54:9<<��΁a�2���s$���:�;\<�4+.�z>O��7x��%�f�G3神�D�x{�C(
B]�����#Ԫ��!�H��*�_����.���XP��|W���Ll�X�Pa��S�,�G9��-^y��&8��U3�xa�mur�����,n%��х��?�l�}<��PR���z��:b����'�A��t����ܽ*��,���dr�c����KQnH�b؄F ��j�y��B���s��­0uJ��&��W���6��S+J��p�����P�jXf�l�e�O���|0.�ƈ�hK�r������C�1�r��oéM�,�|�Tt�U�J�kւE�]]�F�'G��tՌT��B�$�iC�FAU\�F���퐕��ip�d:���(�����[|�����L�߸c^0��X����%�C�1�R����7�L(�C������zjF=g$����t_�>Q4���f�J��;�|��/R8��hnR:�(9FU�����6t�_������[o�����Hɱ�eR����O��ܼ�#~���::,fe���|����t�'�rʽ��z�u�}��Ǌ���s���/�� k)f�� ��uڱc�a�6^�|����(Y5{���W�p�����S��l�s�t`�%��f,�#e�5�AR��̓�mǛag�A�2��R8���9l�0�:j�Ci�����J����8����}�"�<IGJ��<7�a�� ����ϰ�qΔ���!�\}E��B�Q[�������w�mZ8_ �6ګk�B�=���V�Xq� ���vD".Xi���-W������C(i	�"8���3e20���
[/R�^�� �3��O��o~�����[˲���)(~z��r�	�W��я~�֙� bs?�Ȑ�L(���_�Cv��~I��dJ��v��f����>���Қ�)�Xq1�%M��r�$f�r�-�v�����8␘@���Rx3��������>w��W_�����o��vH�?�i� ��0�����}��믣�(�u�{ g۔��ԗ��B_&1E�5�Q�h�@d>wV��R!M(���8u��5�4T��0~�M�w��c�z�����;�������ZA�r��pL5Gܒn@|5M�h���4���%ȳ�����8%+1��L&,)�)�=�'�"!�B��^%.JQ$P�.]�a!)4ػ�u~���?ݾ���_���;o޼o��'�xⴶ�Lƪ��l.C4�E�Rf���g�҂eTj�	֎�1s�g`�^z��[E�.R	���!0Sb"�zR� f7w���]����m)��8{-�JA0	�>}�E]de��%ٛ���!`ܧ������;�ȏ�e�V�����85'&&`� wvv�͚���ցE�P�J+c=��.�Gǋ��fh��C9��z��ɒi#ڴ�i�8�i�IV#>�'�p����=,�X�������㒳A�ŹA=�)�*¤}ԋ�8Q�Ç5�ٓbvS����	h�q��gϞ�ϓp�JM��Q�� �T��S!�(6	v=s�m�9s��%��ZR��E�`�C����5ʜ�O�P����Vg����f��oowdDĲX����@�,]�t���v�<�{6be)��+�0��֭è���|�|����7�m��*����ރw��ܵm۶}�(Pm�>�9��P��e�9�$��a��-bb��X1vB�c�����)Ũ��"R��J53Z��^���ş7k�`1K6l�z��Ʀ�9���5H�'ׯ#>��v\td��+�����tN��j}���D�h�I| W�2-��U�|;��u;A6Q�Jp����7Z_���Z����C�z5�+A-���ط�6ĥ2��������}{!W��H��W���S��d�7�ਣ�j�n'��ԓd��.���W�Zխ&w�q����CC~G7ŋ�� ��)^j�0^P^�iRy��b{JO'��3�d�Ʌ��a��#-¥K"Z��r�,�$#��N�o�[���;::��߄c����� p��	�����ĥ���n2���[��m�\b�P���r�#��ı��O
*�8#�Ww� iLh�sTP &�w����W���)���nY�5�9������C�<��#�-[�S��عoϳ�>�d��}���)eQ�Z��g�d�Q�e��|�}Z/na�r�f͒�]�C;w�|��g��)^0��w��LU~\F��A�-� >0L���[X�}#�k�����5kp�K.�����F@��<�;�0f	���>�����bp�f8��I#q��M��r�����g>3<Y���տ�����E�-]r�������z�����`���*����q� w_DM)��[;�}M����έ޸��H���P4��4�u�������<蠥'�p���|C�c5`^P �49�}��"�ՑG�PӐ�p�֭����:KbDt��1N���vu��RyS��0��k���R�T*�P�K�X�v�~��n���kgLG�H~���ƢN����#���]�p���9.t�b�)D%kI�#�A��6x2���7��^�^M��43����V"lt�[����AE��'|�</��k~~���(n)��(���R/�
�#�λ�lkm��ګ�U?��}�s����z��͛7�v�S1�d��S�����3�5�E��3��z1��4��:�Jb!b��YaW��g `�Ejb衡Y:ug"^H��T��]�����wT�Ph��l��\�gd♟������T7S��& �z�ni
W�(��$�y�o�y���n�饼�X�㈊|(��X�����eQىnn޴�2!y�wW��U-ury��kTit�g`�ӟ�F���q��fö͛�$^}ڙD�隥�>ňM��ɓOx[wG�+/>G��0ܱ{XwZ�?�_��MF�QC���93q (�y|�ӑF���*�pmy�G��$'J@�����+(Ԣ����*A7�����!�Z�>����f�FU��{��g���|ͱ�<�tX)/����t8��)U �VH���nT)afXmϞ=���'��o>��TS`_S)��@IЊ�RW;b�ׄg(����I_�j ���A웸h��a\��9�\���^��~�	'���;R
�N�(�g�V�J�+���\sJ0�Z�չ���-��✥�~���'7l۸���U�+oRk/Պ1W��8�G���	hݒu4�V�f��z�n-�<��#G�ʨ��EŔ����؅Ub�2b�IV�ɛ�CW�M������,��I��p�>�b��b���kq� �k�E�#�o��Z�gah-]B� ��[6nٵ{ �8�;��(%:�b�>f*!�$�X���ɞ�ꫯ��[�SP�md��X�)&�UN5pdx�H7��т8��XG��R OS\�=q��)�ȗLj�Y�ԁm:����nY!�T+���%�F���D@f���6����SF1p�:��hBq����L�d�9C�� ��`���g��\G�u2�R%#A�Ԫ1I����Y�	469�w,�'�X��0�z�n��xLG���P���S���>�4��5w|��f�R۝L��g,���5�;|exh4��Lڧ�]�LF9U[4k&]P��8���tQ:�xkR���5�2��?���+�4�]m=]��87��2L�[�A0A��K�x�+X8<	�':f�RvSǰvl(<��`��A>�x����[J��Y6�m!R��v�j5��O���(���u���b��.B;*E;�ʃ]�mjRP��\�'o��J��>�>��D�j-'�BmÐ�s��� �ʮ�Z0,#�"W�Ro9��F��Rҩ26��s�F
�B���5+�$�[uӊL"f"1�TLs����ή֑J�����+&W=uGj�O*.�xhFF8z�[�a�S-�Z-�����6��'�1Zv#ݞ;{Q[Ilf3 �&����@�U�lF��e�*ޥ0�r��@�-�%ʔ�сG����d���p
�� /	5�Cj�6��
q-5�r}J��N6�`�T�jX��:�~�XP3�.����0��	Ć%f�
���ݧ��Zu�ԡ�T���;vTsVz.��I��/�%jD.c1�d��NL������ٸU�-�Q�Sd�K!w{�"�iR
�	����dvƴK�B���jY�{Wk�Lߦ�>�(���Ξ�(N���Z�m�1���rh�����!x��9ghbL�2]	���\k��u�Ju�@.��v��g�M4����3$jD'����q��j6�΍��o�9sfOG�C�d3&�zv2��=nΚ5ct���[v��M����h���6�͂(R�P34�\��5wxvKF�כo�gdԣM5�6mZ_Ww{��FUo��a�����b8��)vf�ŖPA�ӳ�T�r�� {����(�S5P��85!��W�kO�����^���3UeK�=��ʵ�tzPZ&f��o�喓�}&�S�RL���/~���\}�7�~�]��;�6�w�q�E����
XU����'Ϻ���z�����B!(X8c݋/�Q�b����s��ё���˯��ҋo�3K���|6����ͽF��l-G�ƥ��3�-�0�mC o����}�c���'��F�`Wp�H,j�y�M��F���*��1�#�[i��Y%;��͕F�*��yrM��wK��t-���nN{\O�W�;M��jr�T�|�ĒɊC�<t�=?����WE�T��
^�j&Z�+�e�y��o���+�>�Gɪ	1������ ����c���.� CՅ�Gr�#���Oc��2��%ۧQ�!��	U�@}��2�.�]�B�#��˷n�z뭷�x���͢�@h����iS��a ��y���<00p��8)&�
bS����*)k�c�1ݣ=���Nj�7A�/��³ϭ���;���l�S�r�y˗��'7l؀�
&{H�[�����v`X�b��I��@��9����9ܠȑ�G*�䊳�\�Tʷt��Z�#c�C6N�)�W�%h&����O{&&oG�L�	W�2��r�>��>���E4
��9�Y��5k���`����ܺ��g���f��.��5���r�Q�S�V
'�ݜ���E�����Ɯ���9<��#$Ȗ_���m��ID�@�:&��4S��B>!|��@�X,Ë.�h�C�Jf���3-�5o���+V`�ğK2`�{��Uh�{�A� �Y������>����;��K/s�1��z��O=��k���1�凯d�A4��'��%�	�|l�J�+��s�y���s�g>��.�W�\�o�F &�l�j��E�eU����Hm���j��?���2>I��H�	�ӗ�����6�x`�}sW�\���o߮X��R�����>`�Y�^�{��^��w|݋;��m(׵������ʏ=��f��V��`^�l������i#�DٵkW����nrE���n8<쫕]@0ǆ9-��|�:!����wIʫdj�S ��UҙDP#s������X�p!���ؒ��FÖkJ�$��9gN6#��lۅ�b~�X���>jL�KLJ�c�񶷷����1f�������q����(=�c�0�n��Q,���BE�}.��KĞܮ�����v+��h���I����0Nu����E�QiL���8���Z�CZg�^r��J��d���߿}G�h<����s�*��u|K�^�ˍ� [i$�dZ�B�C�H���*��)2Q�U+� 2*U�̹�Ύ8��+l&e�<V��o!x�iy����3#����s��(��w̞�������IY��!#J�Ș��F���C�i��J�#J��KS䇘�.�"l	��)I]1V~C�j�7������C_�w��Nbyo(���$�����9��(te��l���T7Q����R��� �nlf�N��b	0{�v�ܛ�L�]���тH`�-'K6�0=HѼ����-�[��n�	��TJ��Zi6����&~ڧ��'oN�J���P����#��do�oȀ�@��L*�4b�!�Cbn9��k$��rC�Kj�JY��E���1ρ�n��q2��IG����� �M�w��3D��Ք����P��n���)���h�z�7o��lh���;��ۇ-)�Ǻ��+������:��w��uSK	�2�����&�n�
�`]�4q�S�EҬw�u������2�q�<��͛�d��[�|���(�J����z>�ܺW7l۶mǎB��ԙ��'������x��K��þ��wl-a^��'{��}��pA�'jV���^��e����Ɠ�����!��w^�42��llNĊH�HZčQH�T���/nݫ�>��=�8p���O"�E�|�nݺ�·>��|��n;��S�kJ�_��W ��Ϸ�d��v'�x�S;n����V�D�,[�P��k�BP/��G��ӛX�#"�O$��c�A���?��|���$���}E������l��J��}�9��������.�?��;�_�^H}��8�@T���K/�Ч?���y���-9��d�Cߤ�,�׿����|����Y��"�ȅ��?��_��+H��(���\V��B)�J�O[��2	S���y��Z!6Ma�rس�ų�9�J����ÚQTj-e�J��3������a�a��L�F=^>{�t����z�K��Z�$fƤf7�� uLA�ꎞ&�޸m����U#%g�/̇�6�ɤ��}d|��r@9`���L�;��6TT��\EwS��� p�9hb��_�����K)�j8�^z��K���ZM�V�ب��V;Ca"���3�D�X~����ZՃ��8��T�pfF��EZ
1�ނ}E��tFR�8�NB(����M���Db��wE��uiKϔ$ܪlp4�������nqd�DP�5��{~dd�s�	c��d������|���w�����t+Nv�F諔�g�0o��ͧ�~z�����}��.�``0ŜQ�GI�A��!`B��]�S"5tfF�讯��_sFcҟ�W�������Pb9�>i�9:�:� C�(��Gd@�.jsts�SϏNVO{��~9Qt�����\�_�����No�Z�_�l�e�W��cO�[%Nl�&9e	bgl�j]�,�|��g�,r�j�mcI�8vgz�-F]Z�6W�h_x:�]��b!t�:��.� -��@*�u"���^Nx�u)ZR'G'����~V�*�*���_�:�8�5���,\����J��gO��6US�!�y'���p4��Vr�0,M�U����Z�[[��Z�GA\)U��4s���Õ�b^������nKKG����vQ�����HH�:5�Bfaf2!n;&��uK���ɾK��@�J����[s�5\>UF�tK16������_�,pL�p���=�� U��p�;��|K��q�= ���)�@%&*�̐$�vn��=Cۗ,<�dx�,4/r�J���&4�HI�LaW' ],�شi���$���M�w�];�����B'e���*��	��twҰ1ףc�{��gb���6�	�>�Y�P˗�c~偻��g�9�Cj>���v��΁~�������H�M�AutY8�RUi"�F^4!������r�
�zẼ4uU'Q,�tl)R�&�M�_�6[GG�t[������,��S�3y��pcc �X,�lc~���Ü�t��"�Y�*
{m#�jQ5�[;�BJ1�Tڸ�[7����|jEGP=c��]��E�Ӌ�F"j0Ma_��v�8��h��lƅ:�0�h�Op-%�#���"g<��Dz��?�h ��p�v`�������Az8
2���;:�V+]bu�����dL����,v/��2SO7m�X9�j��]�{7��V�Оiu�4᪑��L��S8&,$�L���WB%��Xa��;u�=�(%��D�O)jvD��Rʞ���PwR�0.��l#y�{Ϟ�9���s<�x0Y�&�h�V=��)샇m�D�]uk�Џ5���p���ѣ�&F+eӶ�x`��l&S�t��ήve���ݹ|���9�V��}B���A����mV�9�Rs�:��9 lU���I��'�*b���"�-���3J\0Eͱ����rm�]�;����t�[kvjOo˴��x�;[2�V�X�4��|��7}���{��7�??������\r�%K����p���*n1�'#e�y��֨Yz��"��L�A6�0	��Y�dG�R���_�j5ۢ�^���=��0{my�(�-l~쑱�qXM[�l�p&�L^�[� /VJU�=��_�ta�k	Ļ��2���W��9�a[vN� /���������;��ʦ�xf���X:�ue�9�.$i@����T NMYH�3��~vb݌���+����P�2���.�����3����_�7q�°	�!p�c[Ę�Ze�xł?>�x.oÚ^8w�S�fώᎃ�C�̳��u����o���,�3Y�g�d�����v��syGICj&d�=sgs��k�x"�U3��z�ԧgsw�w�jǾ�?����҄��A�����mڟ��a^}�Z2� ��:���+j=b�N5��Z�a��Gׯ�R��(�V�_���{%�OS�2���A���|!B,��~p�E]����^�:k��<?���l߶SI��+�VJdKa�1�0�4.]�hW��*�\������;d�f������ǵ���t���Q��ȗS+�e���$j��s�7���~�����4����Uj8���E@�zS���/�� �$�L���l�b$Y��^%��g���%��Tf������;Gp�i'� {�_�v�i��	T��ؖ�Gq��/��Q.�S�����Ѥ���(V�"�6��y���D[�n�$���_�g�gp�����p䑇[�5�����-oyK���'�B���_���s��4oA�Z&�����%V1�|��;�u��G�S�Z;[����u���:��C����x�����{_�7������]�����N8�d2�ȝ���H��@��$��SS�V���J��&|*u���k��c7�x���/ ��sF�/|�?���o|��}�I��Wo��Ƴ�>C�g��O��Χ@)���0�zj��ƙg�y�UWA��?��0��W�h���{7��(fXc�zU*���z�̪øF��F����#S_���4L�)1��rNW����.�4�Y�)7�P��`}N�>]�(ģ0���`�H{�̓P�`e)����?W*�������شi+=��c��&�b�P�
)ӊR����69�����#S���ʔà9?��zg�'���[qO
#?�$�[\���R(��!�`��39Ź4kdd6 6�ڵk��!w ��+���7��R�96B�� @�����̞=o����=x/�ҚXK���l�4�ϥ�Y��<��+�C��B)�I�\�R@0�����R��`@l�?F�Р<���|z����̮]� ��k�`P)�I��KZ���bpֳ:M���̫zN?�(�Rw5�T%���y�QPr܀z�kzC�%�C�E5܎F��\g3��ݻ!<�7o޻w������0�yΥ1n�V�{a&s�,�<1��q�zcerf���"yA*E~�8����۪6>���fj2�\�7�W����e#�5�3�NǊ�w*�]����j(�I"<RM�c����6{<I����!��l�%&:~�rD=�$dM���^58�/b�Ԣ[�?6���dXc�X�PO3ǊD簈QT'�T �^�� ��~k	�5cJ�T�ap�I��<�o��4HI��H8-5���>9=�vj#X��RM]$����}3��4J�%�"�����\>0 ���.\y�8��;���l����k�����ڠM�L�wp�"3Lm$V�r0,kǎC�q���>ʠ.���Mu�0��x֒E2u]]]P��Y�LqtR�R(H��VL>T��l�"\aþW(��k�d�J�"� ��0%�ڐ�:+��{��5��r��-��|���0��l[}��*%���d3yH]By���U��Y��Q��!7�8�tJCy0*�TՁ�jQؚ�5k��bkA�\?��!1�8�i���$�=�L�XohS#0oؚ����Q�_"	ΚZ�Eo&Y(ܶ[��^�BK�8��߯�; �{�����?�9�Ef.׿u�SO=u��c/������ 3��u ��ї���H��~��O>�䩧��8Yh��uo��@A�I� Ô$^/$�駟~����Γ;le��IY�XY�0�Z��_���3���W���"������/����ɹZ^¶g�u����b��FG��ؐ����Ws��� �Z�}W�����`�*�T��lC��.��t.�7���U���nc� E�w껃j��^8�5!�]�M�;IJ4�t�$�R �jʺ�6.Zrp&���?����e��E�/!r�����T��v�o�L��k���>�Z���(7Kh�����7��γ��8f�B&�P�_H�A�cD���l������{ѢE���믿��އ�D^f: @���۶o�osv&R#q���D�;��'���(����k֬��R�n�q,=���S��x~H���1�9b���Ǵ�2��R1�_�%��K���b�L-��X�J͈B!h�4͏B��m��+9���^U�9�ٗ^z�x����V}��.��i��;��
�ą�$%�0��a����5��Oo�	��F�0�DQ�V�+�� G���Т�$�8 %���Z�T�[t����c�>�(Lq�)���׷l����~�S��ᎎv�R�~(�����������I~����ں�a���;'�}���4X��\�G?��=g��eM��&I���̈b�`F�I�q�s�s��M�N���?�R��X�MU������
Gm�\H���B19V��m۾etd�o|	 8��.$EK�@IU��Tu�I�+p���PL�<<��K����D��8��N�|�����/<�R3�g������dղ�����u>�i͵�`-��2V.V�TJ�hkk�l�UK�㚥	b�ܷolw���靹���.P~ow�讽�n^?=�ł��߿k'vx�8ђ����G	�M�A&ׯ�xisXq6`�ٳ&�o�a�3J�'#][:ފŋ��w��Ԡ�
:;Y(
,��1#�¥|!.�-�k9i�2�w�����E�3;C��������>蠥�2��1�U{䳹$�vl�\��9zВ��j���Z.�	�X�'���X�!�']`nq����fω-2C��ke��g��S��e7,��rLw��qf̚N5��z���h봲���y�&�L{qI)f:2R4;Z�&��3�쳌��{0�X���>�&#���`T��f�U;}ƌ�A����(�NS5T�`�t��J?V�fb��I�T�����N�t�892:���/�|��r>mi�Rt�/�[[.�=��;7�|衇z�
 oq|�l���xŧ
1U��Y�&�rn�����Y�\�46,m�z����D��U�Q���m�M����Eu����^ʾ-���}���kr$S��ҕK��h��Ҹ��#Ն
)9>�Z��/[�iKeo��Y��נ}�aE��N�l��YҨ70!�-e
\/�i+����5��1�g�Où��ʎA��Q�����ہ��H�f�X-P�1��~�R
B�i��&D� H��5�Dι�6�{��B�� ���)��TM
i��_*�U�+�ĴLq���o>SpZl��{A7ꆉi��<ֽ���f���э�i�,��`��Å���{���M�(��B{lw�T��cj��1&�}��Z��ݱȏ�wrߞ�j�-�+��GX:y(b����v�DPC+����Y���a�A'$Q�V)��S�&���d�ǁ���s�}��R����û`�����{B�'"B��p�e��]��K��ϝ��v�<'�VL��=O�#l$?��Vkn�ሇ���%�i0��b&���l�r���Lh7�`�}�W<'ׁe�>�xT�Ԏޅ�v�(P�E칯��͒��9���|��Do�Pq�J贏�+7�t�g�C�7��Z���a��V�T�VZ	Ҵ%��cf>gd�s�HJ@K*j�
�[����2DM�pY?U�����TN9Iٽ�c��V�����RL�G�76��r�FDD�M	Y���]��{���s�$BT��n�w�d�}�	��,��Ρ�Ҹ{��U��z`�4�4��=w��KX��[�%N�c���T�*����O8�خ��[���9�O�9r���_�;>�/��;��w�e&�b3@�PU߿�{�����_�YU0�S�:�h)Ԅ �$h���j����_���Jܛ� 2�F�~����W�����߿q�׿�/aQJ���ʷ��'5�lKU��A�s�8k�[s��rNB�|�ײLH�m��L�&��(K�������e��e����7d�Be��҉Baf�J���+��
k�~dtl�+���׾F9��d����}q���(/Ȱi�s�S9*Rv�B;�6)6+���\�kԍ(8�������ȶ�U��P�� �e,���q���go=�ݗ^z��'�p�!u�q�?�����7_��e�1�k�~a��*��� ���w�Ka���s�����<��Yg��Z�0
% ��Ο?dddǎ�y����S*��z�]�wP�4}�-���6���Tc�`���Ԙ�S�w!���[J�;�_�ٗ����$�`��֭{��V�Z�0kr�@g98p�-���/���?>��G���r���	�R�F{�����%Ab\TG�)S(�bcS5WBc~�qq�r������Q����|˶���z�{｡�e�y@_b��$y�t r�u��+</2B!d�Mm� O�=��qt�?�
v��g��7��i��ұ��h�Zꛭ��Ǵ(��ppP�s-mc}G�y�H�S�À���s�p9��+���Y��t�I�
d�Y�Z����>�O�XQ0adr\Z�H��
��m&1��$RA��R�&%*!Kώ��	���K��|�֭�
9�k
�Z�4��������H@8S��j5@Gʜlx֩���|RE���X�T��໔��G��C�=H�(�K��K�8R"a\vHZ�hѮ]�Ȫ,S��n0���̙3��0!{������"?H�oђٜ����6y�q������f.#���+W�,�K��7�CᨚJ=�Z���O�l�2�^��J%� ���I<���I.G��;�x�qj��5�Y����0uZ�}��������%r�6��$�Ќ`4����aK�Y��zQ��b�NHɋ�vu"�D���Jib�V�[�4<9���Cq4m�4���O?��k�J	a;K����f"��0�2C���m���ŪԘ���j�QEF�^����7�����t��i�>�q���^�����٩�K��s}%�[��L6,dRb�4�;�2���J܉���A����L�LT���A{s��m�|��P!��3,;i��ѹ�Z�3m�]I�Q�c��I��Qf&9��$�Ys��,�S�J�I�a�Vf����t}�9�(i�Lm���"~2���)ش� 9���|�R��o�>����6�֢##!g��t�M���z��b3���H)Ou�89\���L&:������.��aΡ�0S#L�I��˓�rH����7<����A�K������E<�:�B�%�)K)���%��uX&q�1�#�uRq��N�@�Q@�V4�#>���[Tz�3��H�1I�d����7�e_I� �!-rv	ה��	��;�R�Re
�4��r9G-P+CJK@R�8���3��E��jzT�'_ꔺJ��^���qi����ϯ}$���q��~�X�T@�AaL	��wܖ������B����j���o��W�X1��_|�E��,����6	r:C<�>��?��O�v���<���ew��黮�gP"d�k��w�oO;m5nAg��ᙡ^;����_K���{�S����4N����U&)H��'J5�c�)L�}����}��я~��K.�����	��a���s��72�p8s�I���O�&����f6^F:���(��N8�֭E��RSNк`ŌD�c�=���R� ��'>�b�rڻ���]߅����Sf�t�'����'F?�ۊ��̈�"��E�p��_��fG~%K�#߯��LMM}�$���0KY�Z�2w4=�Ɖ�s��E�%HZ��t����W_����گ|��Ǣ��{�W|�����5�x�IǾ�Pn>HL�6mܺ��_�������?�w�D���v�m?���W}���W�<�r���;�������+������Q�����`��-i�+ۆI�?"nN*E�����Z(rH���- �!Ğ�����O�YK=�b������;��M�_����nh�t�_��{?��O>��#�;L��̹�}��ኩ�L}��O������������WRs�8j��k��l.�\��k��:-e�s��0P�t�;t� �h02#ϲ�'�eQ�$�xu���T�+���'��:��F��E�T�Pp��?��W]�mЧ}��P~��V�ػ��/��s��w�V��R3���j�ZI=3!2W	2��Te)~lf,��s��$���Q��(^9	S­����N;Lqa����W�����ٽ�����Q&f��X�T��MLe4�ڥ5��S���h�D����{ǆ��E&�@��v���*�L.��y�1��bk�m#�/�����=A,�|귶Q����n@��P[��C�L+�U� �Ϝ�>��GM�������C�a�&Qg{{�J�C���r�j- S�P�#�z=Q�&*�B����-�bTP�Y���Dܱ4Y.�+\��LC�#�7[Yԁ#e�K��e���f�h����~�{�n�Ӧ�vtt�8dV�X��Oq�`�;wv!��LN07��s�S��ܲi=��ji�7gv�ň+aì�)7����RP*Ol޲Qw�p�´^6�vkNv�\ym[?ݽU�p�3�`]ں;g��KtB�K�xͺu[�(��ق'6��i[Ki,_~���8������`5���X}Ǫ%@���X���%�֭3��=T�à��G@Z"kM�z�(��2��h)�8݈�ޘ����C]Ȳunݹi=Ƹl��0k�D9�F��6���x)'P��!�3��@M�v�84��l�niK9W���|H#�lHL�:� ��0��b��J���jԣF���m9�-�t�C�Q����,��H�� �G�	D����-��zO�W�V#)�iZfɉ}䈵�I� ��ML܉fͳ���@Yd�EV�t�Dٜ�?�T[Y����6�$�����_�T#(�%JJ�2)���1{��5Aa
~Y�
��XYx�!���}!�8����<Gl]B�X%��2W�$T���w7�"�\�����M�LN�i�M��M��I�Q��0�*)�J/TP�5?^om��-jiP��i��ic���^���W۾�g����n0�G��(����--���	<��`*Ј-P�QX�bWbovt����b��OL���C#�`���L�u# 45���0�����k���3�Y�Z�m˖�ysVM���p��x�Y�ζ��zzz6�߰�V[8w���-������3�y�}=��T'&�Ǳ`tU�º����tl�z����J%�1�_@���dC[����M���V��V��0lo%J�0%'2D�8?�9��S-Q�h���;�#�#�
1n[';ܧ 5֐�rș-�ר�1/4�@̛U�3�hϑz��E=�[�&�g@�8IJmb�����̠�׊8�1�@۟����)@�[��.i����7����.�jް(g��x+�s!���Kz��?�g��z�����7����l����C���Z��<�>������V�,�]���ر)6%���&661�%��¹g]H�V�$$��+��C0�����-7ɲ�ե��ߧ�}�����K��8$��0����_f��������{�����嬊]�܀�ߛ���K_�R����x���~�Q1C0��V��E1�_)�_u͵߹������w�:��|�o^���FGV����w� �M�$k�ԥ�x_��/����7��Vc�\�TU��Ղwj�����ɑ ��z\9��H�?���d�H��2�!ق ��GJ����}w}�[���o��vW�A���J_e��3�E��r�t �B�M�ttUݎ��������%3Qꚮ��Ȏ��S�ݙ�g�7���-�R#���o��u�}�]w=x�E��Mo"����nN���G�����;~���/�ʯ���9��|Y�8���ݱcGŻw���_�c��&�A`���_)2��n� T ݈ݟ�U�T���F7����}�{���/�c��k~��pٝY�_��W\q�+_{����o*�?�|����}���iu�?_�k��d?��o�p�-���>G�}��w�>@�������/~��/ݬL0Q��s�K7�CqQ�(&C�#���N.����7���f�Z��L^�p������훜���~�����F�`*1:r\~�����|�#�z׻JETx�u�:������o��o�ٝ_��G?z�����O���^o��d좒��4�n#���Ԍ%:�IU"�c0�#x�*�Z�������7�؀�cld��a�8��c�f�����#/,,|���ݱ�1���M��+���`�F{Ӎo����a����#�c�!�C9+�W���m۶�皃UͲ��H���Y�X5�ޣd���u�
K`[Pq��q�?�|��܍J7I��G���]vY��9rD�3���7{�}^�H[�� �\>��FGGWO��������+���!5j�G��%���z�U�V����Ar���"}sm��#nz[�Bt�!���EA.I������'�rT�00y����<C0��w7��j��m����c���c&V�Lt�6W�H�$9�L_߲e+�\ 7�۴�s�D��uzA�922Bsr���/<�e9ykdc�aB�G����� ���Y?[ ?�Ja�=L��<���t�V+�BT��+�lIY
Ut����G�"��Q�Z-������i��rO	�9�x���7�v�Eg\|��đ#��(HXv=tT��3�|��V�^M�:�:�eE�4��vT�`�q)��qQ��[�h������0O��IT��T�4W眹�NUe�����V�������L�<�����������܎W�@�ԧ	.������D3f86_�� %�	e	�;�Z)���m���Dj�I;��r�"_?��Rk?It	r]pt�O��3���E2��<(�'G쑚�J������IB &�1c#��Pe�Q�F��p�Z6��H�Q���׸�d騧x�D���/�G��i)
!�<z��$��d��㬸Tˊ��JWY�	��];9���lnsڕ0�JN��?I�5��$������'(`����H' �f�f�T�	8Pg6 ������3�F������w�^h�'L�N�j��t��2�$�I�,�f�ӳ{*�8Hw�`[�n��r����rM:�K�l$}-W�R�"9L��XH��b��/Ĳ������e:���\�U[*-�	#R龜��Nj,ѩ����E�"��������_Ae �8��ˣ�H�U$SC��%φ��
��1"9�Hճʉ�~��L�M9�k�_@.�r����������W��׃�E1�s��������{.�tZ	Ցm��{��|�{����>}��3Π	<t��@�� Q���f0�K�>z��_N��;������s�NR� �#�ۀ}D�4)��e�ڷ��-��Sh�[�Œ�%2� )
H�}��k����W
�V=iJ��Ϗ����E���K/�������7o\� =N?�t��������u��# 
��
��[�l!���3�%�.u�y��`X~q䇑&w�����N��&��}�o��57݌�:�qB����w�I��i���k�F���D��6���2��&-*�*Q� jC�j�RY-�!�t�|i3�0:A��=�S�r�12:�{�O��#Ͳm7�k0"�>R��B�h#2�M�GWt>S���_Pj��e�ѭ]����~��[o�§>|ٝwZv���K^�������/��w}�N),�b�������T4�g`O=�>���{��=����^|�%d�b�"�K������k���K^��5c�c�W�t�鿼o�b�!�Q��1� AG�&z_��Ŷ�X&��!��n�1|�[Yn��*�:�'C�Ï�ʛ��� x��ťr���mk�}����ܟ���w��Ps<-i�^U�.A�Cuz�Cŏ~���x�;>��?��׿��j�4V��`�����{QB���t��A�d��*G5���ZXrHh��w(���K�+�������N	��$���]���@j��v"��
~-!��1M�5���8'B�Sp
�,6nX��7��s����~�\z�I�#�^ئ�F��(Eˤ	��1I�/W�d9O����U׽)pJZ��u!�m )9����n��C��azň� �ZA�XQ��X�/ �Ch��U��͞�>_��-B�d#j�VD��=P�ꚗ������v?�ep������F��񹹟>��@�{�Z�i��I���|R ���E���fֱ^)�}��Ŷ�v_5���������u����[����]�믪�Z�c�N��ÑF>�k��c��
N�]�g^,�(l���`͍� �z! 5K6U��,�X�[�k�=�D���E��@�A_��qq��H��܂n�V}px�.Xh;D�E�X%�ŝ^\��-�TW�� �:�n�$d���trfz��vg�k���2��[X\n���㲫HO/��Z�Gߪ��A����g>C~�s���կ~5��:��n�S��>Z�Z<t�^�a��[���#�p�X_1Q6n۴�Ԭ�V\۳��i���4)�-�β�y5dm<zlbfzl-�&�X����d�A'�,�
:���n��\諶"��'{ ��E�����r�hl;ck�l9s��A�F7��� �+�Y����_�%��6��9��,�͍T�I>���Ѯ/�0��t��Z�|N�n�JkO��a�1�]�j �+Q�f�
K9w	��G�5�B�X 5��$Q �!����I:S+ ~Ӆbm��-a�7+�Dx2U5���V��8{Tt��O�5@6��^J`�2�`QCΤW�*��6�X)$z(l%(IKP��z%ARBK�M޵�HQ�vL��������bP�LK�&J��w5�A�1�kҹO=Hc%�~T�e�(/�h�(S%#� M�vӌܓ
�J�'q"4I���f���k���rlô��w�&y�8i���U�K��ߩ������X<�D�+�;���r%�Ş!��93šߡ�0JE�M��C(Y<��XD�[k6�������v���h�'|�%�\��dUO�w���B�M�=�+1��ãI�<��#�?��q�b���v?cv��'� �|ʲI���ľ�f֦�w?����m��d)j�P7n��I�*m�#�k��u�E�f=�w�
v!�^�u�A�k��!�Wt}��XG�f��x�m8n��	��|���qy 6Ҵ6b�ı��&r�~�q`[:�� M�Xth"��p�rlT=D��������#�,.&�$��&F�KډRѭ%x4��D��@]%I�'��ǂ�R20����+�WQ,L�!��q�7�p�x����hHwd�ѷ�}�� A^tK?�����>���(���_��6���� ��ʗ����]�j6��p�5�*'�����b�d�^���oY��������w���{ζ�����ӣ������
�J�Hi�Jrhf~����WW�ǂN4��hK�T%�a��"�#~�Es���l���2�<��-��&X�DR$ �4������Y���W�i�q��K1�;����Pb���$��h!o�ڡ]iG~�|�c���?�����إ������w����O�����g� �咭�3����c�g�w~gph��Դ+B\��;z��(�U���k	u �4Ab@3ؓu�
�,�]�~i�)��o��o�_��A�YƄt����V���1ڣ�6�0�����'�.���_��?��_�-2::�����\�����V�E�@���C�"���������_����x�����HN��o��g?�Y�a��M�����e��B"��潈�|��|衇^z���j�y����_p�}�Jd3p�mϕ`���;ix���#������t\��H Y`�c�*/$~��@zrr�{��$Ƞd�1������'?��~���zի���^J$�z�����Ї>t��w�+_��o!���m��e� o���v`�(�˞� �
ze��vD
�a����K%Dji��w�=��:��d�����Ѡ	�n�� _�����'?ٱc��g�-W�9)���_Ҝ��o��'��#�ݔm�0<F�I�Fnӏ)T���F�V�O<�����W�ZU����|�c��J�g�S�1��ϱh��J�,D;j�O�������4===>�O�?�����ȟ\b6���}�)�2��Lk�G�V���VU��2P`�TVq��>Fڄn���_a��
���\.1ByQAW��L�����SƂl�ܑa`���2���mZE`�z��Z-�MvZ-�#epp�O�x�ޒ�$"Kg�9�r݋����L��HVAI[B�/:����0�_x�k֬A�T�.�H�� ��L�U�V���/޽{�a���LC�co���n���"��C��i[RBFg��GD}�1�5����4$��UAnV2��Dؕ��h&�P��J@i:��
��uՁG}t��=�^6̦��0<i$1�<M/�M��߿_��k׮=r���Oc�9��n�:���er��ݐr"!����"�4����^��3,D2ЯzzzV��h�����'��'{��A��k.��� B��%��@+��Œc$ɰ�l[�����ZZ^�͂4���N�F.���}+�S�8,j1�,�X��B���F_E�p��8�-9�X�Dɧ+��ύCi���$�C�� g�DR�ޕ�F6�X�qԝs��.�*K`��5��f����|�+2Z�{Z�E>�Z4���s�)Z�ti�XۢVDֆ����'��)�F�W����Ƌy'�Ĥ��ge�Kut�2�n��<[e�ӄ��������%�\B�<x� �J\J�P*q��D	w�,���Y��ـ>RCS*���˚�8�&v-9�_�e�|Qż��d��0���Ǐ��`��C�K_�Rb������z������zaaN�L�����ꩧz�Uz����aUUjx��2���T�O���sV9[����>3��$=�luH[���O߶����<Cˣ�$�&L�����;t#,E��=�b䖜�U�\%��"kj�0l�>EM&�xr�����t��4r�4�4iϞ��H�bc�sV�,��u�'�d~�CZ�_�O�f�ů��nyGK��*YI��~d<�t=���7o��kiYY$*�k�s'�䪫����I�>������F2�����>���_�������K�� /�5"6�c9��i���y��GA��+KV�+D'���m���Ģ�Dڶ���,N��|�)�la�kF�D���2�8�_�3"��y����	cr4q޸�A.��9:EGY2��'��MC6c�$6l�馛>��ϐ����;�m��:I�����_��ib�����h0GZ����]�ő��k��Ok�3� (y��I�u���~�[�r�[�*v|��в�����؀e�o}�7�x��Z�q����q��8���w���_��}����?�ġ{{o����r�
z��8z�[��J1��-7����nfp��{�f�"��w��Q���Es3CP|����;r����h$�x�a��	0�K.�V!%Veϧ��J���ǎ�$]���*
W��~��?�h�U@���&�	��4B��y�E�[���ϴi��[�/ȜKIn��Y�6�]yы^����n���R��JG��|!Ӵzm����$H-��:A7����Y2%��r���C�e0mF�г3��[�rÍ7܄`j���5A��'-�)*�n�pÍ���vT�6xU��Ǳ�{��_�%�jy j��"]�l�a�r�K/Kbr��LbD/�V�g���V��GN<�`�M�_��o\���/ܱ1&���ԣ[ߤ�O0�$>�=?�OE��q
�7IX������_G��:������������ٙk�{��Ç'k�K�f�����%^�_��>����*��5��Ki�"���#�je��K����v͈�	���0:���~����i.h���ҙ��[Qk���T*s3㓳[��mټ��\g��v�ͥ	r��R&ǽG��y���!�Ѭ�gp��t|��h-Ly%�w��EI58�]t
H���m�D\|����|oJϹM�3y�S�\�8��Y����h�ss��{�hU*I24؋&��,*my��u�U��^E��qKz۪jT�{����G�cyt��!Z6Z�jz�w�Gf�g��t���v��,֦��kvz�.�j�ڍ7�>�r��>��N������07����Q����^.��h����噹�{l�V��Y���R��t�?�ǻ�b�P�1���Q�𐖔 ��U��e�0o��tS'��@&��'X�c�@HN�N���������V���S��m�gO(��N��Oy�&i�Y�r����\�3��P��T�z:y����{��P��J�{�?q&��N�bp�~ļ��~���5U�9i�)���؋]�@�lӲ��$S잕m	k	�[p�����+T��S�1)��mpa��WY�s]�2z��v��^�Z�j�z�צ8�9(b<�.�RX��Yj�P��� ��CaoG:&�	I%����f)7������\�`]%�Y������333I��X�A�GO��j���!mf̌{���wh;\z饃���5��Β��Tz��?P�B�f£�U�{{�,�������e$5�X 0��vO�h�q�&����g膝F�����s�5��h�5�����_=�ylyMK��oذ��4�<���$aլV{旖;�'F+�Z���G�u[��A�8<Y�ą��-֗����G�@�b h��0D��v��y��DJ�9�Ai�>$m�"a�4?�"w֭[;^�ۭz����ĭF�cx���W{Y$�n'3�t�>���F�6Q������J��F78�e����K]	K&⇭V�g������|���v�`=�������!2��6�Lm�<�D
���ǩ��'�Q4\�UA�!{F[�4�����<;o=���1}�L)rM�7��M��r���:W\�R�	�t?B �v���ƻ��=�2d��.)3�"���$e/���}�����Y���dĦ��[�x��C{p��������+�4EMr���P���T�j����~W�4�?�s󯉧�m�^͝.y!��E��dJ<EnJ,U/2�R����X�}�5��GqM.Y���n6��R�������w\ړ�aF 9�>�����}���:�  ��IDAT�w����pBt�{����@{���Ϥ��Ͽ����9}-Y��`&u��V�A<�~�Ѕ�y%�>}*�k�7���u�$S�y$;f�<���|ᲀ��h�R*�~��w�}����>�o�\D��>O/���a�L��0�`�e)0�Y�{�G��w:�BQ"�B<e<`*P��t��ҝ�R~2�-�V2j�ZK�.�r:�*'c���I\��'�1�f��ĲN�nm�r|�]F�H��
v���j-H��T�"�b�'��ʤ��,:e�_a��=�/����F�B;���'E��$ǥ��6��1�>�P���� �3b�������v��-��QO�.0S-ͼ�j7h��Y/ocױ�i.=�b�.�5Uh����ed5
5��Y۰���'�!����lq�+�H���G?������{ｗ�'7R�������4�%���'IWep��ݕ���qݐhY�������S�SSS놆Ɉ)�����'~򓟌�����/&_�| r��5^��\r	�~�K�X^^��;�r�Сm[�\y��#���&�~���O_���7��M��w����u���B�b#T����tOo��x���#6lh5�.s�?�50��s��BRA"i4������L�u�֝u��G�}ࡇ6m�t뭷r��6₪v����y�,Y�d��&����Fz��G�\��S0���,)�^�L9H/�%6o^{��s�>^M�,0F��9D�c�FKZ=I���M5}�~��X"M��Bv�e�������D��!환�K\s�5^xaR�~O_�y��ד�E�.^�ڵk�&-U*�&=>�.���C��.GO��.�S�{��E��J2sݹ����c����Bi��n��z���y�Z+���"�tV��b1�4C<��$�]ȻO���x$����i�$���la���nF(�I����$٦�=e�#M��U##�8z\e3<�ڲ�jz�V����kh���<6M�5�ztT#J���\�x�RZ6l��n6�� ��:���n"��0��eB�J4����_������4�&��d\k��g���g�yɆ�x幤gC�I'1M;N=�5��6�.�)��)i)7)T�@#��7�T+�h�r>����8�;,+>dVÜdf��9�����ݸMD�eK�)*�J%�+���oz_�+n	&̟4rȁ�Ρ}7>>NR���ϣ�X��DD���z	Y��z���<�kp %>%�$c�qJ�X!���%h�--���祣W:H��R:h�mݺ���v����n-��;."�Gch����]�Mz:c�G�PRi�Ŭ�)��l11v���8*�3.@B�g�5�U#�/���fm�v
m|���:�#����=��/ R�gOu���	�d��Ͷ'Ԁ����4�@҈��S*C���H3�ҵ�&�k:n�?W��_3B�G��:R��l�U����b�+$i�䔓w�?��`NNxq$�>���Y�x9I�r	f�ĩU�	7o�L����HQ�s3n��HE~�s�����8���0A�RQ�tEZW\qŏ~��3�<���ϗ͇̒���I�6����~ZaZZt�J��|�umC5�V�ܔ2��cy#�,i�$����u��HhN��isT�2y^KRg�Ve�d]	0iY_>~�x�HӶ�q&�{�=��y�����㎷����G��q����7�������L��iӄ�v�i�����jU��$wGOl���Ȏg�:YKS�j��JJMI_�ţ:ci�I
�]��%�f.F��A�4���L@�NJ��
�>á���q[�Ї��կ~�_����-4G�ɐT����y��R���l0vE�#��$� 09d:�I�C�I2�����J��tV��pa�n�B�{7�t_A|�u��Jc�t���b�����Ė	zMxHx�!G4�6�YB�}�Ua�`�-äp#N��ؙ@4����Q^ĵ�]M��R��'��{�v{*RhZ|�8dwY8?]��)8��Y�d����B��� ,�}Q�(��.�|��P�Sp
	cA"4��%��u����Q(��$����Ud*t���i��N|�"�^W��95Gw��_�µ׾����#���j�� �j��RXNI@��4N�W�$�a҆f
�Q%ˠ{�:�?���G6mx�K_:�g�G9|� �cH��MjAb�v��yl��={��xɋ_��W<��S �4:�c,�͓��s��r:� �zlj�v�E/�pt��Gx�|���ʁ<���`c�WYX�C�(Q�T�<w)*���#����O\|���/}i`�Bɮ�-�Nq�A��m8%�i�n�<�~�K7��c�����Gz{{W��y����~�<v���@u�,�[h����M����rm_'���UӉU�L����RE�!Z�&oƺ��j�
�d�� ��l��ٙf�}�y瑆����~}ú54%.oa2�v��u�%/"{��A�Iƀf�V�ӻ�Xe�E/zQ���ԭcSӳ��m|rni2/4� ?=A6����9�Loq��Xk/������^�˯%��<�����b��Y����Ҝ���N�S�Ɇh�{Lu�ٚ�,��<Uw��}��jɾ�A�RsT2.���'Tz���j��j���|�8L�����p�+`�3R��߉�SKE����wd�J�	"ߵ#��~�(�v���2;��:�_-�왕r_�|���Z}����L����=�493�踓S3^�)�F�Xl��IK�:��$��r1�$I�K�8��`.���ܫ̈́����g�+�05f��&��՚ດ�r�.=�������6�X�
�M$N,��"('�Ų�*�9�U�⺽Dj�Ȼ��ӻ��Z(�Gd��n�T�)�׎�v4�u� (��LB���C��%p�P*#�/�Z��iQ	�)�_�y��p��65�-��Ea��%:U	�>��6![_�v��!���[Z���j�*2+�'�X0
��`I曌�]O�n���z{���شi3�.�7��f]uc� �\L*?\n,���<��ȳ�d�t�]%�mp�ƈ�)E3bH��b�C�p�-�V��<i���cAۍvh������=W�}�)Zv���ǂC2�{{ZmdQd�$I��fӠ�1�Zm�n�D?���f?P$� S�,f��o�0�|�D"� %���� ��%�L����C�EGE~9,XN���W��K{��K/��oܴ��Х�<�0���?��0P͝dӺuO>y�4B�2@��v�(�K���c��'����)�=e{��$ƫ�"]7��iD��������iZ����{d����T��{�YR�V|T�F���(c�Wi�Km��D��=N�#\q�H�����Z��&�ѢQDidο�	MY�BH2�S,���V��m]���i�n���P��{*U:���(��N�#}&
n��r�NbOo|�����^���I������4�H�����u��]�
��0 �Q�b�$f�{j��\*�s�F���D�J+cF�ʨd��Y��~d�⍻ �9�0���Pq�$��T��L�O}�ӟ��'i�~�v:�޾>4PR՛n}�~�6�4�z������It���~Ȅh��k�y��� ���W�Ge"���/9���P<y~��B���%�M�b���0�]W?�I����ƴ�Vk�8��"#�g^�!qK`�J���k����[of�%f�9;R�V�ڰ� ��ddJ
�i��#�=��Ba\��u��	J�iR���@7V
*��jhx!xi}�+d�EI��:�Y<5'�dn��Ce_E����-��9"1�S%+�Q�	I�\���V1��Zِ�r�0B�)
��g �N,�1�p���r��e��*��(�f�A>�*S�{���`'Q> ��ȿM4.�V�W
޸��H{!���Ai<�����TU~
I��g��.J���?���Ǐ���A<�L���g}���R��w��R�@S�)y-Y{*34�ӯ�"mqlq�ta'
�=�0@cn�Q�G�~�mx�����s��8�U���	:9HBD����ؘvsǎW_}5��ۿ�۽{�FKM�D��˸���|�q����cǎ�%���_����wnn�w���oۭ#�hiʖ-[H�����A!�;r��W��2)�����.��W_�>��IS���/W���,�i�q��4��-�[�5$3=�)�얒1p@V�d8]X��&]�����.#Ou�����Wl�F�1���'� �{�E�۷oiql�Q<33c����@MhK�U�xZ�O�
<DOimlݺ�x���ool�0��+_B6�GvB/Յ�Ɖ������C���u�]�m����Ez^��?h�W�T跭Z���qI��9���y@3��!��p���ޞ��'Q��T��U(�I|-�;��G����`�"�賋��9���ڙE�l@�Y��2D��a,l�]�>�ɹ[����Oϱ	ا���C��kPe:�&GZ��<0�,�ršv%a�dW��bfV������e��]������+�:Y*\z	�Q����?�^>)ښo^��Ԯ��"�C6R�$ʄ?rmg�F�9��/�\�lz�\g�}�V1i��U����g?�Y})�~o�6rh��6� ii[mذA�!��Dg�0g3�0[RU��$�I��pn�徫p���q�_��]67'g�����'S�Gq�Mr[�FB�=��6=m=^��ѩ��=gTR�V$�mb��(���cG!c�
�N��~�1JƘ.Z[\���\1��c|����S�Q��5Z�T�<��ei�˨�c����&B�]Z����êDe��M�l�v�x_���d����Q*K�CR��V,���3�#N��Okc���iz4�ǟx]�Ⱥ+�3�8��s.j��4E��ɩ��������^F�rߛ����k֬9��s^�׌���]�WeڦM�h�$�L��}��S׬��88X껠�F����֥���ũG��{����P㦩�A�̿�����zW��n�&���PdQq��9p��\K�TMekͲ:.j�i���M��B~�k�n��Ʒ�|]7���Uz���.<:�(�ꪫ���bD?(�	�����2�V+r�F4S���{�8N(1H�}�\�:�({J*��N>?s��=�D"�\���%�e�]�u�,$�'fAjڂܖ���Ĉ�"*�J�l)R����J��)����-c �G�]	�����TN1�~q�t<����9���5�Q�)Z�ہG�����O�~ZY��Y��ScԼ��O'a4.�("���-�d�
'�/��rL0�9^K^M���uTt�CȰ�]-%�<m����[��b@��ő�$����+l�'�V�F2x���zk(���@6�而�eQV�x�*�̡8[�����]'_JH��!+�0��u��f�᳧�@�]��y��mYif����h����l�h	�P3t�91��H*ɣ4h@H��@���X��dxT%�a�<?8-Ӊ���8�
H�0p6P�6&JURo��2�t7��j*����X�􉺒r C*'�ڑ����C�Z��,���Y9o���7�z����i�HM^x_snx�0 c��R>��-�R҂m��b���`�0���G�L��$�e��v��m���ԡ'}C��]zɚ���]c�T#�����ضn�Ʃ�i�dZd��v�Xk4g�וֵ#�tz{h5>y`����ھ��۬Ͷ�Z�^k��]�T��t5�l�3/��;E��[��U{]����{�K��;z�lD2��[֔׬Vz+3�:9��ޞ��9ur�T(���F{a�F�w����/.w</���� !N��^2&V�#[S��q��/%�_�iy�fbq��a?��]k����X*�qq�3_���ٵ6m<��MVd�O�ӡCGi�7o޼j�0-+�4���nih�K��m�S-�W���ov�N5z����?���£�K�6;;�����3�����a�Ut��C���:6I�}����P�|��?�u`U�KM��o�O ���㢰�7��-1Z'�;t:�n���U�ԚZ�r�S}�RO�**�W���� \�r�Y�ܱ�Xs�n��f��� ��F�dIC?%ˬ���eIv��r�b�r l��*V���~�9��\���A��V�k�pðL7�ѻ�k�`�)H��T �Sdd�0�C]h�W�0R�I�r�����hqCnK�y��k��{{���+�`���E�$�>�������d&%�1�l��.�h�fVK�/�}�I�̘d� �1*�ℵ��8��%��]6ioƬ(9y��>�anڸ�8���ۻ������Y�Z!D���p�,���������Y����y������@��"�(̨�E����0I�R.;�`v��h`I�)}rjH�֠��d��7V*=�+������I�\�SN�PiB[���+vю �\� 7�B���f�6ZOuQ$٭�\GGN�c:�΃��uУ���Y,��t��=�bE+�N��ǐ\M�:�a
�;yt�Jղ#G�[FGn��n�2ɺ0�G��� �ǲ��{�]�dr�n�3I`��~��f[�1.�Ӵ�dM���z�q�<��hj��������իW���(�������y�G���M׿���%�`�Q�`8�zm��tG}�P�+_�c㺑�g���/?F˦�Z�t�yn�����{w�<m�Y����^}�С���������K-�H#Ta��°����=��L����C9я������Ȑ��6�]�����w;�iKU��ӗ�.�	
�#�)�P?>'��8Mwq-t�M���gN9�tZ��r�n2�Tv
��0\�	��"�jVC7�� �n�H���VbctW�(�8Eh�[/���,vNw :��s�� s>R��q�@j�_�#nr��??�^�H'��HVC�T.%��aԑ0J:�Ƅ�G�[A��$׵��4�FZ#��2��p;�f)��IH �b��r�iՓ��\���9m��pR`Rd��)x<�0e��=�5��"Q���g�aj-0iiw�Z��D(����*�ň�=I�R.�����&�Y��)G�e�$�*w!8`��Q�@��!���{) Y�d$D�a!���=���S��l)H��rޗ�t��	>>I��|�����H�s(pvwJw�w���In�y��S�ܽ��#%2!�9㬲��H7�3�V�5��!@I��������LIJ�+s�e�q��)RDf	YS.���8a�M�'���1x)XH�U�
H�����4�8�t��j����*9c&���>D�H��	��?ydN�b#�{j\G��U7uq��00���1);<�	�X.�a!�>�ͫV&&&�}��W	5ȑ#G��]�i���"-��0]kO�'�[.����ؐ^t�B�P'Ŋ4*�.y_�vC�r m9�+_&+�AZG$JB�
��$�)iA��Ҋ�~H+�,�(+�ԺH�d6��Q�#W�È����ԑ�;����kk֬�����Kf�b�jEF� ���m�����۳���^�]�s({X�~���9�^{-٣2�6�wxx��{�D'���v���Pbµy��!�����M+�����y!��Z�V1ˑ�I�n�*� �\�������K��.n�\��
�CBI&��G�#�� �f�1��ue�JuJ̝�H$�t�K�_De��[b1�!��!B!�����A����-��.6BD��.���J�����)4�iI�K�o����,{|JM�MIZ9y��2��v?��r�I^�����^^5s��s�d���I�XW2���E��| ��5��|w\/q�<
Κ�T���o6�ݷ�MD��uYҿ��@{'�|S���sV潧,,��Ӳ$_+PG�{HrҺ�իZ�5*��t��_�m�u����w�R�U�$�%I���4�/-4!�hu\ڡ(�dN6�*�%��	����(�JmL��`�D)e�Kf�����U�b�ڙ~�d���8^i ���jE��S��u!�m��rq��i�'' �m�ޤ��󌏏ө�%C��F�-��pt��cܱD��իPJ�c߾}B��9g˖-ˍe�ߎ?NcX�f#I��@�80�n"^��1�d�&M多�I��s)Bag�cZ武�86�3F!��(�h�I��&/d�|�d\ĕ�"�A�V,; ��x�,�U}��VԔ�OLi�R���zr0�H����e��2Β�ӒF[�$���7��Ż�y�4�w1%iU��ܩ�J5㚖�[.7�ZA�zbR��J�/+���e�RƢ��-�L��Ŝs\vr�a�\��\)0B�b���?��$L������-�|�䂨{T�p�N:��z��-%=���iW�[^�|)|H�%V�F���e0��7�ƣARM�\�r�֭Bd0�x
��K�G�?~�y~�����0�9�+={�HW_6-�e�48���{��J�=fa��y�2Ne�d+�GKK��u�6f�bR�C��pwq>5����
t�<M?�+/[���o9?s��%�1���L�,�L�������uOW>�٤�HQ���]�uL�:Ũ����|]u�����{O�LP�1?���Y;��GU3��B6���� R�g�>������U�G�� P�����=����N�h�E4R��\(F�g�f}�67�055��8��k׭]��ء����FF֭[���|�������AȣA��8�xH�vnr�t�H��cǢ $��S���~�U�j�}O����^���=a�YG�M<��d&��Vԍ�U^?�
K��d\_x�b٘?2Ѭ�s���&���Z(_Xj�F⋃Q*�5�&&��#5��=)D�,<�\L��ܱHu�� �B6�b�6�L�
X�\�C7I����K/�~��g�==9I�(b(�P����<�m��uփ��Z64{�m����A��{7lZ�u��k^���;wn\�k�Pn}�mK�_��W����5�y=���rr��s�#����/#?���#�F+Y�O����CCC�w�ݳg��}6=^K?:?s�駝{�y4�����P�ψ;�ņ$
��1�w����Q����M�g��0ҹ\%���m��d�D�,e���ة*�h�a=�D��tHg'H"*j���N
�`j�طЕ'T��f�Z��׿	^%�c�?t�d۫K����=��Ը�b'�S�m3C,\%2�Rj3U}�>��j�,��*6�"���p;n,6j��KÃ��ˍc��f�/��ΐ%��ܧ�N��%����}9�Wo-�2@���a�
c4T���ra:K5�L]UNȩ��v�T%ۉ�z\������z�5:Q�#�ç�X��U��:��r�ξ:bsssB�3�]��S�+t=�	�����R}A�m�x(���DJ	��m�'B<l��-A��a�F�&��P��2��.4��o���f���K"��_��=P�N+I��J�o����&��b�OB7�h�'~o���6!��!�N�rt��J":R���v,Z��&� ��a�+�+t�&�S�T���V�
N����I>O�C.b�`@�֧D�c��ԡ�J�㫆��K��hY����/:���	`�Ҥ'[�m$�`�V���F��r���z�{׭j�[�����}����޽{�������W\~���O�O֬Ys�U�&�ia�'U�fZ�V�6<<\��7�Yvl?o��w����g�u����O�ޕ���}��-��8묇�z��уt�t-�Z&�zt�=l��峞rXI�J�9
L�D�����m�и)�"��q�t2xN�,��ΩEG�%w��*+�Hj�@z5=f�0��K�|Ӥ_.�!�735�����7O������rɐcneL�H�8�S�*�	�:�$�/ҋ'D��GΥe��j��:�ɑbh�r	%��]��JE��{�d�Y厒t�X��B�9�W����(e����O�꤬Ju+M��{�]rL�^ L�+	�R͂����[��Z�2i$�0<=-{QR:����2&6������b��P������P��}�Ms��Y?Ϳ��^-s0n�PR@(�Г>�n<�X$�Q6�k�B�)�D�JEd(��D���466�cǎA>P���3�}�٠�[���VV@��^\�<�°(���I���N���t����dyQ�3�	��v��
��Ss*7ՑR�ɣ������@�ZF�-��en���MɈ�0��'��?
�<M�@,Q�X+4�*{{{�\333�!�@`����sk�t������d�
���/����gu~~/�]�O�B>����Çaґ�ת��ll���\�N~W��F?�cmAAݡG�o�3�Ư��w�l� ���3�"X��$FE0�ͩ�P� 3�
)�<�f���
*{�Hט���1�y̫��[�Xl��i\��#�JsB�r�j?�B�eJ��5ϴgVT�Q&�zCAS�g��cd��<őd8g�;M/�d�SO�i�-MJ_bf��t4agǐ)���b�;RVvb�ƞ;Rҧ���_��f�
)+��M��3�^��R+��6R�{N�1i.�ġR��L �b�Эћ��g�d�OZ���d�S�
���5�I�ѐT�a���Hɒ���?�|ޔ,��.zM�D�D�_n��>r���vș����#�� ^��Z�HF.��zT:_k+MҲu���$�$���'y�$�S*����J��U�x�b�A��i�I?�-)�G�wyq
 �+'d�'�;{e��ԧ����$Q��� ��<b���ݻ��~��R�Q������J��)�t��D֤�C蜜��Pc�֯_O���䤰({-�-X�䨓�e˖����
ة0��!���mH��z�$jכ�&��k�1y�G�����J��d��TUj�l:5��ɳ���h0F�*����1b�a0v���y�kQF;����+���g�Pxy7�ijNS�;�t���g$+��&�!q�I�FǠ8l�"�g �)JW��H/�Q]��OsE|���<���Ţ�bՄA$T� ��ȋZ\�i���{�Y"�$;H~�1�Vg���U�Es�S0�c�t������|�=���~y���Iǿ��ՕBU��ͳ���Ty�,������fD�9>}����r����q�ٱ��{��`,ӣk-I=X�7�����$"�2�(����$��j�%9���I�!ҝ�b�됔-蠠L+6Qn�n��:��_Tm�.u��rӭ��P��-�����ݻ��.�uۻI������x���\q�o����=7���]�i4�/�5=�t+}���D�gWՋ/�^�<B�F��g�M/��l={����e�z3�,/��x�3��>��3���d�v���=�v>������\��v���69i���O����u���J�Q�L��d���v}�B5#�7E
�B����l5�g�C�v�Lj������u��LOO?���\�n�:�h��NV�s��SSM�C�Q�P&�G�K�E�B�jy��}��:z`���n�1<�w�������y�-�{���:����{��  [��7�ߎ=���A[)�m&���*���m�766:��=��%��!��/����`(H����[׹Vɲ}�|`8Hh�*b��u��hj��z���-&5%��J�
��;�7T&5fǦyz;
=@p-fG	-zB�ժ
U�u�����7����< ����I����%z�42�
tMJ�ٗs�x����c�ɴD��%��T"����D�~W�It2�#?lu��Ҫ8��sn�����8�����5*�M�6;p�,�(݌Q>�@e��kʉ�ZJ���'�k2����������1��su�E}N�U����c��Eܝ���B������mꎟ��ʕ^U3;-��w�y�Y������T��^=&�&�gt�v�,c�x;!���GEW_���)2�
��J�T.� �h�
N�A�/i+䳷�x(�u��x�9s�'L��1I���q���;��{��09�u���̘DK��-���`h�P�����
��O3K=���Rڛ���^ �՘���oM���u�F��PM�nW'�a!�d:v��j/.?~�)Ӳ-,4���z@*A��HI%��u�E*Y�/a��y���:=;9���H=-%Z=A��j��
R�0� -0��s��cC
gVK@��Y����F�f��<77w�Kvlذ��X��<�ԓ�%J���S��B�lyq����y��^zѮ]���y�^Ϙ�0�5�l��f�B4�Г���rΙ����{v��^F����(��j�ǎL��<��^u�9g�����tyy�n��=�(�]<8��R(�t$�w��LM)!�bEG�5��@s��3���pE&�N��T]�GQ��ͮ��2
T��y��JH0kL���,]��.h�`���Ѥ�8
�'K����!=��n'��S�q�`%�ZSa�JO�ɜu)�T�S\�EYy`q�8����$Ir�A�ܘ�� S�@��2�Y>_�pUⳡ�0Ѥb6��
":P�I0_@��g�bZj��V�,h���[���� DN�\��tp�q�e:�4��,���?��M7�����O��}��a쳜�?��?�-��yWҿ�C}V���y?�+��>[���l�4�Kj-��1:A��~Q��_eĶ�<%Ç44%�2k����:i�r�J礏����(��,�6ȯػw缾Q�e�?x���i�P�{��A�����l5��V.�{���Z�47]��t������j����رctN	\	`)�̘��З�gk!��-��k����R�+D�r/"���BV*jEh�[Zj����JMr2B�T���w$S�j���
���[���.J���i^�;p8�#Ghn�Êc�1z%Wt���l�Ԩ��$S~aa��C����G�.hpk>�M�좑���w��XG��yDSғ�/V`q�mh=�X39���/���g�-=�}�uQr`j����ʈ�OZ{i�^�$� >�:7�HR�
C�TP�? �	V�Ά����5xY��]CV�yLl�ХQoCڄZ�4��� ���ʱ�ݑ?eٮ�M�M���7000?	Ñ����ܐ�ב����)�.�󓀳)�)����]H2���gWvzҝ�>�e��8������@��Vg*nA�*[aKvJ��09�-5$�?��M�td@79}��Ag�}�dj���,��eG��f)ԔD��A���H�n�r~���_>���"�����'���8^N_����ׇȳ�U�%9�������F�2<488hq���i�[������{I�d��J/W�����%0�w��a��
0Ұ1TY��>���
�g�}*M���RM.�w�U�N���5/���D_��y�g;N�h�L���U��U:3� +|q�+�@�F�R�@�#�m䡝v��'$961��^�eɈfQU�bf�{'�.u@�cY�������Z���Z�f�&���餫I@��ʶs�<�n��5%#��9��ӏu�J.:�,i�H��ee?�Y�(2]Ռ�,�#�iD����x���[J�Gn��\��a��-����I26a
u���B@���Rv%ն�4�2�'B���]r׹�����M���䱓�T}6ƿ|���E�cc�s��$�l�J&��h�ZR���i9��Ŗ��JӚ1V#�q�0�p�A��Ke�|xS]�A�(�Y�%A�(\&]aU(1��r��s/���W�x�?������Ψ<�w�E��B�ҝ�y������<���{��^q��SG���{�O}�I��t�Ϙ̩��|a�����j� ���r]QX�1�~!^+�����3[���3��P��(Հ�ĭ�����Y�>���,%�:�ی�F؞�����}���.�'v�*�	��x㮻�i0�`h������51{�O��4�^�n��l�Ş���a|���v�����B��n��Tڷoެ��N*�� �־�{��z�N�4�����~��4��f�4&?�?��i��6U����[����{L:ei�u�-`���:T�9/��ЇS�t/P�0�N����/]��?�����R���j@�L�>)W����I�p�4����F�F�/�JW���ͯ�ڭrO��nq�F�iKG�1۶m���#�˴�j���a/�s�����?�/�G.>�����|��\3:F�>v�w�*L�_��O�6Z������h��a�sw��I���H>�0�gap�4n'���c�O�t,J@���~P����/��
���8q�\s2�.l\C3�Ml�?F�)
�H��j�k�M�0@�����h��O`��e��pl+69��x�������ꁏ�a�b�J%����]f%��D��]MI��z����$#�wL+1�ɕ�
g��,�x5���d��Q˚�x�J^�8G��~4���G;g��͛��?:1�/_{Ζ��B0��_n�M���UA-�*:F$���Le��pR	Ak�ъ��s���}��2�n��)�&&�*YEZ��,|2e$���A-J�2+�~Mm�:��2G�f'\�o��c�M:��r؞���;�����[�n}��'E̴ZM,�_�f���$�va��8a٥��k�I���N-qJT�K�BJG�!�}�v���j�O9�"K���D�G ��A�
}}tt��+���#C����`�@��f�������<�jt쬳���,�7m�4�ູV� ����dc��mԔ?�y��ӤZ�!�v��@�aO��`�0�gg���:�Ѷ����Nk/�.Z6=P�@6��:�������H��P�љI�u�znRQ�_)/�T����ޠI�M�W�$��K:�5���Bccc��voGF��y��ڒ�w�={��jd����n5{K%]5⠹�����t�B#�{��F�6::�[�]�v�,�7���݄�SSS���/.ý`:iw��痋�
f�{����[[*��)�cG���I�����dO@O�����)�N�t���9	�r�z�>��S�5��QS5��EQ��:!�G���p8���MKC���H����䈝� ���~���3B����j&�d�O���<���5���j�����NJ&�6��o'�������eɑ�3w}��Wȕ�]C�0s�o��^�T a~Z� ƚ��y	�r`�Qw�$]\����@v)Ŭ��t�=���s��J�-�A)�89Z��LxA�c�m�8�;;��WMi�)A�Ē��"��o�ZϏ�W�S�{,'������oy�����o8��)���}�+j�=u囊�ri�
�{�4N�Q*����;�Tt&Z�

��G��ХQ�䳑ǆc��sa�=�O
��],p���n��4�k����9��X(�'�l||��)/..ڕ*��P�v`H@�}i��S��z)*��l߾������Yf���0�8t���'v�*N���%M�/#E;H2$��I��6��X�v-�S�@m:77C�i>Y��3�8��/�.�L��4S�ݭ_�~ffFt^__I��lxxɺB��f�!�%�F��^�������N����.a	ǹ;!���)���f>���7N���)�hSȢ0��C��s�9iP�
@_W�*�?�|��v�M�� �h)9�ʝ�`d�մ��ג$@�B�o�4��A_��%ޑ(oSc&�(�-�]W�b�V�Tr�ڳ\J"�+�`e+�������=�i]��626�e˖�Ud�6�k�ȝN$Us����q#'�6��0��H�P�����;���Ġ�HL=��:�~Ӕ�G��@��]Xp�hrrҮ/OMM���̪+U[)n �=!8-#��fe6$�$�xGZƚ+{D��I�T%cJ�b�i�Ͷ<��{6��J=���}�%�����*�kf�jؾ��k2�CbY4N�D �<##�|��
N����-k�c�C�"V���T�Ѿ�qJ	W�?�Mj�J�V��H%+#!�MFN�ɍ7�%��s��'�ȍf��U�.`���`Cڄ.'�ŧK�l�@��ʐԙ��������m���=�s�ґ�! �A�FQS4�Db��1ɗd2cf��D���D��(�b��T/�v�m����ޫ�y�Z��{�(�o�Q��r8g�U����}��/w�P@1�n�#Ё�I�K%F1�����	''��,rЈi%�H0ܨ�BK΄�R2P���N��o['np'oy��q����'f{(ˊl>��igtL�=a�1#T�� 3��Y����婪�q"$=ku7��1��eOVy�Ԋ�y�$�F�p\T8پꭕ:��g&.n9N���z�3;�Խ�|�8=`w�u� ��Ȑ(=D8+�R��v'���8ɼ�$��Yq{��������
Ll���i�׆���E�M�f�{�b������/���l��ɟ������>^�����'93��׏U-t�#N�ǂ���~~sZ/���֋�!��8�����	zRZ=�bm�(Nq��w���O�T��>E����!��IU]��<�f�u���5U�C��dxB�2Rρ�YCn�R�?��D�|}�-9�5CsC�^#/Pw����m��NXc�H�Z1+9��]|ayi�Ν�����
۷o�U��s�U��kE�i���a�-�c5��y��&8�g��u[&N;}���Ա�e�3��w^p����w����ĝv�T*��B�!��,Ș娚�f���#��j�
�a�:܄<��z�F� a�Y�/&(��r��v������ٽ�CCy+�YF�÷��P.�}:��3\)�[QX)�n+�=���╗{���u\�<덕��b�F|ż�3s�R*�m�����`��߯��́��(��H����*
D��R�0�H�_3h�%K��*:��I譍DbCL01MT�m[U�,OA�Z41`�I��H��D�嚆�+T�
!س&�g	\�H� ]�_QQ5`u�S(�w�	PdU�0F�Ț��Q2q�*b@8~��؊(<��}a(�j\��^DD���`�IL*ѱ��`�F;�����\-��jn�КB�F��g���BkTsrrҭ6�z�{T4c=�Ԩ1(B��W5<�G�Jt�2+�K�R�g��9�SXְ"_��t�%�Ռ��n{qdԶ�6��Z˃��*X_T()Φv}ף�?���8����9?�=&B��&�bF_�v�Q�q��ƣ��0w�(?NJb��="V�2`	���z̼��&��K��^{-��9�	/���o//�}�a��	���`���Cՙ[^��	G6�S�0`ۛ]^���I\^25b�̅RMgK��,GЀ��U�)*�[�4�m4iE7�1U��#���g���]��Т�fn��UުՖI��LsV�r��h�h��V�X��zle	��x4V���̈���hv��!FW�Z�0X�FA��PT���ptِ�N${mM�[�c�M���r9�R)��[i.t���u`lAVR��>88�+�˷�[�X��J�H�N�۴i��,�u��aK�n7������kТ�,Qb�B0�(�08",�ȯ%ѿ���á+��'1.^����i�.���⢬��5Bl����!)���7���5A<��k�Atɚ�3�,�aF?u��|��'�&��%���ޤ�7�X%=b "!�r�y�F�2�H�g�
Ffj�=)��t�)�"�	d����'�MN�Uz{�O`��8�W��	�.� {!�^@H,B>gy�hU�v�	4�y���1z�����*�LS�z�F�1\\�+WN�d���!��)X��#�*�g��?����ޟ�	�����?���|����>Y�3�������e�rBrc+���n(��G%U��T�}�"�cD1�b��כSSSm��Lʷ���ji,�1tX8�g����GJ�.d%�k��0h�g�q���R=|�p�X���{-�,��F 
���R8k����g,DNԾ�K�4�&5�raP��;���S333�G�F����~�I�����s�
�w%t!��je�ް0=���hp�U��:��Dп�E2��x������
���4|H�eZh�Z�fx�68n�`�)
5�V���+7�u�YG���?\(��-TQٺu��]7����[�f��oz�۠=��_3���E��q|�Gy��'`\�9dQ�<��Oqt|))�AĪD�Q1꥛��a��e��lW��u)?o2�brEbF�A�@~�q3,꣉�Q������N;q_���"��e(v�\��b"�[%�Js��)G�H\����&��PR晴�8��Ț3y׮��������~P�'�|�UC���|����r�0P�uۮ��,BO�U��"16s�$�Pe���\�$������FQ��8R��={��<��]�Yf//,��������H�}L�:88���w��	?9@�M)&N@,M5ap�:�˦�D�v��Ud�-<�s�C���Q�~�{�����0�)��.B.i�Z�4>t���"��[2A��q���J�(bu.-��`m��<�������V��+�B(N�L����L��"���]Y�]����X9�KtKQ��:\^(c�·vV�Uh���������<�
x5� >�x�$���i�����1C��tS�XMwUc:��X�2�����߷m�-���m{�<�wJy����B̔^�f���/9��!��s�u y�$&���K/}�{�ݳ繊��y8;;7
c����<
L$����(��B�}�@zhQ�����pO��v��+K�i�Ɵdy�,z���YlfWq�
�?J�D~�t�b���"�ں���	۽��Ȅ(eM�EW������P��h���9Ps
"E��L�P��*���/�����������,ّ�r���;EI�-YS|7�	ɢ�ı��6^��/|�7�������
�|��_���B��k>V�~���'>���K��~�Da^^���+�9眯��a~�3�y�;�)$c�"&�-�_��wޙ��
�c�9і:���	$ߨ������v%�$㊑����{*��a�cO����K�d:_���[\��{�Z%���S�zrA�;��y�~��:�P���l�^�1�ga��1�DJv"_�!�1+ ~��؎��U�V)B�N'�>��J9ܱR4�������w�rk��/��Aiҩ�����$x6YHO�D?y����j�O)#c:ɱN�6��i��	9�C�I�%��@ �9�o)�$$�}p�Hn'JoJE��Z��v9�%�tè�ECr�c��3�o �k�E&*�����؃L��;�j� �*�=TWZ�Z�D��I�����.?�<E�UI������𦍧���hۚ[�"V�?��*-/UǪ..5ԑ���@�/�*��΃�h;^�Zݠn����]�Vuh�t�}�Ӎ\O�Qo����-ۇ'�w\p^����`c�j�V���@�Q��*#gj��i�)���Q �' ˎ��� �Aa'!����h���c[�l�0<�T��GFG�EE�{��f,��k֔r��Y���>bI[X��G�����~���|C2̳�>��n�v�ig^smX�MB��|�f.?:6��͕|96�%m���c�m��_)Z��*1u�tġ�%���(��Z��P�H�#d��Â�=G1T����ᙲ�+��a�\����#ƭ�8FD����0(����'b������	�����պ-��
�^L���T,E�50�נ� !�a�g�A�2dJ�8U�P�a:"�Ʊ,�C��U��X��+B�C4+���J#$�.����Uk����1f������8�_�|�&�o�M+Ѧ`�o >��T�!��)[ j'"�F�o�e�2-<��$,V���f�N:�<)J���d�?���E]������&L�����EEi�H��0
�1rχ�E���X��&�o�����Y��q�NDUt��h���jVb��i䲌���+%L/���>�۵�_����b�� �<|�PȬ�h|E�b�EI�3��N}U�s�22\��fUq�B�D�`sN��4��X��zSpW���řf�|�͌��ux����.���4��ʊ��Cr���O q�KA>Z$^(��S�617l|����LͥŨXTejiq�R��s+�����J_������њ���v�d�������#���b�Ps�)��DO6bjb�f ��I�����,�3�Ԇ�흖 +n$-��J!�V�dw���D�G�`��-!ߟ9C�
�;��<1������*�I\�1���t�Vܺukq`��S��H�Ѭ�~�0��%#Zi�7���q�xd������M6a�´��: �����v�C�X��y�$�V�+�D6p�_(�t�W}�!�hw����=�d�e�i���������w� SЎ0b��ʺ:55U�+F��G����������^��׃) ���M�ny�_|�c۱����t�vN�B���+�����\���~�3��������u�{����y��
Vs
RcK�w���ˮ�nfz��'�����a���G�����7~���ֺ"C����0	��
IQI�B[��N���Os���X��ܓ}�^vӰ�@$X�̈��0lU����=\d��ԅ
%�Q�:�.���B͂A%�`v��������5� ��D�@��B���o��_U8:6fJ�	斥��u�C=��%�)� ?0u_�8�J�>L�)!�)�����E���)}��_��]�.��"�Ta�I/��	 �G����-�GD/{�/�k��Gbr��ag/}!�|ދ���D�S�.�G�y�����x1��|7�I���!�I@?i&���`�UV��u���V�_�~�9B��А ,�X}����{���p߹�{�e����i�$֮]�E6F���Q��1���V۶m����ȑ#��Ħ)*�'�N�|�UW�s�9{�m@���6@o{�����nu�6!2��3�<�P�����<VY��a�{����c�r� |��M�~�>8�>���|Ǐ?��R#:$�QT�7 m�<11���a$\��p	D�<N~�}�K�F�b_��s{���vږ��q9�C�5�F�(��FA��SO�v�<��ӛ���yP"�//
��/��ڶ�FFF�O�Q�Z���Q�
�5�
"n������WE^��B�'�vd�sl9i�矈q�,F�\�}W,ԛ�nK�T����抪Κ.﵈�A{sL�	�qJ���Q��Eu)��ns���Q ~�����_����Ru�y�Ĭȡ���'����~�(�q����ŷ�\��k
'd�d{'��YW{B+�i@?3f�L�
c������
��聡�>~54 �&>�\Mж1N� $\9�3*�CR`��'GRNZ�B�[�{\�
s�d�5�D�7 4���Qe�{"+D1�j�r%��p��2+�j�0���^��":�Л���H�Ir�~!0O�@U�<�lN��ʠJ(GJQ�8��J���SR��0�G��ٗ����FtS����nC��"�p��c$���ōj�O[y�&Di��r�ر�X��`e �J����i��
)�Ӄ�Z�3SH5��[��V�Î����0�7�����֭�=zV17��o��oAN��;��;���?��?E��3Ϭ����ן$�4�mTe���1���OȲb�AN�Ar�~�lѦe!�U�qc��2DHi�{'''w?�1�W�yuÆq�6�#/Eњ��X��?�p�l���4�x5'b�b��ݵk��׾�� �|p��&�����:Fԋ�o���Ͽ������c��+�*{�b`X
rJYң��NfJ�n�S��z���`�E���$/B!n�I�:�"�`�(dA�֬Y��]�^t�E0:`k=���`k��:�n���/|D��g������0!��LHx��o����d>tW�f�J9U8�[���d�����p2c�������7�7YJ0<{���l,
�Aէ�7[AY7ƙ�a/��MJ��%��ps�B�����9ǳ*;�L��=�YL��^D`@���w���k`�]��~���ŋ=��]X���2t��]�뱣�&�x�G>����wz����`{�*��=������]�k�z7�x�7�m�{���w=�l�����2�^���y�lk��C"�.k�l(�Ao�(����G��	�����qZ�*��K�`�t���X"zŨ�/#{�{���Q#�鉱Ȟq��Nsv�'�q���IY;��ߟߊ^~3�_�'qvm�F!=�%,�Th�����:�_Om}zn�	�/��_���	�Ĕ[�n�Sր���O��S��;�������tw��ĥ_��׷X�*��J\RK���M�׌�O�,,-�w�iEd+A
cbŅ]l��`���jX%S�A�O征����V���c���y睧Z�ܿi�6بWؐF����+���[�(���ѓ���{�����UË<]��RAP�g�����c}���y195u`fjr�68�W���!WE�X���XLU;�RTd
�|�hRH��!v� ���=���,����j���{�>�lP_@� �6�ms���v�cK�����8]ۛ��^�X;�e�Mo~s�n�a92<=�\ZYXX�V�4�����rỊ��u�3�m3q|p�(��0ܘ�G�C�;1�Y���*QF���b.�jfA��������8��NJ��l�>Q2
��X>IqZ��>j��dYQ1L�-�m�G�4U�W�]�U��[�p2��mڲnݺ{�/R<����(��dA�2F�HA���`u-WU1^6
gXQ'c�^bx?�A?B��K0�$yq{RR��0/R�=h|�:f�0(i���U�%@�U;��
Fr����*��5E��s��:~�
�+���+`�]$��H2c!�`�a$1S�x}2
G��,��5$-�����Y�0"MuS�I����8L0�@��Q��L\�fc S������`X	�R%3i�6fl@��	��+��FT7.���JA4d��X�!�QCΩ���JH��@�9�1Y��@�$)�(n��BW�[ŔqA&n�Yp�xN��\\ꮙ)���aֺ1�U�l��T��J��/Y�K��+F�L-�U-0��U����l��M&�6�)�d<%�=D����jf����z]-_�Eiϱ� 
�F��,mt(,�ܼ�[;
F�k"�pGSjq�ap@��;2B�^r^�۝����ؘb1蛭�2
-x�����T�2\X��&1,[Qi�6À�KO�t+�=��a���cC_�p�� {�����[��Ł�>�q�@ֲ����tu�<�U�^�x�E�����DS?�g�gv���i�3�|wiI��.;�R�l��׽�0���
���
�>0a+� �)�Q���C\����YB��K����Z�#\wjva��<�����~��~��Z� j຿�G�_����G>v����¿������!�>�����̯�����=6=u�9kE��&��}{v�j�n�fy��.���#�������Zύ]B��Q���/�}�F�݁e��C����$x_�җq�9�7��M_��=`}����LI���Me�2c��vI&វ��*^���Ϟv������U$s�����M��{+)Gp@bt}o�㠢" �<Dn�i������F�t�?����#����뇏O=󶷽�[�>���/��l�m£஛�l���|��=睻3��z���]Q�P@�P+��&lߣ�4�������-o�����_�2����W�1/��n��z2�˶֏vp�M�/�*�a�Jq�M�l���������	�$�w�k���9~@ ����l�؃b�B�����̓@��Zy쟾�~�vۆ�ud����'� 9uln�E�U.�~<==�cǎ���
l���e�n�����X�{���>�J�N����|;�S3������ذu�M�<Iܷo�jY�|�o<�� ��"�\�#M0�����9��s���mtt�%P59�o��6��Q��ѧ~�ȑ�G�;6��yx�pu�k�y��*�m#-q݆G�O;~���#��ñWR!�P'N0�r0{0���!�-�Y}��aUǶ<��-�������΂v�0�hx��C�ք�òZ��{�����*�ןq�zނ;<��C�������̹�9��.���G6oެ�*hiA�;zgnyrr��j!6Fpae��)&�D�)����vt�<}�ՂG[��%ݦ�5<Z�ģ��Ē���<"1)����m�HY&���]ͭ]�>�xY]�ڵv����@�Y !�f�7{F�؁��>�̹�_��K�t��$l�:Gg�H��$E��=�Oa,�k��֭[��k�'LW���]�
c�t�XE,���XD�l���qSD3�[md��(�)��I���'8W'1{d���;]!-F璃H)���K1c�Ċ<�4����0�OR9����~N�;���m8�;^��l2X����c��r\�8�W���T=���U�
�$2���Hm���Ⱦe�B��9�ȴZ�ODٹp�����'2��ٜ����@�e�1=5{�駗�婩)y���@E�\���1��ǽacBc(&o����%�?/���C0 ����B�XeK8��}�7��F��{�n�4�D*o�9̄>;=��j(�Z��0`����'/GJ�pk�Ԏ�3�����	��<��3��$�q`��������W\q�կ�����x��� 22�,����K_��]_�7�O7�@��YN7�C�Ķ� &�w��������h�q !
(͆GG0�8�A��~�� �	��1�Uě-[yDM��	%f��=[y�'�h����bG^J�@ޛ�C=����y�x`a��e˖W�����-X��"ы)��/I�x�;��֣w�q�/��*\ג����?��3�<���p�W����������7\�����O���������?�AD����G?
���O}�����}�c�v�E_��W~���}I��E�K*?�t�WA✢|?N]a�ǵ�Q��K�1��N��*J��0�1߇��鍛���8�����Ç����oy�[\�(IV�pN!_x׻�u��������ƀ���?��w����L抩�S&%��H"<՘W�&k 72�ҿ�˿��w��s�7��JQ�(}�f�KK��/�Z?젪!D��?`��I��A�m'�B�e�F�$�p��eGtcP^Z<�a$�?�#U��Ɖkou����x�� ����D��FT�ǙU�E⪿P����gq^/����c��3>abG�����B�<1�>Is �So'���8��8����(�% {,�֩?&��b��D�Jo&�n��K�g�r����,�c%p:����pg�	Bmzr
t��C}lz_� l=mkca1�屡����P���<V��rSU,r^����X�[����xB����i�&=�M@�r��j�6��-�n�u���ka$��&��ˤ��d�,�?xxq�.��oކ���P;8�fl���G�(�86<:�f�Z��a쨺
�h���3/�ph���g�0��E�ڜi��\���;R��V!w�Y�`#�bߠ�=/d��ðdrZ�����u�6��r�՚��Kcx`Uv6�J�'�����ʮ��5�(M���j�����?�ѺuSG����TA;9gb#��6F-��O>Oߺ�[�Z;�Sm<�����E�E�rd)"�j����v\9�p"<	�`$�u��\�C�`��kU��Â�<�\)��4�q�+�<����p鱩��s�~�i�X�'�EEn�:9Y��W���5U�y>�s\�M��2�	�B��B�N�ShU(T�a?c5"�#��)V�x|\�#J���hV���Y`;v<���We﬌Ѽ��&=��BUQ.�	DETB�`3����i�%�51�~��
��R@�L!o�`*x���!�<-5Xk�B�Y�UIMTp\�b]U|�$$�(�s����g�0U;�E����Hʶ��?*F�?0���QO
��J;I1L?^-�@zZ�vI�5��7��

(&�`;��f��pl���Ş�4�UX�s���[�;p�@	W�Qb^q���	YPB��ж�&�="J{H5�?J�)L�����ȓ�q3�+X��*�ذB�OX�Qk��W�]B)��c9������%]�]��XU�Ɋߓ_bSUj��E�
�f�xIL�$�1L�{�8@h1�`b8�$��2h��
V�u���Zd�k�m���j�X��f�M�ڑ���Z�R���w0Q�0>��ж�}��q���+~G5���ὺ>�k�Y�
�L��܄,Z��9�5�lwQ���Z��Dx�	c��-�8qI�H�+QU�j�F�X��X*��b�'������m犃�C#�'�~�g띨����t� ���spw�����=Egf��x���Py릱M#��Ѓa@��q'g��b��y�7H��Y����DE���'P(�L�#����aJ-m�𾑌��b��dp
?�'Y�1���Z��AIQavt��23}����ޣx�O��=�葃gT΃&�p����~��w�9����!��-/.�^��_x�l`�����ٱu�E������_��>��n��%���k>�����[�r��|p��K.��<0�+�Cޑu��׫+ 0]u��`�($8�ϏG	I1� �q33�g���y��s�d�J)�7���rn0��G� �@�C��J�)��/�yvy�M��+^���K�i�ࣤp\���\w�k��P�w}�Q�Jk�&>���zǯ������7�xB3�PQ"�N�Y:�[)�b,�a��L����6��p�y<�݇B��� '�D���Z�9^��~�#�g�������ۗZ\+=�]N��Glj���T:�w/����?x�z���gq��w���/2f6!�}�ʘj=��A�߸u��?����?����=��;�
��������@�	��W��VN^B�i����ð�ѣG�KxP�tAU����J�O\j�/��И�������#G8�:8`YX��g�7���~��6l���7���χ;?���ā����K.��$��%{eϞ=+���?�a�o��?8��x�������秧�˶%�Q�;Aȵ«]��I��~�\ڑ�,-a�����}��v�=��*��y����YG�@�\�n��?�M���j���5����=�y�zx��I������\ϑ gT�8��	�#YIڌ̽�;��^�0���!rI��׮]����7o.��U�6�mڰk?���MM�8�~@��	�F�g�CC܏CA��a��b�*����"�)��qQYL�t��2�3p�X�B)A���A��C�"����"�n*r�k��Pj��i:T`Ǡ� q�4�*��_���K1O���m�6��43?�lr�=�ܶ�[y��q_B��)ڃv��6#�B�*�X禒W=�pHV�؋����9��N�(ncd,E6r
�z�!����|2��)0u�XK��$b3�%�B���Ld~-~.��pZ�ل�=P�T�Bx�-ht���T	l
�t�-�ڴ:�1	a!ڡ����;H��!b��9��C4?��Ⱑ�n3?)�J���҆u
s~ll~�
j7�`�R�F�a!���l�-��P��FA!���y>~kR0M�T<�$!F�����O�;2њ�f���횱�+�z�Y��Ё�K��h�.��3�"���ipI��#z衻��ۙg�y�:t�ء#�1q�	|H�SD>�<$�ga�A7;�!�|��n���á�aV�r�-���v�@�v�i�)`��@���{>�Ϸ�i˱��K�_GIz	3�I���֩����	���k.�::< /��=<Vǃ?>OI݈O��0�K3�{hh�2,���h����*�T�	�I¯�9�z8x�I��%Y�R�j������$ezz��0�o���O~�w�u�΋.���������=0��ջ���Ç�u���8�Jٶm�H%U����o�馻�� |���n�r3�n��㎫��S4���b��L��v쀟gl߁�n�N߱�'g�/BfgD�'��I��j�+�|]1���z8&-�Sx���tA2���Z��]�uBB���{v����{�n�	ck2�x��`�F��"�����:�n7�p�?4����7\ww�e��᫅�Ɠ5��#BǑUČe��|ɤ=�u!���x������ٝŚ_Z瓰���������๏n�'�OZQ�})��	��'�2�b�W��R���)��C�X�rb����)���)������p\�[�iLT��<8̞~^bR
F��	uY��5!^=?����P��'U���5���ȑ"�qO�&���tr01]�eE���a����:�ƒ��Hn./���ㄚ
�Q ����_�n`�ʌ	
蔲4�߇~t��\P�U��2�/��n�Z�m���juai��l��b�b�m���ĝ��i������c�!��\W�Y�fVȠ�9��p �*��k�־I��]�O>z���j��Z�N�@L�y/w`ӌb��-������Ȱk���ٿ���r~tbL�8�ե~��rY��N[�j��*����mV� �]�� �N C�Q�v��N�PDp�(޸q���#��&Wk5�څ���r���&�G�8�G)_0"U�w֛%���z�.�|�����666X���նsj��/��S_\�F��`7��JDU�X���ֈG0�1�J!tb�52ʅ@%Cu1Va|�Fkׅ�����D: �lmܶ�R4A1I�xs^�V�k16"۩�L;��{��=�|30�ϵ�쎍�j�R��{�O!��1f|�B��;1"\S�G�x,m�:�eH,	$�Q�L0p��G<-N�.זa�B�ʅL�F�-(�'�+��nU�vmF�9��=Y8��z9��F���J��Łh��mH�>Pyny�T.��կ��X�1���tk���'gg�}�ە<�����b���8q ���J����1��
cD&���-/���*�=�{]EPMUR�_. ��3��4�D5���4$�F��f,� �6�"�=� )$�#�����5�$gx�Sl��L,T4y�����cΛ�S�Α@!�刉��3��E��	��Q7���ǫ;Tt�.	����e[�d�S�%��W]wjjJ��GX>%"E����=�C���F*��sWBE��L*��芑�
���ԉ8%5��L�O�����2g ��ND--)�wB_�XW� M�;�ĳ�T��ɣ�:���h��G��Ao�y6ti-��y�m{n���������l��a949�ܑm[NcZ�\!k@�L	�Q��������	���A�5�k�(�P/�qH� ?V�2��`pWX�uk�����?ؼys����1A�K5�jMHR>
*�{n�x詔���F�|�����eOPհ�H6�_�ƽ_��´P�� wy�u����֎/��9f�ad_u��G��.�A/��j�͜$���F��D��O�D$���d�u�'����b�4B1Dp�<Q*|��d��=='����;���/^m�@Y�#���~kϳO�>�r�-�V���-���r���Z���/~��3�z呧��⅗^��>�>��$W\qE�?���t�����<���������o,�L!�<�����������������5�r�t`�����'�|rh�F!�h���p��T/s�	A�s�_o�*�Չ���k��T<�����Q~C�D�n�h��j{XkE�FVC����M9�q�&ׇ�_�����(�����1k:�UYuu��k���_>-P�(B욆��ǿ�[������Ї��@�"';e!���[��s\� y�%&�,�p��d��?�f�g�x���q�A<�!���h��_q���'���_�-�'p����|�� �?ɹN��	qΘүQO"�u��;I�@8m��o�R��p�
�Z	�5�t�ݜ����h$KH5v��5�Z�%(m���Vg��$����#X�U����9:�5G�(�X�3No�G4�Gyd�: W)�}���c�i6��C��M�6m;�c�mٱX�˟]�v������h�h#�2��q}0(�qJ��.��0��9ʴ�!J>i�z�*|�������kׂ�w��ah0ܹac8ŋ��l��3#�U�Vԭ����v�0��m����y
�W�<�m0t�������,����^��#0���Q("{�c�{�[^Y��S�~ⶮ"�⇛6m�nʱ�UL*r�#�3���IF�(O�r�x%p	V�<`�id c�(�긄�	��FP�l�ѣlC��~2W����<��)`Z`;�=��&���c�nB���y�*�-��C���k�ǐ-�(�`�B#� #���ajy���E�y�g�J�N���<��r���wh������'��O\�lo�����ړ��[�V�O ��M =�T�~�0�����&�HI�	�"�Sv��?�0ٓ��d�O��4�Xm���@��2��������01c6`�Fb �P���O�'9�;{�Z�J�)��60
0[z>!��Rf2͊�$R7� 	�0�	-=u���.rDK���"*<��xU���4�K�d޻w/�m���S��8p�ȑ#��:>g�?��ə��;�����>�Z�{��F,�'x� ۖ�#��v1"����t%��8�1��RW�,"������jH���|����-p1"�c ���bW��
��8�g(����%�-�'*��x��1
J!" �H�	-X�0G������1U��Z����J�rٹ���N��QIu������흘w��m��i�\�]=
����B����m7��͊�qH�pK�\���~��OLL\z饳���U��3������۶m[�~��={p
�����G�=��6i��.�������}B����>W*�W]u����B��ףGzh�Yg=��wu]SB���~��������}���,OA|�a�; �TVF��4�>KE��:�����b��f2s�f_�DN����C%A[�>�EMM�<�+��493cZ/�x����#�|��0��G����q����d���3��c۰G��e���"�?'�˶�9��֤أ�"��Ȩ�#��J�){�d����Y�p2q���~T����y|�ג��$�&Ӣx�
���~��Rʩ��0N��̧��i�n��t7<#��`���(<_� ֍�H���9�� \&f�Д�H
��D>� S���6@q$���@HT1샪�x"��&ٌb�PDG�8I:H	Uib�a�*�K����@�)TȎ�DP�L�ķD$J�:�|����جrbp#%��ea}���9I��g:�Ú1���#����,� �̂F��ZA@����L؉RTD2<$Ղg{5�Qd����{�b�П��b�@�h���v� E'�ǲ��"�����r�����
�����w�U)�c�ã9#�V�̫q���u�!�%
�T�`nv�+��6��@UL��EDK6�8�ߗ�Mk�Fơ[�"&L�.��G�+���̳Ϩ7k{�K�ԝ�]��-�=��!a�y�ê�(�5f�1?��`=� '�[��P��gCA����
Zȃ���n�\>�����鉵뭵��Ԃ�d��LQ�5�i��˺Z�7��Vm�0��P�e՝]����&i�	f�SȅOpR1M�ClC5y�Ga1��N}鋟_��Qo�q�$5�:*��~��+圬�b��S�DcDcN��cZ�G�hj�'g����v�{=FHq/��H�J���<�����Z��鈅}Q���t]�ZD�2uD�����F./���&�"�(����P>L0�m.��et�Zh���{Jv���0R����u�o0��r=��d	�k+[�l��������������������m�����n�������X���rh�QMZ޴�:�m#���������"��� ��.��`1u*�z&O����y��f�AY6�bk�uU�V���t�0�[�1�j�AKA�ݱU5\��t�?dU�:�l4;�(�e 2X�y��a���ѣS��@��ᕑ4<�I��q �����B�>{��!E�PC㍜i)�2��E�n��A�\X���`i�ל�?�ug�p���&�s���2h�	Xza�� 
��r`��$�in� �0�m�]5x����e��AA*6T����$Ib#��$���¬T��)���������C�x�2.�ks�ˇ��K~T��J�����J;/�j�����������,�;�>������w����}|T���:�raj������r1���Q��<
Ȓ��n��x�m�S|��@�Ra*cڶ�9�'�%ύ�"��y�L9��q'Fq��t�š�A�[�
6��I�b�"�D*�����h/3c��nY�_�_Z��t\�����u�U#�:���j�P,���#}o���A#��������\Բ���k��v��Ib�-��/�C��Dx;IJ�)5Z�llޯ��+eS:�o8�UB�a���	�]q?�d�X�|d���/x�����X�����\s�-�{`�A0���,l�vFǏ��Q�;o��������2w�!�zl�>�>_э�;L*U�E�T���}�}߸s�������v���������&� ��.	-�Cƨ|�w+Ośn���������c#�\�š,ɫe�"��q�%�~@�\,F����&)�?��z~�u�v2oEoRL�"
=fp�d���F˹�jb.1E�@<�{﷧����˱��v$��;��+�񶷂��v���/J�����y��"#����{��箏����]�6u%Q#�&[<�i��"�]�E��~������}���@f�Dזpʳ��D�{�+���O��/�Z?�PUHL0O��� �@�C�C�3��@�Hb�9�-���1A���_�{ 梀��#O�y�L����M�0e�c��S��(m�l��UHb�d��!
�E�6콣t��q�AL@o0��tM��ƈ֫af��ɸ;�Ƀ��rf�@!~U$�1T2�0Õ	!�:�i�(������#<P<I��W��2�a�&1�)ϰɱO4
3t#��^*
'c	k�����d��φ�@���C8�jZ��N�S��N�X��`�-J�^K8��'B	�ý��P_��ײ[�����CCC�
��W�Vp�Mɍ0��@�,��C׶}-�C[�\.#B��mrʟS*��'��ϧ��-���j'�z*�@�n����֢�CSUBߊI�S�R��jp􄫘������
0aA]��y��������i���w�.��֭[7���6����L���P%�yi���5�[Vah��-*1��&�3ba��Cк��???�C�S@�œ5cݺu���J��4��Y��#���5�+X[������)[6�qQ'tDN�H#Z��D�8�dQ|���|0r2*<���p,��a!J�k�=��U�<���|Ď��c�Ac���t���*Hfʸr���x�O?�s��vR�2)�
�a��]n�k�p�hoBt���f�	��!t
�i|𑆆�&7�b!��U�``ӶY��i�q�ق7*�����	ǎ�0�<
��)t�g���oz	���Ȧu��n���`o7c��E�b��̋SHv1����슂�MW�ex���%����\X��"�!a�p���tlfQ��<
h�L�N��ےɣ�&^g.�b��Qk.�U�EYR�rL&��,�ѧ��\~���8�q��c%�׽ͳck���k.4��N �3{##)�U1�Z���2����Y�����|�'�������I!S(��l��h��N������̣�{+�á���;�m����̧?���G��o��V������Gy�#*0�V��?򑏄�"����Jex�!Mh���(��4s06��_I��u�B@�f��"i嗶P2�Zx��\��N�=�����K>�f��-`����8��3L9�z�NNd�G�	Y0��C� �	��t�#A�����0��<�0V�r�*��!���'Qy9�

��\0�����o|�T��!���Q2Uһ�6�O<���o|�[n���h�B�cǎ\N�A\
�̈�AJ_�*�^��W�+��_=��s�}��cG������8Nძx𪫮�jg�l�bs��bV=�?�*N��`C�a�%�]��Ybg�s��`ToW�)a"�(�%S���, �
�H�RqI*Ůӕb�R޴i|r��w�{�Q�k���*�B�y�~F�am���.���W��U���'��}>�/)�١Xbb�����;�;6�����{I$p��?^��~�ᅘ��
�]E)���x>�$P�"N"Š�&c.<����sF�w7,�\� >�0�h^����I�2;�aapJ��T�u�I8���=�f	Y4�1�Ae5��bJ�	�Mo~�I6�H��
ؒ����Q�#"�/�!Hǜe"���i1���ƨ����M�.h�j̈́5�Q ��#���M�% ��iB����=x�X5BxI�I���*�A��C�d,��]��DD�R>[��X������C_H���>U���e���P�[c-֐�����P$*��p�<z���Hg_;��C*$�R�
7��IR�����󕡡��y�_&����;��Y;<�t�QF0�b�i��X���9�*�VN�y6��`M>��Ӈ''in$�ʾ���?0:,�-P�%��#���Ɖ��0@an�-Yb�<��뫝����U���%4��$�8U���H��T��@����A!�-3�1��������Ï�+ �eb��5��L���������I?����d�kԚ�P0�&#"m๪�xة��#�w�S�.%9x!,99$�]5P6apA#�&��u`J,/.֫��۷�OLlܼ������j��#[�UEڲeXe3�l�b�A��EL�j����|\4A��d�1=�(W*���+58ӄ��U &�p1aFc	�*�~!��<�pn�ck����!ж[����֬��6�P�3ѽ-�]7��CUAc��EлA�� 
bT��YW(���W�����Ԓ�n��i\}��+�z����~��kv^�vӦ�-kTw�U10WdA75x]h��[֕���W$��n�J�f����0a5�?@G)Z̇��[͆$QLL!:� n7�Y�1e�I����&E��n�Z��W��[�ծ���o���[?
�%�\�m۶�{̃o>��+����;����l,./��Y���h���x���rQ2��.]'��#�%g䠝` x�Q�Ć�|��a���֎#��U�Ě%Y ���.,��ζZ��={`
5��.F�4E�
2���j�9b��5���s�]¼������B�i�A:������ʇ9�n4�b�\(w�
�F�`ǉ�h��-s߯T*�x�3==�F����Ј����m��%DB�þr���%���Sʣ#�Q��������!z0}�	�y%��Ȥb��]�W�ۘ��(Sk����k�$wb�EuY�(��&V���;Г��GD��0qEbIT&��T.��_,$)'*�1���RH��>��EnN�=qz�h�!���Ѩ�:KK��k��Eì�-KWj��ŕ�"�
3s �NUe��q�)�wT8k�O�	RGE�,[�W��)�4��ҏUy�.�3}�"�8H��e�鄹��&"6$�bjǁu����*���Hs�� �>kp���{Q NY!�z3/`'�shg�S�]\�!��[����<)������G?�����wq��%�2e]q�� ��c�_�hߗɺF��ɚ{�'?��,+�&&Jj ��I�. ��N���L��1��yU�/8���>�j/��w�/^�n�~���^�+�7��`� �U�|-m��*D^H��2��֎^z�yw����߿�λ�>��k�]�uW�8�� ��V>��\�Օ��Y#�޽�����a;CJyU0f/F���%Fl��bOG�ȡ�J���4%>�\��c5�MG���Sd����$ɍ�ĤTM�
��\_�L�� �~��������ܴa��z�j�^�D¾א�3�����.Ef1?L��O}�^x���?-�,�M{!l���``�kz����}��֛��^�:�qd�� ?��˶�9TEu=WT��j�LX���<F@^L�=�`!RD�M��R*"�aFn7�45�L'�ōJ�8�����Rx+�籉��H᯲�v��\�KV؎b�JV;��v��z��b�rE�0�lAG��FX��7�1���uMGՖu�0����BB�G	T4SIf�E �0q� �"��O�2d�`)�v����A�(��5k.13}9�� �6ZY��ђ�[�N�h����~�ж�����:7X^`hY������i�\���g�D3�&.uΩs���(�)�b�9©�
Or\a���b�iݖu<�@J���/�l\�Ojm���Z�T�'�f\�f͚͛7�66���h+�J��N���_�#_B$:I/����juaԌ=rN��]���WQ���8og��74�UT=Qf�l��~�V3LhG�6ll-U��^�k�.��}0��u�� �,h�����޵�~�ŚC�}+^�uxh$J/�|��.zD�՜��lc��83�@=C-��0��Z�ȑ	�?a�aD�ʡ˰�233�hBCCC��-cdC�0K���@�n�b������b��PJ�	�v�wY��(�j���-���a��?p��O/�����td��8��Lv{�b�� /4	s���	Ì/��8c}��O?��`��۷z���ӌ�,P�� 둎0�9�|�֮֯T�f`�x"��A�ar�1=r�.��؍a�����U���XkV4ԁ�K�<:�i�U�P'�q�
D]}D<�Zlii	f��W^	{�F�ۃ�
ܧ�Rk6��~���}��g�l�y8ǡn�/�e}�޽�jڜ�`TDq9E\��G�P�%1f#tц�Q�&&��W��q߸q#�X}�n���>~��PԠ5m��@�%E�~��!�k�r0�ALa��
��Q�x�D�����,� M鳛r$}c�]�;�FxS��!������Ckm�����'a�pj��R�h^� �lw|p0��ĩ���DĿC3�f��4��.����c��ؓ�|�x�h%�$K-�$JC��Q/�8aa�����"E���*t� R� A��%�Τcrr��}3M��v�vL,�r�<�,��sND�>2��o��d��|&|H�x��m`hg![�����R��9�S�)�� t���wm�b��e�p�v��1U	=�0��-`#�O0�퀭��8<��:�&<�0`i�#K,��K���R�<7Čw4�}�yNF9��"g�*Ac9 ��A)^���g�[��Q�$��?:6���c���믾����J
^���������ʯ������SO}�_x�[��oI���
���G{�sχY�s��9t��ra'��'�)'ro���"������0%g��ĺ8���;���_���q�q��$�F!��ż� 6Š_}�0���[/��_��_������{�E�T�@��ka�p�4gQ|��u��iptt��o��O}��]�+��/G�v���Ga��|������߳��n��Pe�)�T�y:^��~�ڂ����U�Z:j�"��G�!���N���T�八��ǅ&��n)X��� ��Aq��P�|���ȗ�F��S�e^fJ�~RNERnH�;��9��N�ݎ�w|gN��˹Z��8��9�q��uXQ�
M�:dY����!��I��)3�`�� ��]*U����j��LǸ��zS]�5��G D�Nׁ-�j�WƷ�>��Wݐ}���� �	聠6��=Do2�\I ��Ʊ�Xt�����4���n 3�b�仂�tr�q�O��ˎ�ė�� � �@f�ĉ��5��0ڒ}L%�ѽ��H��
�B�����Q��2�o^�n�ƪ�mھ�@�Ǘ�GWf� �&�t�BeA�"Ce�����8gj�1�	�<��y�N�HV}]-��jy�T�V�1Tt���#)NH��\�X(��BA4�Z�hd����@T�w���I�ռDO�8T�t`#1�lr���%%ʩ^�)�ډ�g��--�&da����`l_\U%R�e��X���_b�/haKc�X�f�p�!H� RM���`xg�vqN����&��Lŵ �f���m#��+(��f�AAd]R�0^^Z��{�fYU��O7Wխ�]�]�� �A"3*�HRt�10�����<�4��i�A��)*�d��s���n>9��־���:���|����[�N�g��׿¿TY33�v|�-;X-W�x=�vj�S[�68o߾}p�h�� z&��5�a��;*Mz*��c��pf��m�B�D�p�Tf�A��t����:H�J-��7��)pS(E��	"率�j�J��B����}����x6�YС5�(v/��#Ts�j�ƕp=(���.��hkgQ�7C�);���r������oW .�)C�l���aqp��%K@�E65>566V�3���3{��c�h���t&ڂ��Lʣ���P�w����]|ښ^!Nu@���b�]�������-D&MŁ�9�m
��ǎ�s���(�Fbg_�E4d��%��aj!C�(S���Hލ�Ս�rc� ����s��C��͔��Z��r�\)0j�4��8����U �3S�uEk�#�DA�@�O��/Xn9�5��"�sɸE��C�`��U�r�e;�;"6 VIL(U�'Hat[1��ԁ�	ȌTu����Ct|hj�4s_�ɝ���X=�ikC�k�� 5��9(}h�эfm��� ��P�RM�l[�$@z�`�ގ �y��M
4)�#{��3XG���6�~v�n��1�xy�A�GT��8�Q�Ĥ�"�c�x�.��2ob}7�'a\��ǁc�t#-�4i���l]S2���������u$ ��)k�H��w��#mz�%����A�D)z���X�pc�s�q�Qy-����8@�`p�����DK���b�Jg�)�j��QАG�k��h$EU<�hct)�P���7��ܺ��{#��gR����i�Q/M!H�3°�P �04�/���8
�9h�EF�y^3a]�7�2q����J-1O�>��$��j�4-���;�"i���~`��[�n�ć")�F�R���@<��ƶ]~�������t�I��蕽ł��z<#����r��޻ed�M7ݤ�>R:y��D������ܗK���pp���Q@7ML(�u�!]n��������t��?�<t����ν�v�����%� ��=��x,~/��"�R�6�M����Y�1��2�S$ZGb|O̵_%���9�y4�E$h,�Q�S('JU��׭��C��������o� �WІ�O�z�_��_;\醚v�@�@��e�@�禿������!���z��Fv����_0rI;B[���~���UL�A��
n����	Y/p�����඄���_�ҿ�������`�X����\���W���?���fr#���s׽jrjR!��%˗=��S��,�ɞ%�FAd	��Oa���$̓9�� �/Wn�N�*�=�]��-nh�e�K%�8<t��ϝ�|��-1:x�DD۸H@(�>?�s�w�x�*��""�a��ޏA�r)��P*�7���o�P#$�&P"	�:��|��m��iM�"�6<4�G}�45��#I�v��+���o~��qWx�kϿ���f�2�[�~h  `��u�y��1�K�����ٛ��F=��zL~$�A-Zt�m�Wвl�PAQ�[}u� T|8�Ǟ��Vh�r=��3��x,(�~Q����0#6$���]�vi)v��˗�Y�fx�^�����4W@y�:]��l��z��|Ga�Ν�<����(U�;d�B�����es.���'b�����͛7oݱ/�{
�ɥKO��EΟ���{ ��Px*���j�#����^G^��^k��]����z}�����7,Fydx>��f	\;�[�ׯ�54��3ϬZ���/�����,]����dfdFd^�c```|����ll��対ږ�) :���߅o�·7=s�i����ك������0"7�۸�oT-����*����vtu�Q�x��`AΟ?_�V��-�nY�eժU��Cp�q���(֜n�|�	����{�r g4��dr�N���j�J1e��6��#�"P���1ծ���\'��m�첀"l��� s��B?W�Z>�d�2�M60�ԑ�
5E���_��݋���]�������۷�MڣP1��h��bE���4�3%�Ea���DO%:X�k|v����T01J�z��ǽ��l��'?�A���믇~����G���/r����[?���e��R������#����sϹb w~v�p&� �iFա��*R�gcF�w7��B>����ٹ�_���wn���7�a��E�WVi���D�$�6St#��޳l!�cձ8��#�</�90���sV��5�՞m;@���;v�ׄN:��`z�*u�}�{zz^��+a>��.[�@�2���s�}��ٻwoJ0ЃH�0�2����344��K��'Sq>I8WS����;���𩩩f�n��(��&&&`?�[���s]Ј��G�����4wI�/����G�<����pN9��`tF�߂��Ȏ�w�!����En�;�����B[ʙG��˚9�9
M���. Kɾ��&c}<���:M��NT �
|[o'�����"����l'ZH����1"?�a-o��ـ��ẗ����b�b�U�6ˉFqdӘ���9v099�K�� Iac��"��=��c\X)[�����@D80ر-�E���޼l�����N>���I�W�{�����������VQ��߈�11���/9���Ð�(
b�]���(
CBԅ<�o 6��&��X�d	\��cO}�S�eX�	����F�(���W䎾K/���q���Q�cΞ^�dɺu���e�O[�t)��
�M�D������b�p�W`���SO�y��ȿYާ�����R�u,j�vBt����i�I�L�!$!B�$0Y �P~T�����Y��m͑n*��̵��:�zb���9�YƘU�E���}�C��G٨���4LBNLJ��J�|�󟇭��e/"G�L �z�ˈQ�>�ɏ�㷑a�����b7����ov����{�Ix��T,j���ׯj�g�0٣c�a�efN� �P+�Ä�⊷��׿\)��55�U[7o����'�9���V�\L
E�(�L����
{-�P<.7=&QC��[Yk}r�S4g�`���n�cBx4H���He��R��%�"���<���bq�%��&����9��W�
�+	)SE�+�Lg�[��I�h���3�Sk(R�I\�/����q�Q_�섟�{�駟��Hj<�nI�<d>d�׿������"�+h�����5�o����-�����T�5'��w��,�:��o}�[>���}�����b�N]���-���L�3:C�@�#Q���q$o7�T�f��Ԕ��ta�U,�-N8H4M�k�D"J��u��Z��Q�t�LNN�<�,���Z���N���L��+V�E'�֞��V볬��Rm��'�������v Ī���*�����O�<eM=8>�����4�e����r6'�vb�_��]A5;A��;�ci�T��V�<!��Ϣ@b0bH��}�ͣ��z��b��BF�?G��Q��a��狦3*�7�*�tՊ ���fน�<<�FL7����s3SR$cѠ�x�c���|���cdSZ�T���l��r��ܹK[HX�Y�bE�d��l�Q*��XhD�x��#l�"��J��ۉ1�����3� �T��ɏ�������H��EA��1�+��Y�&�O�L�{�/�|=�3ɍb�f�:b���!7�˱ّفf�r$�U����ly�-�3�C�'?=�����E1E(Ţ��-�m�8~	�_|	<$b�E3
h�kȪ�j^����j9��.�p˳�zOi��x*�$ø^�	E���1���=l���*��R�� \!7��	G�f,AF�8�������ʼ9[�l��+ʴ���:��N���8cK)�Q��]Y֕-�t�539�r�������ۙ�7�������͓��@�\��R�2��ǔ��V�-�&�NX�ժ����y�(��e�II�B���`��I����"����.� Mj��� ��l��'�nW_7�f�Q_V����ݳ�Nmi
Fsү7|��a������ѝۗ�3�;�,�b3��#�B!O~(�^���WӤ4�1 �*`��������C�@�*T�9͔��a���L�� J�:@b�a0%\���_Ŧ2G)�HHBE~�0j�I��
B]5�MMӲ��eRH4�|����1Q�(pc�/�:A�"�P�WRN�T�؋&E��j%�g�g�蘳!�2�j(���h�Z��D)����I��;����Ua���#k3��!��,��W�B�ܐ���6}5$U�YpOLcSⶆ��*܅0�b#peM�xf���HLհ�ar|��H�4���2E�ĜX�6T���Ti �׍h�n��wl�8V�v�p��.�L.߶}[���.)ƈb��dQ�*�B05�0N�����v���A	c1�o5�BX����c,"��UD �
 ��k�@�xo��Vm�?��^����H�m�0��X�-���:R��"2��A:L��p{�5p�@�e�c�(��&�`s���:3�
J�F�Q�#�b�8�o�S��B�y���q �^��d��Fe��9�����F��"���<�a���5����KސEKn]S�XT݀�rn�L��m���O���o]��`ȇ.�s����?�ՠM~k�J".e
+
�28�}9Вe����X[�-���8<@��t�$݃����t=jSs�� f�=�������/����Y���U��&��~��0�����T��!���)�K�c��o��gn��O�e�C*2ds�W]�η^�v�0Q�����\{���Ma1&�i�Z�);��E� ��jb�& 7I���o��z	k���=<Q�~��?��@�VC2&*+��fo~��z�!����М�=� ����W�����?���Ů�'���t�r	��i��Y�p�$n��%��&�.n��ШUG�_���u�o���K�Ј�?��Y�V�E���5�q$ƿD�	�2��B�pG�Ҁs�x��W�╰����'a +Qa^4<4��W£/���GyD�$׈B������_,�����(�{�����/}��x��^�dd�'�%v -Xُ=��_�Շ<O���Kxם��AR��Ǿ�����[-Zt�[���<��|�_�@�5�\r����e�֭�����.��µkO������s.}��~=� �*���:^@u�����|ls�#�-Ph�F�3��8"��w�O#���iST7�3`_�6fA�\rB�M7ݴl��S�8�ԓO)�˳�h�>p`zfff�v��ݻk׮6LL�
���nx)_�����l8;[��7mBް����;Ｅ�Q>&�T+�+�1xix���SO��:p���
(�_��pF������G��&S�W��aR����Ø>�e��w��j�'�h�
hip��cײ���u��A����=ccc��o}������^rɥ��������{_}�+������={�<�裘������w�g�7呱�N;m��E�'�χo:Md�sm�v�C+��(�X�p����4��֌�O>y���6m����2���'�\�da>��;w.�R�K�R���+vv��6l]�|Ἱ�������K%�)�,��2^ŗ� ���)-^�L�z�
w+�"�����~������{�`zL�<��ݨB��@4��1g��[�0����Li�0�� v,+2�|ٮ�e˖�MLBN�����=���u�W���:���=��e�φ�e�0���\�cpk9`��:�]�����ss�]{��ui����.3�ρa�������1��(c�bQU7o޼l�
,��0��s�7����M�����u�]���s�ܤ�5�(�Zzӛބ�'KC;�L��037nV�+�X�ײ�;w�|�Yk?�яNϔ�����Yx;m���!��G�Y->@���g����Y�����P����ַ��ٽo^��~����Y�����;
P3����4Ӱ:`Bں뱿�z~��AX���n���<�
k%�q�bN8.�����ph6w�b6�8I�:�M W0�9���ll�!���}���<��OJ�=�R�-���!�?�}B�O�A��l�����P�P"�I��YNP�~�T�����]d�o��V�b1<�\m��[�3�d�'��rCB���yԪ��	��6ܦ�_7��1�m̍���zX�<-�ai�?���Z/�����n��/���]�j �+n��ե����R�w\<VeGW'�`2���i���[���5�o�{�" �rO�H/��a��ۺu�`a||���O_�v-�,h|�R߽{w��®�k�^�eW6mرcf�F����+�G��YRHM�6
��Eݥ�Я�)�g� �ox׵n��(�� pHA7j&2a�$�I�Ƶ�r#3�}����ݠ31K- ;���d�G������N90zwo���k��&
��k[,[ܿl�O����� �����k���ob��d,�p*d(a���;���o	�X:�gc���T��u��0���Z��q&��+-gk�"�h]��6�EO�*�zż�~��o#⻒�$@VHOM��1Q��i�YtZc>�T��?��#5e�͂ �^c?��@�|Ѣ$��8@}�ޱ��� �V���Ҍ{�/a�#�v�+��t�jj����W������y�ɀ$aF������'�o���ݹ��5��կ:M#|��f��OAw��ڗ~�����-7���xqM��Ϲ9G��,H�M{�#ke'����*��;ǎ����Wh����܍�Ҥ�#�Y��Q�cM'�9��3���R��"��*׾�u���˿���W\Z�kiIe��`���N��������7u���	f���F�c�+� �x�g�������=|�f/(�>�M)-�r������*��[��6P����+b	�u_Ҕ��?��W�p��g�s�:}݅s��m�~���)Ʒ��-&���_�������7j߾�sN�k��=���^�j��3�~��?"��U�ÈB9B�[�(撎χ�MK���n��UQ(�N��XW����*+�Xp.�0�]�C?�/P��{��7Cݯi^�.�C�o����ONۏ>�qb
���� �3���V<gdvz��ضk���)�d5��z�ېԘD�L���阽�z�6ﴫNW�?�Iϛ7Oa��,A�t7=;[���=t`�W,*z�I��*�Z��3�^@t�&^���~�a�y�
Z]ZSƴ���k�\6�����B��ӫG���� #�X3��É��!����&�i3��D�r`j�ɑ����R�{���riz���ڹT]kB`{��T�ӓ�Zk�)�d�
㈙W2���*SP����!�JD�B�B�VK����t6�h����i;r]�PE/l�Z���I�0/`S��R�r� ����Nd;���u]��չ9�%�īa=h&bU%���X�ȱ�3]�5ɐ��Gz!��bgz��ɉ����
�?�����"\�������mߕê���[��0�!oi=�pL
�(������K-X�<�V�̨�I�Ο��L5�7�V�E��E�[�L��:�b��@n[�6DQG���|��|�6ۻmKŎ���:89��y9)5xE��7s;��b�� R����),5Ԙ���è,J��w�4_g��ςR����L�Ss#Ao�3�l���.�[v뉂-�=�=�����@|6�ͤaID���{������^=0�LM�S�r$�� uX�����UX�q�,��iO���j�αr}������(���g��g����R9<8�M����e_�Bꂗ�
#=�`0�W>LR�X����̴�Jw��Ն�?p}��J�
�AbQ1�	bL���f��r����`���;(�dL��Z6L�ت�
����=F��R�"��
虔��AYK,/�A���p1�P�a�]%B����W<'�]�Y 㨀L@��ze �ǻV)���ZlĹZ�h�WtA!CE0|�c��^WB�GV��aE�V6��ŝ(�E��oRU)���1��D��V�,�E��碱GU����XhDP��� :-��$�$@?�0� Z�
V1Y%D���F�{C
��T)"�h�AxA�����(��JFr,i"�=��Tdׁ��̈�E�St�.g����i]�Z�l!�*�}phvjXTd��P����^�
;���ê�9n`�=6��Q��6Q,`�8)��H��K�`L�@w�ժS��$N���3U�X2ǔ�h�����jg	_�^-��z��A�{5�=��U�4�*�#5��V�� eāb!�b��cNR}�����T'�g�ܺ��͚iXw��-�m\�3�� 9�f��˃��h���JW	Z�L�1���ad�A����#��@}��	�I�.���0��v�ƪ"��Q�s\) B;E�j���x�h`q�/p�j��)��ڈ��&�AKq���	WD��,O���0�$�#�����I�y��g�R?c�H.gm6\�@Y��s����x�ʭ�anr��BSbTS|��a�8�dYIE��)�\$�PR1z' +���Kh8D>�S�A/�1E�]���+B>��`Y+pP$6RjkM#T6�n�f�%w -r,v�#q�%ƚ!�{	k���	����������|ӻ������\�`F��%�h�|�=�����G>�M�$���|�fĿ�˿���700���?���i�X#\��G�\&?���yE���?�я�g�����.���ݔ�B�B�C3��7�|����	'��H�`��t�V�ѹ�)�pν�<���'��]w�;�����O~�c˗/�4B�9_W,�*ɋ-����������|���Ok�O�SO�٨/c�p�`���4LX������]����瀵؟�8fƼ��t�PT��Aα��>^���u"�!�	I�������/s�������c�%̼-��Ȥ�L&�͡��f��ԟx��H�[�H,��֭[7>��<�+2�M"�8��\��=;��)�)1'��p�T��)"1�`�"m�F�.r���G�*�I̟?��裏r�<���c��ի�v�ʷ��mi�9�k׮-[����r�4Э���b��?22�q�F+^�����a����΃w�ڹ��՟~���� �&�&������+��8$=	z����?�F��۷oǎ}g���|�Rڴi�m���3@kY�p>�(5YR@I=p� �y__������$�y:��^Z�v-��~=�x�)д�a%n�M��|�tTJU��r\@Cccpf����n�ԝu޹Їw��Ї�|�x�[n�0�����c ��d�t�gf
]�lv �5:::=:WUKc�E�{бЙ>��N�!��w��-h�_����~�ӷAk	yƅ���[���q�Zy^������3����H�Ri4����X(����HA��A���N׷p�F"��0���D�Q�3�aӾ�1���޹E�ptw���A�[/8�<�a�@�j�T����|�Ü����4��a��[n��\4wHE�g+:a���(%��.�	ot��%�������S׬�������P.o��3�R)tѽ3)av����@�85��Rj���<�n�����»G�	yX)�Y��
�1�m�q�ӈ�������V�L�x�$p���pN�ZQ	��|��,��k���u,���	�U^�7lx�2�ԆA�3%�+��"��Q�wA5({����/hյK��ܣ���ءZ���{ C�����m�&���X����8;D��ϡ2��D��g5nܸ�cW8t�g�̵���4[PuE�!�����SX�j�R�y��XBOc�>L�C�^ä/Q��q��'cv��0�Ҍ����<gpp
+}� �F�~�y UӜ"����7ƴ��b7:m�E����O�|�է����F�]��W-_�h�捏=�X��d���B��]�"�33c����iJ�;�f��(`a�]h��Y��;$�{�jE^�#Ch1�6�mKw����1�?�=_@{>���5�D�em�}�$�pxƕ���>Eq�	�y���*�K����.�2�ǭ���9���OZ@+�ا�62�8�Mq[Ϥ'���=O���8�f��\m����q���(��N�^;K|�С����J�҅܁�^d�KX���XJ�
}s����Ͻ���}��ٟ]�$-�-zQX�-�L�6m��
�u��Ǌ�c�1��N�,*���hYox���M����U�8�q��<���^h�bGc?�UY�OR��wI
;��3@Ɋf�nJ`��\����ĸ���x�q�rcɋE����@7�s�Ѫ!�AԄ@�=����>eMyH�'nذA5�\�F5��n����"�A7���SV�r�M��s}��@��uYUPR6<�̵�]�j�������R��{�z����I�ǰu�FFGg��[ThM`X��|x?rڷ�a���$��c̢h��m�8
���Þ7e�A�t%*�.�}��X�7Er[�5j�2��k62]i)#и�>�Ѐ���cJ��\���U���K�V�*9Q�-g-�V�O��%��神 ��4�p�1^�Ѷ��Z!cFB :��H�NAĤ��O�x,{
��SoĶ�V�͂JÙ*�F'cEܽ{������LF��z���04ר�ʅμ�Vc�)]��D�lʲ@	߳y�.i3��U�ڵ�dAͦJ�ZA-0�C�3ҫX����,.�(j2y'�@�c0� ��"��U��K����_d9\9�[%�x4�
��Ut�5�.��*��x>�j{��z���f*z��b�Ɓ�9�YU�òo1C+{u���Wd�s5�.�LWA���~�|�*����;t��=��:3��j�!�M�.#G'V��cY]p&��-ǔ瞰(ו��e]	{�ҹ0H�QNb
���-tL�Ad�z�V#XR��{0(3PB����N������^C-�%]4��̬S�x��q��¿Xp2*��(@��6l)���!Q��D�ި�����9�Ԉ�9��ʥ9��|j���q����H��y�|�rDAyׂ����(AϼbG�z��b��,L̊H?�P�(�Tb̍DB�����~��BgG�W�-է�j���,m���X��r$��Vg�����S�c�@���Z�
8y4Bqr ʚ��,�ЙN����jC�d���Z
ĝ�)�F �R���ȪLs/D�ʤI��a��!��L�D�2��7�$2r��1�H	r�[�<ݟ�ȓȽ�bꐤ�9���"dR䣞���lX��Z�j\�:�����Tx@3�R��nݙ�*k� K~�̎\�J.�lr|��$�^�&1�
ؓ��#�R($[R,br�'F0R2tA�K���ɃG�ڈ��	 Q���y��/��L��ob"E��.��
�?��GT#���'Ʌ�C'pN�T��=�z��Ck� *A��d�,Zd�BԬ����b� ���~��4,n�vҦ)`ᦪ�y���i�GlS��F��Pp��Xyn�ٟʫ� d�?2h�������fjf��)Y43��-�jO������5�S( �ݻ}��m���/�����O�Ƭ(�]ł��[G���3ي㧸4���]C�|����9W0b)��q)��~��Q4���I��Z�$���E67E��%{pDB�I���Ԩ���V#��l^�0�t��Qa�5G�Ϸ�(���pk>�'6�[�4���pcD	ԉ�*���v����� P�-kuo���T��0��x�ݏ	�8��?�2�;
aғB����E�����(�b����x7{�P���o�<�A��g�a���!JFfw���<@��w$&Ȗ'�����z��'��ʃW\q�G?�ѯ|�+_|�F��03xMz��غD ��	����0L���{�hE5t�&'j,~a��xq�����nu�/ѰJ*L�0ܲeL�E�I"��j>@H�`Ğ�X)��*@C�Z�J*���<�8�M��|��?�ѥW����)Dհ��:r9���|M���V_�r�T����ܹs;;;<X�4�R�犴���G?z�57F*[�j�=>��b"�$K� u�vn�?�qt�m͍Z4PU��ПhwT0t����zΜ�[)"��9S���;�n�h|	JLu6��h�v� Ō������ύ�B�)U#"��X�:H S.��)�/-/�9_U�JB��Q���� �,���p%�B1��	##�]߳gώ�[���{{;�`'T����������I+��&\��u���|!��f�p\�;����Ȣ��br�FY��t2 qs?kE����"��p���,X�o�>2N��;�����ppg\56:�C�x"%�cõ��r����P*Q*��b�G�rEǝ*===��� �4P�
�4�?ܹZ-�;����i��ױ�1��.����&ihԈ�]] s�����c�"�A#gJ��5%�^L�l''�����Ex��~d*WM�������Ӛ6�r�)@<�qǎpN^�
W�q�F&���Fc��-;���^*������SH��ӕ���u�k�fcz�'����.���]@���ð �*6�	�
��JcM��'�����"L�ʖ��
FF8 S}_�B��ix��j·���*C�t���0���V�ځ��H�A�S�
��lV�v�	|��Ք���93;��%�-I�4�H͈e:I>)��e�x��{E��˨�/��*А�����N��H4T\<>�3R&��D�J<B\E=���ɟ��̨�9k�Qp�H �AZ(п�+�,t�g2�L%���T����%<23
�3�:�0�p���vt
L��J�j����B2|\�1��L��c�R�0�9�8á�#�B��	-�R^�Ój�V�*|���Ďd��)(�B^X_�a�1�$�!�Z����7;��7��ayr�}��y\���I)�f�|'�Í7�|��\�UY���X��o�:���m᪡�{`tf:a]?��� 6W�^y�)��L��Gab�is��s(S9/�Vz���7��nh2�5q����������$�ɯ�QC�}��x�;�;6s���4�9춇�N� �3~a�ܡG��˥ɡ"�Z6�I�@)��F\��^q+ኃ�$9�x�c�8kEp�s������טn�%���B�Ǹ��V�c����Vɇ�\@x� B�f'�6O��S)���%��G��艒���������+������O~��0�u��$����/SJ�`#�d&����� ���Uc�X����Oy�;��g.��	|ùk��G{��z�۸�ĥ]��Ԭ1�&����\�.��#A�4�:����C'pc4�w_s����AQE߶U�i�	l#�{�u��0��%PD�zrh��[�6<�y��e*t���F�B �����.)}�	���э><�{�"�ߖ�Re)�mۖ�/��W�����N�d���}[=9r��U_Я$�Ij�8����L���FP���F5�.��U�w1��خ��� ��߮(4=s���Ύ��t�������4�gdz�Gd{��e���@�|�$oR�HR`"*X�,DAj"FYV�1�a-�Ю�T7+J���WMe!���ЩR��r)�\�����FOJבBM$I�����n���_~ѹ/_{�
ǵAY�� �07]��/up��������ix�7^�x`��M石�wڪ�Jʘ�?�{�y���@o�۷������iQ�N;�,��`y���<��c���۾( de�!�\Al�Js*m�	�R\�˕K�rʒ��r��Ri�+�IM�M�6�%˗/���'h�'�S�̤��g�}z���S������.�<�BN7Y��?�.�\����7���h�FW�TC/�F����7��w[���.��φ���#�U�3#Wk"�XX�L�\��Ū;���-� �E��Eg/X�dI�ܾ�ҌGn�H�!�X_����ԕ�s���{�����ГG<�t|O�S)1B���^��4��\t�Jd�Z�ܓ���tJ�b��ddr�]�����7�\��7��^'��ʬ�}������_6����3�-f#S#�v�F��g���u������'w�<�L�I�Ꮌp�m��~O��\�t"�n�1gΜ��������b�xB�>������i��Q���׾�5��*"���:hE9%��
f,-�ۓ-H�����OY�J�Ǟ�N8a�cOa淉}�E�J�<95�
�"l� -�U� ,_~�y��s|)E�Nun||����A���aM�<��&a�w]7L�@�>��������j-r�C�T5`�l�̓ua�a��r#�jz<��U^�W��J~��J���sK
�"M��Ke6bQ�B�z����/j��lUJek~$z�TuFS���r��7m(r�(t%�ӥz����KB%�0P��MDJ�ZҲ�ЧB�A����x�<`}�$#�иg�2Ck��0����n!�	&1b�$�`Ll�������a���1^ZK�h
A�e�+ر�+Mcd2V3Uδ(�4�ʼ�L�x�rc���U&'F���KO�@ˋ�ж��:�{/��T�yǞ���g`�v����NMt)�����*$慢c�i�Wf��Yh~���]8g��gw8vm߾}[��R�ZV��~;�~���}�^���۶�*OO�[]�2���pɭ
��bg>�K1��Q� Y jܲt�J�����ј��_[�E�s������9��{��qS����n)"-��ά���X~���9j��A�N����5�byYbR\�$�Ӓ���"����BԘ�	�X�K�j�S�_�\�n�8���_c���l]o�g���Ҽ�E�B{����l�A[���ɋ1gH�X�0����aŶ&��G}C��I��o��b���Lu���߄�����֑�0���Xk�\v�e��y����+�s=�-pm����B2e�@�g���)��ST��")��S�3MY��?��<���?����89� �	N�13��N:�G��`���F��͗BZ����Ȁ��\!��rΪ��<���9��'�Y��n�~�ڵ{&�f���CM�`�@V�p��8B���U�xE)��eyW]u�5�^7��W��񩷾�m?���_�����2ڀ��L}���L�c���k������m</B���T%�;6l8x�!���݃�}��C�) i�S�M��K�ꈔ0�y�EU1�>���iQ��ᡨ�Q$:7�sLQF"I�CP�''�O�C[~!D#�=����Y�����NLc���^�Lq��B*�iQM��b�hYu聞��5k�x���
�
B�=��BA�է�~�<�5����� �m[7>�KV�Xw��O�����Ff����V�~���{)��B��`
�"�wZ�40\�	�x�o c�*@b�N�7�ɪ�0�q"���GMS��}�׋[��5�p�����ŋ�9��o�2fLٶn`B��L o�v�����|'\=m��&A�ᒑ���ga��)tNLL0� ��~N���B�-��WHY	�v�B3�޹s���p�M�`09qx�/��p���,*����R-4qfC����q��3'_100�p�tw�7:MLҡ�=���*gT�Z ��|6U����%�=�\��߿oiHez޼y)�Hu�NXt��EJ�^�� �c�TOOgW/�~ >��;��X��F~N�17=Z���W�*�����r��S�F����r��3oW����� e���o������O�*��݈��LK�l��ڏ.������U���9����:}���	������Z>�)J��V�ĭ�I�=�zM1u�H)�iDb��@Q���V�0c&g�7���%��0(v�O���%n� ��]��$H�1I�b�z��4��ׄ�R�����<����%H�2�E��|$$��5֊��Rj�9�S�w�)+����F:'g#?1�����#�}D�o!��%� 8�U�|�Hp	�RX�0��ΝH&�����?v�ձZX��LG�q
Kc�+W��-x5�nR�=.sp�U+HsBuà����=�p�A����}��G����0���C�g��gn�g�Im���Δ��#�Mf]�2�̨���C���q�;E8���Sa�?��m^��֚0Ǿ��o[�2k��;���lF�K.�k�ݻuL3w�۝Z	i!��jϏj?�xcA%��gvU�G���D/�VE����h�W�q�MSu������%��3�L���w>�jI>����^���x	k������e�6U����{�?����x�;"&7l4]Pg�/_ȡ���*���$Y����|�`c���t1�Du�c������G,�����L0�9����h��52<?X�d��������^�Z�8`n�_��w��;��.wZX~�:צ�0��������W�)6�ɸ��Ǽ2Y
a��K���Hk��r��'���+.�|OR���0�[��C�ԁ��'�ڠ�腁������Oj�4X��k�x�|��G~����t��t+ˏؠ��Q z��X�5Gh:����|���I��dT���HmB�y�"eć�U�k"v��iX��%�����ݽg|?C�%�FcI�Ss��|�j�L	dd���Xp�YΏ����c���D̢��7�">��8>��#r�$�IH̦�
���HG	C+������ׂn��a���P����
P���V@'�:l�v���=�F^r5�%������!P`0��A�T�6h_:�L�4]k�ض�����ȋ�}�Pw�LOM��O�V��5e|vvϞ=���=�x��@/u���ݶ�ڂ�i��ډ��x	�xN5l懺�"EH�>�-��/���B�o�u8���&���7�*��W;x�� xw��a�J�
h�\m)�~�(1Q�%�Ά5�r��� �ܵk׾}�V�r*�aǁaP�Y����|w�`W#
7n�&��SP�zsy�f���K	��7�k#m�Z�����jT�(|����<��\.�7ch�6<����\3Vz@�1������ϡ'�H��G+>�s[2\A�]���"�zG(�:S��A\Ǵ�E-,V�)�*�9�A����Z=K�Y����IP�ry�8z���T-Sr���w,22�����Y�.T`_�7}�?��ӽ����i76�.h���\����)��Q�-��<.'d�TM�)����s�3S��o?�	xh��~ǏW�Z�{Aq�T��0`�
���QO(7�h��R&fV�:8�Y�����ņ:S� ����5g��YSb�5{��V{�(ٰ�����)U$�y�~}��&���T�px!#T|�q�Ȯ�Al�d��ߣ�,�Yc׻p}���4����7�	�i%!��� C8/l�kI�?�ʆH�FS� 0�yJ � �
`t���-[�#0
���FN� ��q��׾6��1[s@d�!��M�*ꂮ) |C�m��UEJ��Ұf� �Df)L��~�	DT���`���5��\8C��H�@�l!Z�1�*D^C!�lYI24P�`�A[�,�����cMB�̂~G��t���n��J�������Ɏ�s'J3�i�0�D�G��α`S#�z��"`�ݞ2|��o#6Ӧ�j�mO�j�L*�If�N8ᄡ�X?�.y��l�\Mg2u�r��0�}�T�����wN9�v�ݳnݺ�O=��Zj���L�|'�k5)ߕ�;г�;��&��jÑ$�Q���<q��u��_��Y��[,����̌eY7pkU�L�S�:]�vuu����#
�-{�NE�� d����H"���=�tA��ҽ�����K+q'eOqWV�EO;JOi���þk�`Ga-�q�Ck�����Q{yV��y  ���}j�!��8>4��{��#x��2Y�I?�=%n?���u��Oڃ9��������z�N��C=���u-Ϛ=�,�1�����0��78��ؼ����<�.��aȭD�㹪�u�#.���d�8W^�KX����-Ȉ�N?��׿�������7Z��c�ʕ����|���/����b�����0����5;;����|>-�rH���?h?;|}
X��C?2t���e˖�7<��ڵk#r�����]�f��؉���������ܗ�4�b��#j�c�=s=E���2��O�+��ϟ?q��w�\��y�:VD>� �|������d���.15t#�aUY	q�f��h͚5��w�2����.#�[��]���FLw�T3���s	F�����M7��(��{�(��c	5����r�#^�5�˫�5A��4ٰ�%���m��9E�>�fO�c�PMT���gNfX*;�E�8�t*���;�,��(ޓ�4��:�-g�\��H��
���x����ES�ip	�C��&�R�2�ر�qh��i ,U��C��x?�� ��Lŉ<l�B/Eq��z�{�C#�_��x<!ui�C#b�0���FGG�^ ���xN�Qk�
����g�ʧ�yY[�/QM��X"�A��%===�K�c r5��0���'�|z����üĎP�az��e��7�\��T�3��
2RRՔhR��[�r\՘����u䐚��9`�i�9>�c'�+�S��3^v)��������jc�A�����z��3'��r9������~ZP�5�%��KӬ����CbD���y�%(by� R�T�4R��<�ϳlP���t�Y��>�sr�廱�4e��N-x�H��#p�}B_p��� 4>�v`�C��B�^A�IH�֘|�I�p�u��+-�ԈC�R�gb𡪦1*8�9^.��쥦���&�"��[!���EB 9��	�1�x�84/�8��>���2���<��ͨkxdsDg�t/Si&��M0t�uڻw/�S�S�a>��|����Ϝ���:��G����V�W�&�x�X�B	E@`xB́"U���*�ե�dF;Etȯ�����4-X$lTt���6����K�p.d4�I-��3ZX�蘞��i>�~��g8�=MN8�'�xcYAd+�H�E� ���.���#y�4>`��O�V��Γ�`&��ʳ�xULX��	յ@��p.:��T:�ӌ�ꦵ�j�{��%�O��Q�P.�`ΤU\���\P!/͌q��5%�*b��!;e*���-�8��Jj��l�B�T �7爋��ߎl�Q1�G��	D�PP��=�?��ݞ�$$3�x��W_;��G�x�nU�G��"j��>���y�a��v#��ټK�p��~������
��J�6u̓yz?G\\������6/��?(�V�1< v�W �1�75������>���	@9�|�fp�u������n��K��<Xv9���؇FF'o�ĭ�l:��[����K�$�m1Z!�3�i�lsOse�Z�y)��7&s��51�$���!q����1�
����
3@{�J��A=���^���������U˗]��D,j���|�Y��h��O�]K���"�#�B�Ś"�1C�	I�@t)�?v=��ҋ$�o~�U�����y�k_	�N�2�J��؛���壟Qu�}�QX䕖->��{��?,�cQ�$up��η�:�8���� �R
��`2�ɢ��(�"��@�����}�M�-����?8Ol�n�"�F� ��؍D��d>Y���!�:%r�-%�"�&�+O9	���݅3#͘��)b�Pvw�ȇ�b��T$�ª$�J[�Sm��(�'""3�����mTѱA���,�3j0��^G �zW�b d����E�
*�[�V�+��TU��-���Qoؠ}�9�s�M�h]��*����PL��؋��SDQ�Q�Y�	�R(������|�0R� FF��d�Νk�*������P��ς"4#�vt)d���+dF�1� ���<c~��P���\���0ÃG��uD����킸|Z�HU,X0�O.G��j�3n۶���8�=#�;ȴ�f�6�An�2��^��RM������#__ωo�����rkN=E+v��r�
�٥cզ_��3�y3��a��Zev׮�������nݺU��˗��baO�����H�B���B}�ϡ�8L�B+�����Ó����h���X3*Z25��40B���Z:��T��/v)ݝaOa���IR��`�Nz�+O<��)�D�Ddj��3<�ī����?H�l�E^:����㳳Ksx/�1���LiR��-�*i��~G�z�Y���bO7�s%SF ��g#:x��Ι��5��;���w�g����ff�e}t	u,Ax>�}�*�L��Ɯ�[a^V]@s��3#Z�Z�t�6I�`N�x4N9`D� ��`}&�KV	\%�ugz�Q`���<FS�%]1�1�;*��dx���pHq����i��M
�ļ�F9x�L��u��=["`@1�
y߱�N�*����J���&" 0R���]�2&ʇ�K0�3�PU�XL�̉�F6�Ũ˼WQ��eAF;�5������U�s5�jف���R�LcBk����R�4l���0y�PQD��V�8��<aK����|�O�Q�z>W�z�/���ɪV��3�Y4-��յ�kG�+SL����m�&06/W�4�#[݊c1M1#`M��H$��+��hn�
ac�<�(�aא`�7�cQ`���@�ҝ3�����N֋��t�k^�j�-�aZ����=�)������|�3��\��n���tQ���m�<EV��lU�WX��Ry4����S�ž��}�'�F�[ˤOZ}�SO=ՙ˯X����u�ٳ{ߩ���|�ܩ����驑��\�wqD$2R��M��R�� G���A�rr�OB�V	B"Ŵ[*6S�'=������6�4�Op;������i��!�qs&_�0��V���=�uuE��&�5T�h�e	�8E��.@�`A$e!	�%*$�"�j�'+�%�a��$u����a�%��λ+��X˘� ��	-�$P6�� ��5t�$��4����}r�P����*|1���7���@��GD6jJEO(S�4�He�
���Z�Ɓt�[E�^�r�[6�8���I�����.�k#����b��>�wO��_���c�^T�TiT��aI7���9s�\��_��XT�#�%�d��7���_���bq�###P��������/s��W_�t�C�D^���|r[	����W�O��K��^N?�[{�/��>��g�	[E	�3�ɶ��H� ����1PDrP�5t4%2׹뮻־�"x����m�N#���֪U=y�J�㮘h�}�$�h��t܎&i�ي�U���A�{��N;�M�]��|�g>�D�Pn��3���)���w�[(�����_v�e��O_��������|M�@������0��Y�B3"�q1�X�0T=��𵚘�@�ZL��3��`GBԌ��|B;+W��k��g@w�'vqtM���3y�
�̦`1��a�}�$��)#5===44��zњ0h+�2͒����Cبa0��^��G�%���ryr���!��9�6`&wuu�s�(��s��GG>*"0H�o�{ �:;;�>h�Tqr���O?�o�C�Z��/�0�/�y�Lsi43Ż�'�.xG���6�f�3�Qb�iМ��8gT�v78d�m��h_V��
��AINf�:�i�����!W(:�j(��~633�@/K�L:b��7]������y.�O/��^U��H����	p��6���8vܓ{rCbLl���8$v�sO�@�$.$�1Ŧ�APC]�[u�������YKKB����'��1����k͚��������׋z�J��uu-Y�D��IӓS��L{,;;��iݰ��V,�fd������!�27���իW/����UN��[1�IP���&^�1�� "��T:�6���2T��+�T��'r��x͖eK���D�o������95�(&�8��QU7,�m@|��E*��8���t��SGBL�� ��?:J��y��7���v�㚩���s�]�=�� ���Ĉ�xU�*F�]]��Ks���R���!�����O7&��b� �$�I�4�\�֪��:��a����-�됁=��C*-<I��x�XI!���K!��H2b�<o�)k#���)JksQ�h�3y�z"�����&-�*R�?w��.�X+F�c-<?���Ｉ����Q�M��L�k�q��"%�ۄ� �LC�E�Y�/rY�}Dv�Xx�@�C�c��?!�)�b�5�qw���V��������\�5l���ץ��Epy�ܳ��3ܦ&@Ŷ�p<409j3�'<�6b�d7C1U���}�oOr>Y��K��פ7���������N�0�.���I�^���E'�
��«�=�ݍ<C��[�.6A���g�#�Y>9+j����^��)>\��
�^�-[���e}��^z��yD{z:��+��bll���ee��WبIR��*m�ؑ4�z�Lr�6�%r���xw	�ѐ�YNvq�f�BR�ZM��3��"t�b����0i�2� �ES0l���:LD�O��t���8��_��-B�'՗NaP|��r��!:y_\iaE�����n~k�N�x�[���@n���t�:od�S�����O.A����^�-**ZOAA�l��c<3�� Z����}J)�������.��WN��N]�mU"�d�xW�Z������Pv�����Z?�-�|�$r�%X2�c�#����O���e��XV����5~��#�<���]�ZR���"k�O>����=����r�14K��g+����dʨ5i��D#��
����D����725˩����ft�.����i���?#f��� �$$]�v�Y{�E�>�h��v��&d:���T����O�z�ퟏ#\OٰCI��!��v��A~�b�wV���<)d����s~���W�����ݬ�0�~˪�JB�.>󧷾康���q� �����{��_����~+�p��.V._w�ܝ�A��_t��x�P�XX"�.BDT�j��{�!��O+Z�4��4ꍄSQ�9D���	�&�XҘ��|�7�Af6�C����ޡ����"�Z�%5仪��t-gê�<!잮�^�#/�U|�Ы���TD���˖b'UQ�'�p&ĥ^q�C��w� �]�8DxvvNH��K�7ܽ{�fe�̔� W˖-���� f��1��Jh��@3�twv-Y��)W�gf1w*��`]��ѓu���Ӎ��J�ٰ裇�� g�Y-Qz���P���$�q� �q��޽�D�c>b�U�]��B6@t�`�0;(0b�[�c ���ʼ[Ir�÷�ɕq��f��a��\�t)��H5QsxgA �Ո$1`KB����l#59����n�\9���X��Ks#��6-��7��.<g��_��̙�����337���(�N��v'R5`~6/e~y���=�Y)p�Yu�����ڶs�֭�v�;���L��BI�@�@��P��HI�e$���"��,�bv7P�8�љN��궮�Hނ�U�]x�UWU�ϒ��F�U�y��	E.I�|z:��<B��crW6��w��)UpD_'�)����ƍ3��"�*���!i¬����#��^l�P8�MbKk��0#��?s��׼9��o��7�v�ڵ��mW��{5� ��(XN�k����� �i��U�W-zr������	Q��[�םW��Z� �����n���E�c+�nk��ҿ �b��� �2t��ˎ�2�4?��N >���KH'��_�]s\l�!S�[��`8�t2�9-r�qj�/l��W��*U�cr�8��~R�!�M�ҫl&��Fdy�8<��g[Ϸ�|>{F{��=��<9��H+N'.f[<D
���G_��p|2�2NsvFVhH�=����V��PuIG�>Ӏ;ǫK4*KcD�����rUk
h*��ʲ��y��p+ c��Q����܇o�	�/�A������y晕�;��3��<�����aS?��uI�>�\Ӱ_?һjټy�8�z��}Ua

��&��h�xRb��B��6�S��Dzԋ|]75n�S��W��~�᩽�Y+���I^1��"
<P�,Y��H58��`�l�G�,ċ��mz2[�Ȟd�Zc��=�~T/V�ek)� ��v�'���j^����u������@w,[O2<��[�����խU���?8|��3��G�T�|�5oZ�f����ߞ[W�tϞ=ɱqx���4K�pg���fs�^�:����BF�b#+,������Ph�b�
�1�Ĝn��Bu�Xi3���&�B_=C���0*Nա<���^�`Y��ګ�j@� ;|I��H�I��U��`�{OdE� F�[��F0X��V:1k���YL8����&�\t�=�,/�]�z6�1F�[s���dl�Nb��Y̡Ӟ�x�g�q<O�k��:������*e�"����Υ�
��U�Ñ��.��s��[cժUO>�c�pb�46o�|�������}�q{Ƃ�������{��C�п��7n��&����r��᫮�
ܝw������|�xUV�g���_9����^�h��d���p�`���E���O~�O���F�8�w�w��/���+q��*B?���x�	S�0*a�ď}5�r����3ar��4��E&��l}��9'��O$��~?�$�o�P#���7ه�J��d�0����u��ֵ�I~�%&L`T*5ƫ�_E^e���g�����eQ�+�p���g>���S�
��Бܜ)�)�w��VD�8��@��|��a�|��_��?��S*����+/z���SP�;�\�c�a���w�ɇ�B7y�ۮ��wv*>(6���0&� s2OW��Wm�,�}���o��Ե�f�Q%n	%�3�
��O)�B�/���)Ŗ-[FFF@� �C�?�*�w[s���>����ö@�Ԯ�6� ��� B+�	 �� ��CM=�=��U)9�������z:�g��p��H���`���U޵�Z�6000;�v33�����Q��h���S�c�y��/HQ 2�˶�9a_�]LQV�	w�q���"JV����$}pSpwBS���}¥����ARf�@	G��1����.0#�h� �@�$3}v�3�i�591w+��E�~��^^��~�;Z��\�8�2�S�62�h�P�V�4��H$R�1�}z�O�����ݽ8?W�:���!�@���9k�ym8?��;�����y �Cd�<xB�o~�g�c���V�vtN3�F2C�ǧ	.|JM��rg�ڵ��v<o�x!Py��oDu����W1����Bt��?�<���}G���h�Y����4jH��z��aX����)$���,���-�P���ū������tM�J�L#.I��O��]���+sU���3�E��Mjb����.�$d���7B��7�i�:��n�YsV�h�6�-�����uX�y��\�r��ց�8�)���!�^��*��!ǈ]����E��O]�L�Δ�BW�=Z*9~ �؁@��`�WL�n�B�$�AG�18�Af�v�#�$��/aS�K����"�j}�4��TM��(֪��0��,U�GoK��[�ϲ�����u��W^"p&6E��-�Z��]K�:���"d���$*Too4>�p�
Ir��"�+ ����5�Z�� Yj���8v�  Nm��M��s�����F&&AzǦ�A��!������n
����`���dɒuk/ ͹a������%,�7�ذ����:��?@��$3@ a�\ ����ĹL�����iQW�=~��r��=}\9lXз����HxX�A�Jˈ�0�
���j����5����'ا���N�W�OPP�ξ��z}�H���  ��IDAT��88~�8\�̙}���s�Ƨ����֝_|��K�$+�=� <j��4}�$�JN-YX�������G>�I���͇����+��m���|�~��_��7����61�Sq�-�}��_:o��?��O�d�LDnؖ�[^��K���w�ۿ���߾�c��%׽��{�}�(���.��ބV��\teqf������~����Cx����w����(I{�����v�[��U�7�F�F��j�xq���^LR��}?~�\s�_��y5\j ���B��F�+��s�R�*L�b@˴? '�k_�'‡�T���I�����S���LZ��y
>����;v���O�t�R�P�(�P:�!�5����l ��"���XӴ��A��(�>����?������B�_��m�����hJ�����}���@9 #)օ����}����{�aઉZh�F�%9�'Aݩ�N�c�j��Cき³�+&Ga�LF���k���ng�ƃ'$�,�F��ËM_�Y�b���L(��x�s9�����|4�^8���7]Q5����9� �c�A�bR�D�u�׹~M��ȋ#+���t�Z�Q�l���~����[�qŉ���3xS��u<ohh7�!��B�y8���8#�k_�����/��K,ya�^,�(��{uǰ2Z}�{��E`i�B{6��VN�2�9�h�a�����{>�a�c��'�j�҉6��H�U��2����8�����$�B������(�ÕO쪋d�!M�I�f��БUe�R4]3�(��I���Y%g��=�gvJa�W�Ñ��*f1��X�xqg[���fK/���Бc�,Ym&���M`MIt[��P$^NW�w岖S���ٙ)�3�ҟ��|��������m۾�g�)����Cm��榢��i�v�Y:^Iq{=�T������Y*�2�p��jczn�L4&�%�q�:�1Π
��r �"�C��mk�����c�>½�ݴY%Lv�"r*������I5�w?��,����Ny)i��?c,��O�O���DN}X���qDU�x�2�a���Fq�NgG��&]r�N]�:�N����<wfv2���;Vf���Q��1�{����J˗�X��YX�`1��t�x��}��]�ޱ45S���B�t'�oz�0�4���m{aO?��%m�Έy2a+���po�[�+��%[��q�1������Ƞ=6�9b������iC�MY�*|�;�>؞�O�����o�����σc���%���ā�1��u���֫>8�G]gG�v���A���zJs3Sy�"Ej`�dŪ9H�1WD������(as��[�5�vǊٞ-��ݏ=��8��lI��}�y�T�M�DN@Dd��*hǤ�!&��&S�9/X���+��Ҷ��~�c/�3�����_���#�wt7�g4�sI	�8)��	crlɔD��+;��qT� ���l��HW51Z�����9��yb �a5��f��h8l��i�q;��K'��'��&'�#
#L�G�$,�vh�ah�$�1弢�x9<��(�a���e�K��M��HZ,gtŭV�#�"9�����&qXwm���UcD�a,b��1����������<�쳠�E�m�ŋτ�9�MNb�-S�AP�.�b�D�0!���}{��$��ji����'&/��R�����������K��<����N8ߞ�1dK�a����^zf�f{��g��q\x��}tt4�x��tv;��f|�\ ��TB�0NS�7������C�\3Q뾴'k�-蝙QK�sh�5Q����V���s�Y��l��}GG�Q*����Z5`�O��AP�V�*���᭫�X�l�xuk�ĕx�NT�}'����L���3�E ��b-c�B[g�����J�&��5ؿcߞg7�/�捅�����0�a	�\�ĕ�W�V�s��ed$��碝'eDL��_��f'f��y֣�>��������|�+�v�u=�����n��|���߻{�+۷�>�@p�
�vp�>�T���j*bN��6m�:],wvTԳ�	���W��8WQ4!�����Wv �	�U,_�|�T�$iD�����;�%�ЧV���8�4�4���W��I��3��
�A�)iW�������~�1q3��a�B���7��?~���׿�4�x��g���/��_^s�%\pa��?�?o��O������:{TD��[>�/��߼���9�iM����J�2B��p�슺�ܘ�	�`���n`4��s��뎏�|��� �*~�NZ�t�6��YO@Y'H2�� ���jn@���u�ͬ�un�4��!��]E{��>�eL���59�Fa%�2�͛Aji:�.mN�5��H�L��,��/&-=Р�Zgf7�b��d��+��=&!��5�}�O��s/u�aDBK8�~ǲ[����⹮���DF���D�a�{І����J�r�>�GR�����Z)��eizRC�`�s�H(�EsÈ��C����,*/.V�'�Ȓ�F�"�ȁ���X��(Ō�赤m��U�,�Y�kc1E��7f�獅�X�O��%L1&�y�_��Vl�9��2��<O<�D5�J�������-�w�Yg��~@iz�"7�7�V:/������:x�ܮ�g��L�C="Ap��s��СC��՘��v��8{ﻯ��{��u7�pÒ�g;vL�ؑHk��4i'o�������!1�i�[�����w�=4�L�^�;I<�UƠ%���&�#"���G��;�N������irW�$���k�dԱ����6��)���#�5h�"B�a:q?~�9���;߿~������	TӁc����%���`�iV*��Ws����[֭[������<Q.��Z$����;��\r�y���;7�s�_�=������M�����,�ףV��/���]	��T
=�P7`��Y;ǎ��:4�v�50�p�"����?��Hۧ8x4�'���tq��N�B��8k;�������E����4����fgg}7���۷��`g��j�DL\|��h3VP���:�X��jTɓ`d�7-w�l�1^bAGqlvӦ=�Z}ފ+o���j���t�w
�Q5f�<i�k��s��Ͼ��7�� `����Q�� ���89MKaEKF���N�O�կ�8p�j�����<�!�:��EF�ǖ��i�R�^�%$�D(����N���ʪ7ߣ�����H(N����S�X�xꏘ�́j4��(�,Un��A���I:8uooo;YS �VWju��ᠺ�gsp��,��_q��g�y��Ú8."B�B�eӦ]�v޻�o(t�0QԺa�����|I�8W�ȑU�Və,�ڰa���	�+싹bqffn�m��E���B��B�=����M�ю�)�i�jEp�E�!0��:e&ki)����Ҡfa������~��###��H~l��Yguv�[�n����{����%�>tW��(Z�듁��)')ڶm��/�^���W`CUQo����p��y�7�t��GpVX{;\ �q܏�,7�i��[���������A���J �9�(i��`4���'�����Q�X�q�S[|�����o4Hq$s�o�����/~���s��ŋ�=��c��r���9B3��_~����7����Ç�[�]2��7m�_O�+�x�ڵ�?�܏~�����F���^FǢV"8�h`� <Κ&�MЁ+W�ܴi�D�5�xUE�O��y��M��r��o�m��e�?�����������6�W	u��;�7�xh��aU�L͓����6��ަ�6���A�&�X1�o}� {T�Ûٰ᲻�����!�-
��駟����+�������������/|!R�/��������6Z�ұ(	�ǂE�<5��YM�a�	�����~hx�S����>�9�WY����"�߬㷱��94�p�аp{T�l"&SH��GS��!�q� K�\.�ƨ#�c��ʂ��=��$Tc������&j 9�|��iE�2�U4�X�A�+�*~�_�?1R���i���i��_��p�V���it�qU �ݲ �D))�Ov�r��0�9\iT�����qh���	NG����H4X�85%�,ҘT��H҉^���=�0�.)F�BM' �Rq�;Ԛ��}@�@(�>�&�.���P}Ǫ�����vl�-`Y�	d�$O� ��K!z����u�񢱻�l#l9N�4�"Q�J_A-r�ފ!(���R7��BbV����g.i��si���ӕ�Z�dX�e���#{��p��!�S�)0d�:w��mٶ�˖ɒ��Oj�6YWB��߫�W�zq���U+��/���=�}�]�׮q���}x0�����n���l����͗_�eص�<iI�ZF���3&&����5gr�}��<#c��*��H��s��U%�go��6���1L-/i���{� �N}x��D'���K�Bl�o�4+Lc��
&~�XJNR�A"�=�	�E99��{�{ǓR��\���ո��x*�耯�v���&"��8L��Q�F�1',��q����x�QXv��6%>:}|f��ҳ�ß&�w��? g��1�o]{��Ҧ����<�F+�(����\��2q����dk���Ě�@0���ӕ�OidU7r!��i�k�o�Z���%��L�\9E�Jb��)"Y�H/.%syE�ok�eY��uSq�`�<>:��9:|B��|��*h����	�݇p$n�dS����r�ݟh��.�J\��,��'���X��%#��=���(��D5�
�*������M�>l��Z��+j��^�{�x.e��$�@�59^�w�V�z{e	���ģT.��S�w�%���EW���T���ZY���=�k�v��xp���	��꾖5z$�XF�A�A=�Z-�foUA���(c���ڲ��C�Fyk��m^�c5L�.�	u�'��ɉ!bmM��q=�)I)i��1N㚐l�z��kfľѝ͂c6`���\����?�'ݮ�
Ո#9L�}��~$��* �75
��n����������#�0:�p�R���k>��z� o
$(c�B�R�lƒJE�����m��ʷ�k������y��rF��f�V�GH����^������965y�޸��K�^v�:r�X{ow[O�bX�WՊ�|��ڝ֠��a&(
'��C����m��"�i�x�;��T$]�9��p�@��N�'e�h��:ɺa���	��#9~6kV氛1׹ԑ��_�!�[��b�EkK�#G�A|�h񲎎������P��}����;?�Vk�މ����-K:�컥�Y�ag���Gg�}��5�^w����B��5ˢЇs��?�3����z�%ú��wںm��A�@h����UkVò<��S}�Q�������m���>�zz�@t!&ԋȓ���o[c݆���l)O��`O���P@�@F>į1���|�'�?��}{�>��k�����/y��O<�c7��[�w�ޙ��O|�c�?��w�����vj�C���C�_�漥������-��W\��CG��������MDЌ�:���_:p���?��;�3_I[�����z�9�$�@���p=_o`=xڪ�:�
-YK���yȸh���Fc!��P�S�2�R�<��Kl�BǍ9�1�;)D�Kx���9�K�=��&!J-N��4\Jb^$d�J|�C��|?�u�^��_����C�ltk��I�]�V>����׾r�����|/�]�P�a�Ӵ�C(��&�A�HxN�x��y�k�����E?@���i�8~]����Z?�H���	��I����Z|M�q��h�h6C�d�����CB��<�	12�	˵J6��	�)�pp��A�<��T;�$����|�w#��k���s��'�I�e���޷RJ�'s���8�ɧ��(��(�C�ͲM��bK�\�eZ�a�������b(PT���.I��=K� ��5�>}QB�t�j!(��*)�0m�sc�j�P�i��GLĉ��G��\UF1C���2Lp=}W���B�<?�
V�I�=�?{8/Z�0��ĕ4�R�E`�ʂ�N����l�N�`����<�yL�+u�joow}��3��DN���z����A�Y);pJ5ܖ"��Yֳ��*>����2�S,���d1�ַ,na�Ν��C����:��(&��s��tt���֎9�3�jy�|m��(�F��j��rmmmLx�,��Y$����O���u�zq�\��h��Z�ڔF�2s�$ZV�w�	[3��
Ok�XYS�K�A�,:5R��NP��N�c�|���E`x��LMM�,�Ai*� �=bZ�Z&#���6 ,΢E��z��ѣ�y�B9�����.]�����H����|����
&��`L�W"|��#�.VlB?�l�˂�0��1�I�"���gR�G�`=*K�R�I����'u���L&''�cYNO�C �cke6��"N4n<��Q��K�vGBW�?���2�͞[��y���
}�eX^�8�y��1a^���x�X��PO��	�ϟ??o
�W���:	�|�������]$�.�e��p��3Z��GK
B����o���ji\P_.\9������R�2i��xIZ�D5N,j��8C��~U��� ��r��X�UCµ�ӑ��s=1yt��vQ%I35�r�hָ^K/��;?hUr��o��FJ5UWB�m�~6�I?U�@���=���ī_�^��w͜��cE�F�K���UXOx�8���gmb�ɾ���(ڽ{�����?���:>���AD*��,�&�Au��kŉ�[D��<��R	$��- �y��D�}��ǅ�.e��1̀�={��t~���\b|��pBl�M�msm�FX"'�k�Wq�s+%�a.�������Ç~4���{׮][�΁�wta`��`�����o�~��q����(�l�M�3l�������������իW_t�EN�
�G�2�Bؿ��C��w�}p���lG&'��I���gx����7���{��m��O~b��Ű\��ē6;ܚ�����%,�x.(��q�'���E��Dx���,Y���?�>��O>~���U�����x .b�s�=���>����;�ݵ�^kk4�.�<��{�R��0�����-K�ꪫ��.�;�f��v.Ar�:\IY�c*�H��o�<��vc��!�_8j�d��i�%�u�8�U�X0�&�� l�'awEn0�%(#G_�A��b�d�a?����y�{?��\��'��-�286b��k�hA��S��Q�y��\\.�뾛0�>	F�PFܽLW�����T����z衷���w�}76��F��� ~S�_�X+����Xr�pd�+���0�LsD@�|	g:X�,$�蠌a(L��-��[���!8��jhHG������3$v�hK��(X��C5�E7���cf���I"��0�4���*�C����%�l��
��(%b�h}����Ywf�AM��1�½���P��T�B9	��`so�F@؏Ќa.���6%2��B������BQ&nnxz �M3����?� ���	��BɆ3�B5n��V\W�lUA>uŊ��Q#x�G�2�CV1����
8�b��j"TٔBW�`[a"��R�)'�+�"�ݖ㋺!�#u�ZH()���c�pHT��e%��\�
�m*J��������d��ڌ�&�"��[����F.��#CS�����5��#kȈ;��%��u0r�\��"z
�mfnhh(��8djb<ȑ�3���u!�	r9��3���j��:+�1%LL�%
���! ����ùdep�'���E�n*!�(�����蓱�i���]���=oZ:q���1��.+�FҢ�8���j)H�m�l������m$PM�n�.UC�O'�n�u��c�v������p�%kH��A��z�#O�����1�N�W��`=֒�`โP8��TQ!%L��7���D��)"_q.��y����Cc[�f٘��~�H�0���j.�R�&��*����qHSvb�sQz�߾��*�5W�9�7�Iql�7�>�o��;K�*x��d�J�Ӵ����|��7b�(��wo� r��6�N�����|�`����G���8Xɑ�P����j�	x�����I�/�CkGiTC7c+�AŽD�(M(�b�|W.����=nٟ�6�����8 ,�`�;��&�bŕ=��Zqd�l��z�ǎ�Uˆ_��=�y���ph$p�X,תg���^�[�������� řH9I��Q���Z����7��^~t[^�^�ƥ��GFJ�'*�S��==e�=t�X��:�E��삀v��~X�M���p����ao����;��\���A&;�.��U�e	 �&����E �#K(�X�|c'U�仪T�U<���@�A�A�(�H�h���D	|�n<q�A�o	$9:[����8m�6yj�_��!c~DDԚ�+ئ��C��G/)��%�~�����P�h�/���j���V(�+�6u�Ȩ�Z��rU'�J9�\Y�Er=Ƃ@�֨����O_�������֪��a���-R�N͐�p�))����x�2
	��#C�+k�=m3�{��M[��۷odj��%-�y{w���ͷ�
�D�����z��:0���z_{.�{��+-4�A6�B&U���� -$c��p�����<��.��DӇs8� �!��9TK���	�~|�w�o���ׂ��d�m��0�]۷?��� ��������-&&qCAX,�bvC(�]!H)m]�`�����m������oxCOgn������?>6��/��}xrrrj�k�YL��3D6�KTK�]Т9U�;>R��]һ`q��O��V���Le׶ˣ�zq.oB��;��;�$�$ܶ`�t �]%)#+�k��5S�
�����(��x���yX/	"��Ȯ"^9>�ad'��|��������p�9�ׂ6=:y���~�?��d�o��=7�|��]� v�~���8gՊ��ł+�]fr�[���C�?��G�]�G	�n?~���]~ݼ�~�<F������c��.]�䜳�q�d͚5?޸��k	7Lw(B&�ͬ"g���?r�Dc�C�2��F;_(C�O��fQi�W8<KԀ�q�6�ɚ$.�t7(a�/�|_䋴�&�P�����\�:�����������|�c���~��J��G���K��F������۾��s��DͨA��u��P�`ʡ@vUOO�D"Er$	6YwEu�~HPVC/R�l���[?�����������؉�l\���u��%E9�O��Y5�R�_�����D� #1Ii=<b�4b��o����Ks��4�}�$�Z9}f�q�1�32����*��F�<��hv⡳�EF&h�jRI7͸�F(�4A��M����UC�L�r�8���/�)I�u7I��{_���O�� ��B�m��S4��2�<��U���nO�K���v��r�K�| ��(|$��ڄ͑2��i�_�8\�$T��&��}(�Db�5�3F�^��V@k��h|�̎ �+6�?-��QGt�5�#�pZϫb'���b�=gr1Kn�3��!	���L+T�S5�����V��� ����m]�B!8|�ل�JYS%§�Xa�\jٯ���E��m���)�;g�B�-�\��椚Nf��9�9�R�����@�0<<�����"J�qQN��db	qhT��:0�}�YzT���Ö��Xݢ��B&�d��`c���e�h�J�1��)��t��u��i�w���y'"����Tw������L��|iq�L�L�N�5�"�w]&�fnC��j>�	�f��}||9�h�C�u#��)2�̶���
-B�W�4H�8W�ynW���:y��a�GU���1��԰�a����2pU��[D��"���e��<k�I�ZQ�adt$d�2c��s�_GTiX�s���vV\�ý�h�r�gS9.f����2�g��剙Av�Z��s���E䎣Y=X���5�$	V�b���J��u�֑���l��fq���RǙi.HV]�\�/��1ͪ&�&8��>4�H��O��IHהh�OĆ�T47 5M�+����ձ֫S�'lP�'�)3w.�����G���%�� �şx+��P�����ɖ)4
RN��L�FZ��$�8�R#P��hc��X����4h;�C �D#�v���G���������j�V㔿X�:Wڛ�g8!�>�t��?��Y^�g���w���u��# ������8�0>)E4,�k�̮$8�#�*��Df���ls��K��hf ��?m۶���Ӊk��A|����,��jbf�D��j�nƍ�Y��4��k؉{���;�,xb ��V��۷��w���$vS�)^~�e6a{��Yy�9ȍ�V�;[�����æZ��I��h�W?��V7Z��Y� ����[}�߹��`/D4�33-~tbb�^��ϟ��X���?�����5hh(�5.��"uJDTj���K{���瞫ox3-�g�g}��7�k���D���=7��'>�����ξ�>�k�9�y��+��N���� ��M�v��rc�&5t�#M�&̈́Ͷ&V��>@�v6OQ�r)��,n��|:�Q$����6�����D��RMV�0W_}u-���g��?��`��&	�y��xE6��oY���˳,f��!�:٠}��UIe&XI|��_������}�{߽����&k��I��I(�7�����@�I�h:8&��a!k���%14/tif+��^��+Iх E�=|��/N9�i�&�ѳv��h�K�������R���)*Nװ3��L^�s��Ƙp�����֡�����<s�s�~�pe�q4C�	��R�ς�S�k�lD�-iD6 kv-�NH/�pRr@w�=���Pz4�Rc�B�4��
�@E�z3�Z%�6�a]ײD�o�6����j����4b`,"b���M$^��R���D�J� ��'_)r�~b���ErҜ��؋��ke�R�*H*F6�7U�O�
N���摍�38����U��d"{�`��sCՔ�Ilt�;b��>D�&k�����W���:���$�k�_*8�H`(�:h79���X�U-�ݗ��B�4ʎ�+�H�9��A*��0''f��ƢP	u�� ����AI��يR�������C���l�iF0w�a"���	5� A�,{�?61�oI84�D ��+!=p#����L�1,.�x{Ad,�=���B�2$�-$dK�����!�	xH�N�H������&�WԜ8L4�5�iQ²�25�A҆Hr�E\��q���H29I�u�ѧ�|6~D��w���qnI8g/Y��2Z�`/�}�v�K����vvfj2[���N:R�����/]�8����	i�ܖ�/�I��������n��$M��a���"j�A�,0i$�G�
-��!&\D2@��a�`�e+[FF��ƩQfћU���z5|
�����:댕&ȸ�v�;<6W�o�=r��/W�Ǽ��2'$'��7 �&9v|�"S:6�hs}��3�]`�qNƾ{�crbrɢs��#?:�G��e1>��ARO������μ�������}�ڵ��w��O�=����߱W��-�Wq���#EM,Z��×�[���,�ކ>h�
W�!���{t�Q��mo�p͉���_HY��2�{��E~|;L������(��/�̵,t2
��(�ݑ\����:��j��Z�|���BB=�*�^K3���;M�uB��ʛy\�����l���*���G��H���#�����o-&�L܃����A)*=A'��iH����f��eP;ut�q���~���<3+�j����W̻׼2�nn�ṏO���ձ�1N��~ �5V�`�O�.v��F���� `�Mถ�Ý�&&���:t�@��h�]�J��N8�[{q���cǆ_~[�����������ի����zh���k33w�y��O�f^�rew[Gmb�& ����3���0e#�{���af�M�t^6���f>�?���r������CK�Z�񥽂�  ��=r��	���	|������Zp*�bxnT�]����8��li׏~����mk� lrΩR�Ԇ�c0�qB0[��L"G��zn�<����o�B4���u�\�|P�Λ7o>D����d�����:����1�$E���?�{��aK46a�����O��S�H�X�7x����]���=֑��W]{�+{��_~�2�m[��\������1o�j:�l�x�c���/�s��~=���tᕗ::�uS�,Y�b��R$�����}��	]��O/����?�O�t'v�ł��P�w��5�[�MI��TU�~�8��"X���j��A>�=[�V�GǆXn@��t�4P!��Ԑ�%���L�4d~�0IMQĠm���4�.~�[o��<����KB1o��6]�]�(�ma�H�n�BI9L�<	��I�z./�ы�{P#~5��ơ�IP/�+#�[^��;7����b��~�;߹�ƫ�����B�&,&�7������R�i�V�(�BO�@�)Q"8���oi�zI��tdBzp�������a#V�\�z�Gܢ�$f����}�ʉ\C!�\��0	�㨔�K-���ȭI\�4����w2׼���-Dog5�8~��4�0�A�Ĥ��D����0�	��!A��ز�,�Cj�!��)y�MX��%b�O.q���q��9�R�$I'�;���;��d*�Vٸ��s����0��J�!U��B�\�f�i�(�����>zΦϢ�M"�A>���z9��𙓖���@�K�XA�n��	t������*[��''���">�й��4hX���j�H�2�;��d�ۆ+O�(o�����գs�����C�3"��g�R��8eˠ監�.F�jyS8�T���ȍ!�2҉z�ir%%l+-u���x�:�m,Dy��7��#&(#�Vp���R@dq�ᤖ�f|"5^���~���>��l��!�����T�c&�F�bG�*1g"�G�%�?�q��/�� ^�,2r��7�'�M���$�i>���IܬM%<C)I�L�L�8�F��y�M��U=�̄���F�\.��Lg �-T�2�q#b1P��^E�>Q�A�E)L�e��!�E�Nc��B��y^�2|V!l� H�y�-E���sR#�5����t�333�9���ƸjQPsM�"������j5~L�e���q�n9n0�֩4=`ۨB#|d�&�ii� �:d��I)c{� s	��)�0��8֒�ɭ������bI��%��sR|u꩒�f3��u���M��M����\~Üq�it�5)��P�lr���IX�^�jɂˉR[��Y�!��
�QsG�E�)p0eN�4)c��Y:4��\I�`�Y2nd�p���P����#�`��5���f6/������%�Fc�SQ���
���p7o�l��:����~���1OAR!'i�KXQ�̍&��h�s�3'e@���*��d���K2���DjnU.������ˢ�:S�	��Xx���Xi6M�c�O�H˕�F2���F�Z�tlqx?�ƧbV#Y�
�I�?��9	��Ei��.�ᆈ'��\���U���<b�Q4���O~�n�z�Ek�o�γ��$�+x�{�{�?�91:Z��/����?�a�etw�p�窫�z�G>���[w���ַ���ށ�]{��{�V�{�B��t*uC^x�׾��>��w�-��I�$��K'�ӯCs�4BҳunFM͹��5v}�/v��6�BY &I��O`1��<�9À��>�Q������<߽�~8�7>����r�-��.��'~�"ʲ��6�U��b�-���=����#���o��X�5,-aA�������m�y�o|ӆ?��?x`��+V�j�G��B��߈��>��n1�c�$�6�DlMh��DH��?�SO^�.��y*c2{!�H�t�=�X��B�ƭ0�W!�� �n�zssn�3��:FX6]`�{H�1��1�HV9!r�$MfJ�Z�ʝ<�f~�u@����f�uz�������"d[�����1��jz�x2�fpR*�X�?�R�J`M
���*k	��ä�f�1�J�0D�8iJ!4��i
�L͝�70�%cB�J�3�ΑlRc&�=�(2.*XC	.XָM�X�!O��|p��K��d]E@��c�$�<d�"��c�IU�t��(8��ØzN)k�6��X���d�����@ǔd�RC_g���^LEF�z5�e�H�5t;�����&ٌ.�e�wuh�X���#���I!)��8���ӌ2�j���l��,�,�#�0u��E��q�pi���#3������
�M���^�����j.	����[4@Ypd^�#��~?x~��e��/��$��M��RW$�{�^���Z5��]v6�>(��)�f�%"��%�K��C�Z���J?�$I�,8n
�B�R�مl�:ыΪ
�=�T��6(�O��J���Ra*��B�?ӃG�P�ZF���jc�-*:�4Qe*L����A�5��D��Xj�P�z���ZĖa b(���Uk�+;v���{zz��;2����X_W/�wUox�`www__��+����ׄ�k�vX���d?�����"��	�F!l��c䄽�����?�V�0\��'nڕ���c��ʏWf����kRl�%�K��#���|��n {a�H
I������:z:;;G�39]�moa�#��(a�Vpu�,/�]��X�paO�妦�wBYp++Μ?�u�R����'�3
����Aq~�F��5����Zvޟ*�����\��XHJ��wF��Xݶ�BNҍR�*����#a���,���ġF�=��n�o`�-c;�<���;wj|��M���J__�⃆L��A��@�E�"3��,tI�Up���h��{�Ȓ����1W=C꜑OVэ>���NR�鎴�}̠Q�J� G��H��J�K�Q�%%��NQ/�X[��礦��h4��vM���,�r�m�<��/V�7n���9��\a��	e@�c��TsL�9̡��
�b���?ѢE���D	�J�EBƱV�>c��3�+e�ڦA�aݱtDA�颤��������j��=�c&��)��`g�Y��q�x��;�ɡC8��d�ݰ3��,�T��c��b�4�3>�r3f�ҴFDK���4<�<����u������.0'N���uϯ�Ub����eFX��q6�����F2�re`�`��T��v��uϲ��A�Yi��]�j��m���}^�����(�p�����L�V�N�;�Ns��5-[��KYE/X�����<U�b�j)*�j���-�pI��Y�H"�B��_�ƻ�}��a��Hԟ��(�Z�N3E����X�
���ȡ������G�GrF�'~�\_qր껥����1Zt��X�erqm덺�q]�k���k�x�g�g}��k6o�96S����P	���0�"k��dE�$z�X�����x~&�PsJ�)���i��s�1����͝��쒲.!�8�@�㮤�I�<�͍ߌl�F�2�p���4ȁV��P�ӢU��`��A�u�f#���+V,okk������*�f&	\pI7l�lÆ�����R5�c���9ӏ=�����>4/D�O�>1uu�KJSǆ��z���AR�^w�8�M�AXbLF�� �Ԍ$��|�3X�W���[n�����;>������ժ��ڑ�+x/���
���oB��|*��n�'E���Z��$Mi�f-��X�BM*�8Kڛw�so�F���2�K��Z��'�|�c:�0��4bU��'�;\�a䯰�98`����N�_��4�)i�H��TMj�D_$Z۱�գ�~"@O��4d���O����ޑ��I^�Z%�ή�p��kQ@� n
�;|ICp�*�Hx&i_M��h���.��CQ�h ��*'_�|��R�K$ ��P(�v�!�_>|�����Ad��w�pp�>�K�`/']D&���Z��ϭ�
�k��f�dp:�������όOr͇��%�����`������0ݼ<�E�q��M4DU��
�����^,���9"ak��������;��ש�#s>�R�/�5�2���5fL����u�@�(�C�KI��M�kթK<	�V1�ǽp8r 'hє�n/`動�	>k�&ju@[��)��T茟��m�$R}��s�����E�4�		m��S�WI%V9�Z�	�|�`§���{!���`�Kݡ.C\�&�O)Q�g���e˖�l4��.�AQ�PN�ͦ��
W]�9{���N��:
��!�S��.�LI�Ć�,���jn�F�C�h`T��0KH��N$�Ra���#�֗J���+w$�Gc��s��v[�T�1��!��g"�/����NbO�^�ŷ��GR�r*���:�w�^� ��:y��

�)pJ~��d���qR|�ʪ�'���]�ȸD�+)�8	��P��8s����M����d\V���RJ��q*
�U��ӧ �S�B'M��>����r��F��Z�u�`�|��gfff�o���xru�K�9�Q�L~��:�>�]���Cv�Y�_�x�9��a�\�0�-�b,��J/��[�tމ�;��+����3b�lf0���Ax{���j��J\� cAe?5�i�PE���H���B`�)�T'.W"J���/NK�7o~�\f$�T������8���)%��rk>6@��o�HG�S<�������i �&;e�Y�N�E��*VP]��fL�Yd_L��ɩ�5�Y&į��>�Va�
����C	�$�l&��Lxk֬���صk�1���7Û�@+�\y啰���w߸�}��7��Ͷy=Q�ʢ��o������������\�j���_/ۄHG�	Q��NK��Tl��4���(&8������t���q����,E�B��nZ�4
:��oh���ؚ(�i=�ڒL��������Tr�RV��B��g�yf۶m�>�lq0۪�޽�r���'>����?�㎷����AX�	�������ǎ�Ͽ�,�)��؃�Q�*!e�1��E��F�h�M��8��z�Ν;|����=���=^eN��߼p��>���r�E�8D�4IèF���Ğ�h����G�	�V��f'ݗ�Ý\=b��!��XJ�� �l����}%7@\�yx�Ǽ�"�dLue�0F ��?"��Y[d�/��
�I�]�d��W��){�9V�徕*��;�G�?q���{��e+V-tk�v���2K��p�8ޚa�i}-�����Lj%�8Ԓ��7��DY����D�R�T�)�#�F��!>_"Ֆ�YT��Qh��e����J�O)M�G7B�I_1)��hX��)_J���=a;�a������D�4*yD���غ�j�T�c^|�y�֭9>v��w'ˋ-���߃'Rh��g���g�7\}@��a"���L�w]׿p!v�.%��]ٌU�=~|ǕW\z�@q�E�V:xdjʫ�=C��+a.ags��X�����09>>95;�L��߄�ʛ�;u�R�֫��A��+'��3Ǉfg�u��u�	(���[���ɜ���6�VuM±d`k"�Pm�F	��n����h�9�	��d�k��0�|p%��� ����>��E8M��������K�]|����Ypx���?|�ȱ���z�3����Gݹ{��W]�`�K3�_y�����mo_���k�.���ۼq#��:��x�cC�N8�q#4����;�Һ������{���`���U�0T������x�1!ל�s��c��{Or��fAP�M�P�����{��W{������f0�|�_�>�ݳ�Z��{�����M�x����5���+�O5ZМ��GV����1���\Cl�N�:�8�5��c�$DS�TS'�v9D(�$v��Ztuu�v������uS����Bul���U��/?���3Xdcu�Ɨ_�ك�:c���o��.��
7��2VR�eQSո���Ħ��1��O��`��U���ط抱FqF��P���.>��\��)�l�p
�Rq���Øqh�o�{s����f�8�Ӄ�"��c�,&�.ـ����5�7W���Z�fif��gX$��4�`�ĉ�A�����չ�������ϙrv���PC(�f��n�46��)fbu��X����aݭ����r��h"WCif��X�lfE�uYNsr�e-=묳^�8 �ڮR�Y�A<����*J�]�����?Е���_��X�i��p����� ~��� �}���2읆�}�$��*�Pd�*�����7m&��K�O4%�lgH�P� �k�"�m_K!��N�ؒ�&�q�`�<�%�=O�aR"�9��E��8�i���*�����V�KnR���(�N놲���\��,y�bJX"�z��U̖X���3�Ȗ+5V+WJe�e%J$�Dy�e��Ǳ���rKA�@�DL��_�i���7o`�hR�i��3�(�ɫ4�r5���ޢ�%~�kڒ�[���f,����%��󍅪W�c�X��)�O&���dJts�+����<���9�X��D!��	���띙�G0� ��F�c�z�sǫ�Hpɿ�2�l`,s��jX6�E>˶��u��(���$�g[8D٤ٮ��G)�硇ܕG����`���(	�F�۝t4��i�uYOV/�i�!pL�p�z��c#:��������?2����-�-�R�T��� ��&/����:���?���_kT��h8v�*P�lRE����3�6�1���ы
�9�<�A�>�݋EFJ���c����x����W\!a˪�'�Xfv
	gth��矗U��ma�g�K�,7m#F�0�&(�8-R*�Gyr�1�4׷'-�ZX섈��p�~�pX���zu�gl�q��+�HAlp{�Y���؎빗]v�C=j��/��a�CCK���7ހ�))<v��O\y����w���O>�䙧���Xir�-��������o��&�4�!N)F�X�*I]SU�`��7��@(�Դ�7��z��S��C�z�K.�Q���J��;_�z_��� b�*���0��u���F��j�X�	S��S�0��Q$��Vė�w��޾�mO�ڐ��(��5U��F�{�I[,8f�ff���!�����/��p���H��_�ЗI8��l9jq6�sDG��k�Gn�ƛb���m�q+��J�F��iI�i7��j*$���HT�Ϙ��ס�s���IZ�I�:���|K��GF�j'EF[��-
�����)K���}A"���H\螞P��*�-N��<<<��(��M%��F&_@�$7�.�M�6͸uI��Z�۠�h�| �_�c�׊�">F�"�˂j��P���0'����"��M��'������@d�$pg,�LA��wu!�;86\���W�a= ����҈Y�p7�b```�ҥ�ET,W�l��\�e�w�rY�2�{� ���:�c�>����U���c�{,����#���B�#\
��z�j�ܘ�����h�#�׎���ɱ�f��cb�R�k��l�0��E�0cN*�'�5j��Bn�(U�g�	U�
V�Looo���|���:��OLL�t�#�4��ǁ��ǚ�#[�1�������$����s��[�qw�s��`,\�|����"�l�v�(�Z	S �.-}6�Z0
q����"b R�N�K� �)l���Gi�8����]��^<��p�ʬ�M��3]��z�����ǑH��b��QV�d��̔z�T��v��v�ۏ-[��؉1�כ�`ܪ��g~�z+R��
�E�mxW�+����I){VT��g���8m��U���t��^�#k��DP+7E��t2�V��� %EEk�ܪHڑ�)##F"�T�r�������?�4Ͷ@8��Y\�(ta�wes�[�Y4u�Uu�s9��"��/���b�����h�.�'�#$-\(��:�j3�پQL�M?h�^��My�L>�eSA"ܣ����5�gی��s��2-�Ky|�0�+lpp�s6��'���s#X(�ed`B̈́^� R��s@.�C�:���l0�)�����`�@3x 6��bmO[>��7�p�P�؏<*^������!�ycI�̛�UuUQ-���5�?�-��A�;�^x�}��N���?��Y!+��׹��+|��W�w~���-���I�b�y�T�����f3�'<x��/�}[����4�\��^��o|�{��Ki����۷�K�����+j��j�*��/��w΃UH����(^��Y�p����~~��EU�[���TZ�s-1�.�i�k��h��a���m޼����߯����J��6�� �h���X�I�)�����v�z��Ͼ�����3I���� �q���o^s�5�/��J��jhL�q�w7l����	�=(H��`�|������n�������[]=���������8�j�'���z�Ga�ၐ��>p�/�QV� �e�Rq�e�q�}�A�6gv�=?�ލ7��0�Br-�$���t�E�s���S)�p���Ο��爈Kv�< 6T0\~�U=�o���?�ٿ�ӂy*�EI*���СC�#�"~�6�����~�S��_گ���� iY`o�!�:R��ou�"s�%ʙ&}BL&5d�X§	�2�67�����S����b�d,0��o���K.Q-�:�T�O���o�h���K��r��ݻmg��4�=���e��>���l[��\��0�4]�媫����~7����^r�]w�	���DV�v��p�|����n���k�P8�E,E���G7~�z�J��.���(&+fK�RC�`�?��Q��5�Tf�,nS=�U���l81���9=Y�*�]�愚��1v���oj]]K׭kl�Zq�K����V^�l��ۛ�=�+7>9��o���,N���9�)k~ڨ�k׮���𣪙I�sE�fd��nR���f
]u?��+%��d��ʏs�X�|a�` ,���8!�y;�"qmEW�[�l���i��ᵫ�]?99�pC~ȵBQ�$$��h��f�m�T3�s5�(�5ᇠ������B��D����0���ì�����kǶ�8�Y�]�=	���&Q3����KO?�ݞ����#��=��k��6�x`),_�T����U����}=���3;����c3nFM���	b�F��lP��M�u���yj�s�Z��{��K�ZiÐrV��`G�)�w��֐:LGk�'n��X�� ��xB����Q8����!a]B��JT�s�]�K��驤�������m`�-]dV�{�q���h)��~����}�/HF����xh�>a!���mh+j������|zMHE?�Uq��0�-Vs����h��A�N�b]W|>K�����6Xe��@��8��YE�`�T��)��n�@Lĸ�Q�-T��I�Q�F�fbX�`�S�M2F�6s��)I]F[ZF@P���F��d�*v��
�5�c�3��� K��B�S���$tc�p�53�������+1d]Xp�-n���@7�^[�|������T|��{�I�������5���3�]�y��� -TۏT�֊a�C�}0I��U�H#��"�e��z�DjhRQsVJM^��M��v��8�;�$H��t�L\K�,.�T��G"�5��h�iR�uC'?�$�E�T"?QO���w&�k�$��Ȱ�r��,���k9ð� ��^�����}��=cu�� 8���g���b�D��-Ն�{�j5�
b�j����$.4�'i��P(Ki�a�!؝w���{^C�3XqA�U�v�e!�5w���y�r�*f	�RC����@�O�j�_���ý^�B2�C��	7t���J�+��N���F+�R�[�J�g`<�U�����~��g��͛������Ջ��ȶczI=�"%J	a`���;	��b4LT��;6�}lu�f�g��Qd��&!D�'��<�g��탯OM��D���}%�v�L,�n��م}��HԀ�QVTI���,�@X=����}�;��j�1�B�l�řC��������0��%>���4��%�w� �^}���^x��,�������/���].,:�΃�6������奺^��=��(���~�ُ>��qǜx�	kӨ�������'�믹�{���k����r��}������_���r^D�����d�p�Єk{��3n1�c,:�|����ç�R�NK[1i�/(�(F���y0�";�S��Q�+�ub_�Rj"T������~�?�~���JY�d׋M3����c���Vd���C=��Sϟw�
���?�S�7�m��V&^��\L����|$���:�U�Z��}�xIj�-��O\�c����?^x��^yn#�z$��K;��]�z��Zoy�2L)'5~���p��Ծ(�&(����̈[n��O���[�
":`&�m�SPR�&a
����?�я�tn6�����F�$��Đ�phM�t9P~)PU+{��U�����0����S�.��Hp;��Wn7Q��+;��4#��n�#I�x���T�ґɝ(J��7LDQ�'����&�e�A���^{��׭{��� -�E0�2��'�j��S+,�ǟxy͚5�ea)HȜEW6���~�����'xLà��0�m�'������˷��_��_��m	z�ˎYf�aP�~(��ul�_�|L�0a��w�w�~�۠<B�y'�����D�S��j�曦�[xڮiSs�>�{���^qhܧ�5_�lݺL�h�^`/Z���>�9�l�B���_xm#rn����Rv�|��'�,^�j����bqx�����r	�!��ËF�.]���m�v��166�0Ô`���a>n���O��`��t��_���=p�����*�ާ|w���2�:77���/�;@�+�q�5�/r��N%�@�khD�@x��������wxk�c��
��ʕ+�O�?��;7{�W�^���=��c�-Y��P�0�s�� �d[�ly������|����.��w���WNX�r``  ?���}���q����=�^x�C_���j�8i2х��`���H�bׇ�����ISX-���Aju�X�V�!�e��%~g�l}�jg4��Hx�u��9��i�������/Y<z�g�1�'���zF��N6���B���P0KӳE���EC۷o/�J`�r�	�{DO�s�b'*����%N��ÈS檂O�<X��ަM��ߠ���f�#� G�U2��Q�����Hh3ccX�SUL����(�cw�J�OF;�B'�V�4g *���k���=(�@̴J��z�1�+�p�k��"#v�'���r5Y.U����A�3�����E�� �_�J�|�������i�;oݺu���0ΡB����y"��?|�O/�B�:I�l�$��H�/��Q���'�"df1.%E��*�U>�V3�h��o7;��p_�f	~�2W
9!�jTT��٫R1�"��k��Aa��&h/'v�$r��<�{__�<t��w�wL��t&���6^$&LH^ .x�#s��@j���"�%`Qܙ���v{�I�Vv�[�-�A��a���Bj���(���:�OR`B���	R�l�&�c��5n�-Ukp��^{�Z0��pk|���<�/�Ջ�9F���k�/�
�t�'؍�E�~��sE������'�PȄ!��5�N��r0Z>���[r5�Dy|�K{�����HZp �OnUU�c�#P�qB����A��u����7W�	�܆�|�\�=l�����|�#�}��2��� "똮�����z��~��z�P'�B\�^z�<
�a?��.�R��v����7l���#�ƶy!��w_��W��;*�;����/FD���S:�X�wx�ðo��r(����M�Y�a�;����>��@j&E;Z�9�_28�*��cs#<�l�4�ilVrE"p��C�d���9��|�,��>Ut�`�_��g�}v�9�P�L�!��,����p�7}�&��BL ��E ^�˭�����u�w��ե\��/�_�z_+E�����bj�!HA)��W6n���ρ��c��q�VRAx�|�K��o������ם�a��:�*,
WRq�=?�7�q�3<o|f���Nz�g���ڶ��rf���RķxǕW^��i(�WGlnI����\��J&w�y�W]'B}�R=��� yMC��h��.uh�Ј�����Ңga��w�����&����A�v����
�+��Y�Æ� FR�T=���.���҆�/cWOe��)�ɲj�qp/�pѯ~��.G34�1���o��'�����y#*�D��[�˷��ݿ�����;�KB�~��ꖆ��#Yӟ��s�]w�l���������z������o��7��WnYu��>�G8#�t׿�;3_������ϸc���g������?t�{N����o|��VW,��]C������=?��5]t��۰|��#��YU��*���/��Na*���H�U	5���t��D�����AC��*������{px�V����]?T-P�Ϲ��\��� u��ʉN������n�R[�
��?���g����5[��G�>1=6>1;W
��,�-��!�NNb��v�������}I�����B��Yq�R�;���2�f�`3�ι���3����L�̈U�q$� ƺl���5�1�m!p��B�
�t�^�]4tҩ���X�,$�ހSj�NWW-�b���IK�6��B%��^�*�<6>{h���;������*��4-�=<�
����2�i�if���s�R�z�~;��ȧ��m���53Z�\�
�h��g��.���S���!,��V�L��IY-�D�F��2� |��ˮP�5t�R�I��'єJ�^�א�8M�8�;)j���,��ڄb�lI�p�`�4
٠L�4Yp��;:4���-����gAB%�����#�8Y]��ֽ{����� _�"3���'��Y�s�*�"&�m?M��^B��n����'��f��l�֠8�[��a�)�,XX��U-�W	Gvogj!�=�.bP���2W\��󅥹y��"z�DW������r�ED>i N���fVK�
\lAUIl������)�������G�}ꖷ�"Ӌg�6M�^��"�E]��]I��m*D fQ�MQ�uw��,2������B(�y�^�S_	j	�Te[���
Ey�dqn�\-W���"#LM�.����5��f\����"�$P�a����bU�q���lcʶ�AɅչK���m�U���DU������S�ծJ���݋���aȤ�e�����26�b ˺�苋AW2��^L�%%Q�8�R�DD*��z"�N̍������Դ��;4�q�}� 1GϭKX��H�`_���8��Lz��*�
I(�Hq)�{)"JLI�)v�Ы�AF%!!�r��:�h�(�-Q�<1�fD�f�m�Y�~�;�д|&�J6<�e�` ��O)sx�D�^%�w*o�d��-b��M[P��poщ+��L��|ġ1��CE�L6#�I�l�A�%jiTkTY��/�ʕR�������8����q�>�
Ìe��-W���M�5|_�����ـ�7��a�� �=�or��p�Ta�.$>F	�+�^�жyk�A�v���m����y���1b<c�g���>���E����Q������(DW'�?x�Pa�D��&�Eh�c��ݳ �c�)�2d�������O�p}�Vx��ʟ���W_,xj��Z�y�y��jy��P[B,ſ��"�	�K?=b�.j=�qa���BN����8Ң#ێ_���$ȴ�/($ǐH썷�]\���y��o���l�-y�Yv󷑮�����i3���c~ ��q��mrՊ4H��8`�8�;��Ho���n�i"�����m7�O��C/ar�X3�j␜zI��^�O�)#DY�à�-��#|H�{��=�R�q��y-�7�x��8=��眚j��h��}�s����N;���߷o_o^�:��Qi�!�'�����O����������~�\����7���L+��҄	c]χm��9D��s��#�Ț�	C�h0�h���B��q<��sE���7�G�h�a�w�]n�aZ�o���5�e��a��`�ӟv����~��W]J�s:H.0A�J��/����<����<���m[2��D�\U1���o��o�n��ؓO�J�EC$�>�1�� ��r��k����G�8��ӥ���ꭷ�|�ͧ�}��?��'>�!�����y�0��|�; Q`��-[��o|�/�Ͷm��:�WWup�){����(�����O?��aÅA��tS5=�RG�o��b��#�wF|��@�8�e���ț�k�]Pu������� �V1K ��ر�駟��k�6m����I�=�?���?�����sβţ###pMC}�����MOOoݿ��W^ٵ{\?U1��G1*l�6��S?33S/M���?Z���uttT����U�`��*�_��#�<23��hjg8ꬴ(A��v����W��q�P�.������4+W�tL~��}�{���-�MN<��30]�00�\�O>���q�*��������/�'�8�#�%�"���1EjD���AB;�s���[M`�#+�����Ⓤ��fs�t�^�7n�����Q�RW�O�72��FrLde�;fe쟬�O"��hU֗���N;����W�c��� m���C�v�ٳ'!����<�Ll�%K����z��e�x�U�V��v�ޝ��ID��O)�B��H��\�YJ9S,��l�c�$U����&@{H1�$��L��,�9����cԠ�_�hqBw��:�_�N<��c��0ڃ/��*ϗaT~�����_z�6�-`OZ�h��}�S3��ܢ��ƹ]�"�h>�G�\Fd����f�Y�r�&�$ށa�A�>66f���͛�����$V�����\F�{n��\����^s5��x��ñmF���\j����i��.�V�<�ǒ���ꔽR��M)4C��k	b�;���l1h�*X�%�P�dO+�F(���$Zi�fΊ�`rĐF�u�4���Φ#�4�F�[��_\Xp�Pd�L�^۸q#|k�`Cb��;\+%��~;[�#�i;�}T���.�>���w�1,pL��&<�Qo��bm&�p3�}���F��p�r3��O��p�W���<����ۋ�SD (�=�T��mq&;�\~v��lL�����O,8`�SGPʤ|�V���v���I'�\�+3���� ]�>77gY]���g����i��(�@D�}b�6@q�䱔([�m?�S���\���*~����h���5�#0�+㡚D�-R�A���0 6�fO ��	��3e/[V�ĩ6��K]���,���Q��Km���r1�/M3���{�j�X�L�N����'O[҉�ٹEi���T���J���ґMYo����#�oW[���q���m��O��?!�7Nd_P���P?2V��y�&�@k���7?�Mlyc����+��r���}�>�f[j�`M�r+~)9L0�X,X�v|��Ŀ�|��}-��d� ?Q�Xi�ܟ���=������<��S�065�s�&2����l��7������/�������us�E��"��z�t�ʸ1�P�T��S�����gb'%�G�	�L�cpU�C ۨ/�a�t���L8%J��j���e�2���Gj�:v��e�*&��1��)K!GY:���V�ρ��;�cIGl
5l�	`���{�����3��_��ꏁݠ��
����8�������<�ӣ�����؏-;��ut�娛���z�8$T3�kYC���?�����'�g���/�y���"�):0H�вE��o������������_x���G�:�[��<���~���j�|��?}��S�\}��~qYR͞^�=笻��OW�!��,B�aZ&r@�e��a��$���Hy�&Aֱ�39]�9݁��s����S֜2w�q��.)�[3��򂣚Յg���O.��$4O+��Jz��݆�����s�R���q��玎���w��hb3���>��۲s�Lq�=U�����;�1g(�#v���ƭ�Z5Ԇ��<��޾��ﲢd����^�<>>~p����� OP�#��O��C�-�Ƒ���)�Iaʌ��'�
:H��EK���k/����u����Y���,��3�ϖ���M+�k3�jxe�23�_�8�K�V�.�j՜�����nٳ;ok�Ff�i�&�ɹ\��eXP%�#��`��ĚhA7�Pp�wD֡�T��o�&6�{��Y�c�O�������Z�C��/,���	4�b�Y�,˰�zO�แ���ېb���������/c�+Ӄ���p�X���3�Z�x͙g������=�����X����E0�
��F�\���OC�j���`=��r$G7nټ�2h(1��'�҆ �I�,U,�XLkg����&I
��(f����zV�R�Vu��$����[��9�Z�+6\U�M��"�K�dW��!V3z$r`���-[���?����g�UİW��.��PW�1_��J��hj#{�GU�Ky��[^(�e�rB�A��>���-�$�O<�M2�9�6W���˸X�k�S�,�?Vj1�=�aC D��I����7�O[x�P�zR=t��C�2��Jv¨��M�=3�UAeiĒ���PO��z"t�`c��	DQ.�BЬ$���3.�밗��v�K�̤�f�hK�Ioy���6y�h���F]d�>!J�N@�*�ST�R�Ja�F�PI#id�i��T&j�-
���]�?�x	X�ഫ�+	�.��V�3��E�$�&�y~�65t+����Ga��X�ٗ��±S,	qS��Y��WB*[��	��΢ݎ�|2��9��tJ�#@�:��P�� z���"&�"�`	]�:�eɴ�TAb+�';�s�5{�8��[�lt�%<khn�{�+w�ڵ�G=��/���i,�%
���ᕋ�T�=�H⁌Ō�����ЬՅ�����+��BnhՊE�.y��;�������t�� ��o��O?0Y���طw��f_�95�G���)y	v�a�	zt�� �"�M b�F�]\-?g��l!$�Ζus7v��V��ӓ����sᴇ04$�L��N����P9�7�L�@D`I	�@79R,{^h�7VP�Ć�J
��aŇ�"h���W���N'�s����d	���4�T��\��VO"&��Ӡ6a�ն�*�����
ǵ�V�;K\U�j��;�v���`\^NY��]/n��tt��\�z�A�4X�$�[˘@!�1*2c�h��*��6��R�
X�B���h8,��x
�?	����`�`��jĨ��;��6��P'DaC5(��ς�7R+k�W��)�T�w�½K_�z_�-/�U��K/�v�̷��n�Ȁ�B��/���@6�{��7e�=)�ӌ�J�H��OO�_43��.��|>h�B2!�`���]ʹlY�)�)���oÃ��At��ǰ�Dr�����a'��ɸ:��Ÿpr�{�Zi��R�����rA���u��������|��C]C�Isq�T*�ma��cW=��&^&�=��s_�e�%�#72��fK�b$��Wܵk#1Jq��"_��7�x�hÆa�y���2AU��?}�+_��~R@S�#�2�<��{?�'ǞzΕW~,N����Q�x�b	l���@��'��HN�>S0��Z��-N#��K܈�����W�Z��@����/��2�_,_�b���b�׿�5<�������9x�3���8p`���o��#�ُ>�}�x��<�FI����_���k�r�?�6��ć����g?-1.h��}`1`�̄0w��l�IX���w�nG�����y..�-�'֐ႆ^ �ېh�U�~�&�,.�eQ6�����8��xꩧ`�N=�T�@܈Zy�ouu=����m�a�=]�j��'������G>}�駿��/|��\�bEoO��1|�K_�������N���T��_~��W_�R �$�R�B�IG����[#<�]*���oܸm۶�+�Y�~��;v�x�Z222ҭ��х!b�[�r��� ����j)k�z���;�l��s���};w��.�����""�4�B
p��%�z{{�M�r�X�lY�ma�{�~88�	�3�¬�/���v�Zx|��knٲ���Ƽn�:�����?E4y�ǝv3ߴp(tJ̡�4�?��Co�\����BL;Lժ2����w��R|�F�XO� ����<[�$
�~k[�+'��W��lxͩ)��"}��}kj���.��r�0��E�ɐ��P1��7���G�����w�7Q��r5bo�@&��j���4�$�3���G_~���.�nh&�E�P����%}��:Xw�%s4*��5�o�?#Z���[D{��̙�&%dȲ��5!���Y�&�}�#���V��wZ�����a�B�c���RIj��2Ĥ}4R6�����F���V�Y��fM�8�vo����ʘ|�A�8x/,>|�����9�o*,2�C�s:�m;]�f�j��O�[���+�:�Ң�b�Lh�xq�{H`�%T���)ؾ}����'`�ds0�O;�|]QY���r$Tj���r�S3����<����>�y�G���+b�����NY��"����V�iQ��7B,L�1�Ũ�9�ʇ�SN����OڛE�T�/��Y�l	���{�N�b�/'�x"��;7˄�	����R��FU�R��{�!9�K�:^M��w��.o� a�Ϙ!g��xҘ����0QE�	pDz44�V!��D�6�+���W�����DM��%���)�%��^���h�r�kJ-'�y����#_�i�~^>\�o[\�9L�TI�?�
�����|���֮.i'��6 بRj�T����zI�)�0��`�Z���f����a�P?6(��x���-�X���ᦲ�L0-��r�!�I����\�����q�����������20���9�J��>��҉��z5Z�d	V�R�� [\Bځ�Ғ�.���k׶��/��	��O~],ʫ8�HRCG8�}��O9AN�cTC�'q�7\����'�y�qj�a=��/�>�ll�\��5�|2��SQ���A��:���_��|"�8L���*Ha7�Ȝ�g7O����G�3�G�*�[��lm0�CܢN�Z����a�%E�A�Ea�u�D,Y�԰@�x;�*�<�1����?1-��Z��H��t8����\��*����'>���2"-J��NRKSFj�{l�leF�Y��y�
�p�Dϰa?�%kK��\��泰l�&�X��_��'�0o�:���^|&�3/�'i&�,I6�^b*5D@	�:��(:��H�eY���ᑨ�G�HY�P\a������Hrͯ�ӢT鑵�NWP�?���Т��7���:h����bvN�+Uҽ�A���Ŷ������OrNF���k�2�w`,,Uf�v�t�l��_�&�Zj�%��-�gm��FCS%F
��C��T�4R1F"��$Y�'j,)��h)P�����&�-U@��s�L���g+E1����h��%�k���=�ő��F��t���9h{|�]��F���3h�f��"5#�^�Q���p��t�sƺ0nd,k�po�W'�*���`_����2�^xaӫ/��.����|~�ɂ��q������8�^;?X��WK^m�i��z!�2��F:�3���?��L�BJ��[�(�ze�{��Ʋja0�P~u����8�l�S��]Nyz~j�Q)=�Iy�	W,�o�م���
����#�P,crrr~��i��$����^vF�o����3���H;��dp���3ǩ/��Xa��������l&s��!�����:7���uvif6�rh��� Z��d�dQ�BJr,!��ly���n3���?��6X��>_���-���)�08Q���jK���q�6�)��dT�����z��;��/WY�'��'���dB�rp���m���.��g4������FQX�%�/���p��=�B,^�Q�~ ����M�p�#���Y��F<</��R�(X*GXB��]*K3��.����t_.g��u;�H�,�K�_�,�%#CX-9_�$bέ��шZ��`LBAlR��<��i"L5���b��b�Ѣ���Bf"ʷ�m{�Mn,���� ܏tI�Y-i3����T�|kx3��E����䱤ܗ��+�ŝ�-���p��;\鄗�E�6-n�Qj���@)��؞���HI-���N�细��(츦����-��;d`�[ Bd���92���,[�C��$�LWa�3� �[28�2,>�<«� ��
�أP��%&\Ӂ�Zܜ<be��aJɜHJbC�`���Z�2E__��d���It�	Ճ��蝈���M�o�ޥ˗a}�"L)�X����d���m���ԕ-��ꥅ0B�F��՝o�5��48Ru��vIn��_4Կltdz�P�������P�v2�e˖�^x����r��T��h8��$.<Q&��H5��ۤ= �;J����Q`dɐ�bך�G�v���a{�V�k��B��$L�&]����a�(�FA*��O�T6�CM��E�1ѝ �\G~(2��IH"\�%tɒ��QT1(�+
�-�}I&&Ub��4`�)����~0T�6is�rG�_;��FIn� Sg���͌ف�����x��������9��6�&[��h�[�:�p����@�jpK����&�@C��o�Z��d��;����d\"	S�@�$��Zp����j@��Ӷt4zbak��U@�
/�[�$��������1-�R O:���[IH;K�M�x��{��=𵚯�T�6nܸfͪ\.�O)^_�����L����W�^������a���fBU�
St��fD��{����?����j���.��R��9F�K��`�۠h�25A��ݺm�1�;������86rl�Ԫ	>�Ex�;�[��m"<>�A-�w|Q��,(���K/�*iE�Q/�X�뮻���MH�*�tI��G>���o�bE8w7�x�M7� |���X�k�`
�z�y���A/8��\ޫ{/���ʕ'l��
�S�u�bz��)��r��%��`% �!�����_z���N{��'%�g
2X�'�čdjf���F^+.~�ZŊ��������Z��cǎ׶�D�O{�O�1޴i��͛Cbw�bj����0Igff��ك�U�v�܉-lX���n�[ضm����`/��u��.=W�ƗcM����Q��~��G[P {�*s#� 06b�kT[����G$�1��Xvp)�d0�F	
8�~y3JT�/�@̨��r��f�k�=
��I�ׁ|�'����,vm����;�oO���!����p�w�}�yH2�}Goo�L���o}�e�O:���<x ���9s�m��_M���t4���o_ҏhr3,,,�����[��(G)M�BR1f��v����˖�?���=�㮺��V��	���+�C�G)m6� J�ҕY�v�kV�`�လu�	�����د#�c�D�{f�𭌉e��W�8��S�w��gO�l`|�7�zz����[:���B�,c�2����]�`�OMMQ	36|�`���رV���D�T��\�i(���i˲`9�9
�+���I���>��S���-��ك�`��2�3==}��u0*���>>���W^�Z����vM<����J
��Ip��+Wv���Lpe0x[_�O*�"�S�!N-U���g9��f�\��@�L�K e��}��CH��pTa��L�9�w#Xk�=�����co^Ԉ`MA�`4:F>�cs|7[+��R��^jp7h j@2<A9�@�j8e�b��#y�I)y_�c��3���[^
�͝���1�TV�i$8����e���Y�ȿ�ӥ�X=�����q]�&��CѪ�j��4�p5M��_��- Fs#���R͟���cJ��.�{g�K&��8h򽢟/�8
i������/���>���^7C�����;�~k����}�������_��d���(��jDSL�5P{�RC�ޔ��L�1! �n�ҥ�S�9�8�p6�|�A�S�s��}=x�@G�w�y�V����0`�6�pӯ~��Ri?ZV[�7��ӥ<Cr�&H	O ���D Ww��V�X�sz������^s^������̦9�촐�hc���9�#�>jYl�����w|q��O��q_���*fG�O�BU�a,���%�c�F�;�d~�]C3��B:�
Ơ#�I�0�2�|����n���a��P�ZA�_/�uM��'P 8mji�D�@�0$9q�~LLȐ���{�넨,Z�UGjKjQ6��,@8���c�,Yh����,�޾N����uz1!p]��Dn϶-ZXe|~d�ZD:�����J�@�� �%p~USA�9�[�9A���-�QL�63���p	�;�,�Dƨ
y�DG���
l"{�������TG�'�cs]�ȡ.YFy�ڕ
9�����An)�0�|�<�b4�[����o��+���1I�����?��䒏^Z�E#�m3uÆ'%�$�����GW]�au��T�˒$����Q���M+N2���]�\�D���W��p7��L,�����S�iP;ԣ�`�ţ����-:�%�bEbhM5���o�@��G:�rt�ig�%QL�y��n�,8y�F����mu��u�ԯp`�5�Ԓu��ӟz꩚ DH�F�3~��ͮ f�����_�-3+tQ�׺LĘ��o!r���IW-̍�\�?�PxDv�W}�����q��w_{���꛾���b.JOK�)p������0X�4V�:�
�"T(�<��{����G�~�L�T�����~3��	eGE���{�霠�K�UB�g!�:Wra=,�5��)\�X&qa�	�`z|�,�"�LJ���#�c��[�O�� #��f4�\��� �ڐ@V*I5��'US���%�z`�-���*�l��X\0u��oqD|Jq�04�7H1�q��c�B# ;L��`Hu����(����L׭΃����<��G��v��i���(Y��;0���W����m6usS��ݻ�������� ��h��O���#oI��v�Z�pw=��V�)��BBtce��20��'JP�W|�L�.2�h&�#/Z�lx��7�gϞ�bfr����s���_����)k�QY��;_���z�1W_}��x<�y71s}�^y��_8�`	�ۻ��0q�k��݆�.Z������/9y�P�$�ʥ�\r�g�1r��9�ߋ�-��d�x�v��������3~]�����\)������S����ɚ�l���1���$hĲ��0�Pp1��`2� 1%kYD��I���-�#]��ߨclh�şZ�xqv���n�x��^y�Q0+����r��=g|�3�� ����`)���o?#c�>y�9���hLE��_ڸq�zp/���^�Œ��~�V
�bq˫/�g�Mz2��6�W�v�P1T��TU]rE(�\[���Տ�D��^<�y#U\����I��,l���^w. .6C?�Y�fͲd=xS���K����0;v�Y�V�9����ˋ�63��	x�s�;����`~B�b�ښǆ@��l����0Q�4����$��Z�G���a����%4Y�_�UB����Ha�d����Z�<d*5�dD��Qb[&U`�(
��H���y��h*�8�E��H	��]TnEy1|�L�#>/8Ē6��P�L�����(S��B�$5��Zƃ?�[Pb�o<��੥���,��pc͐bËEգ8��s�N�����Њ���L-��PM6�7�19]���g�����i� q��\� &��/X�F��� h|�\E�E�ęP]���T�չ�ٰ8P�*nc��Ӗé�nT'kz_�k��N�g<�w�S��؄9ͩr�`h�Fs��Y�fI?4L�Q��
t�f�1�p����e2u�N��î|�ٗ��\>s`����ge�(�EN7
q(׫A��`[_OA��³�׌���*��HS9�gF��=�d��j���ת����~U5���J�L���R��A9����0�,[P�H�֝V&y>�ĝl 3�H�ё!c1X(�_E�C��ꆌiDTAQZ���) �G��؇0�j{�IE	�*(�����QL��>LZ�ʱ�ت�����$K�0��IGND��ɞ�x���ЅPul���I|y�dtqtčͮd�.a�N
�s��J��hDBI����VsA�:.9��.Q "�#�����4������B�vL���n�J[��m
���R�DJb"� V:���%���p�b����+5�`�P�b�C�N�&6�HRG��0�h*�f>Z�0���+m9��)MI��!Ņm�2��):b1!�jHS���,'��ƞ�fJ�e�vF���L�׻��j%j1��Ѧ(��͛����W�6t�G��L)����=���K�,��Ă��]7ֱ)!���֮]{�u�����'�pL��:&^E����G��+$��d2w�����^�@;K-���qJ���x�� �����,1T�j�����+�Vr�]C��5RZ �D�zE�!;5mQ!��A�L��uE��8^�l��?�o߾|��(�;H�^��F�g��ݧ�w!�&�����y�4��y��ob�T��s#Y�
)��1B�n2�f?޻wۦM�N;�x���Pb"�[�2��K%��_VVG3��?�V
Y��ɥ�^z�]��\� ��I�^�~	JSHM�G.2�*�����Rj��P�ȱv�G�8��H�v��EA��I�b���.l���x�1ҟ &�P��U,�N))�)m�ϫ�r�G�R'��4A�H�GI�̓���3�/|g)I)?�p���\2;�#�|�f{1	F����j�^ǂp'�bA��<$l�p�3�B��W�6�^wW��$[�RE^�����A������ᘪ:��đx�W�z:<���G}���_�.= ��9���O� 9J��4����h{6��q_yz�J� 	��x~綳�:��SO	\��۷�hJ�P���bC������KR266��o��+�x��@I���+����X�K0��OZ�٭�Ix���nxRd�"�csT}vv�������"s�ƪ��n��V��u��HnK�f7�>�m�B����|���~�¾C3�2�#i2|��A���ƫ��G>��GF�ݝ�����\�8��p+p��}}v� 2���lL�/�INh0���bybMMM�q��S(�}�U�	�W�謁^QĠw*j��@?Lc��J�1?4��D��R�F��3L�[9�V,?��U�D.�j�|�޽{�8p`׮]��6�~�i�j���^�t)���g�O�m�w���G�s,x�*bkI�:(�ZZr3cЖ�ͪ�����_&�&R�a<ئVk����ivd5y;P����r�X��:�{���FHm�\������R�6R����W�b��3E��px���	TO]6F(Rl��B���7W'�iR�8�G`�	�m�r__��=χU�W�Ēb�͖���QUp�%��í{,,��.�Z�ی*��Џ�5]\WT��c��i.Z�H� sw��@Y�ᔨMiB�Ɣ<#��2�d�F3�7e)�,LЕ###�����۶�	��q��I��b�g��'�Q�"���X1��:Y�O\�3�(п0?T�(�0����5���Y�)�	G��ϵ�����o�� �1P聻�VK��E�#EUh���?h��V��@M���{�H���E���E�dj^���	�$&L;��0�� ^*�,��>11y�R��bV��!�2��/���� ҝ�NDd�l6<���mX!A4.W��-&Ӣ:nL�ؚL^*�&5�ĭ~QA�I����o�^R�{�S��s�Z��n�O�W`�m�uF�;K��
U}"H#.&��C�j4hu]�LMvZ��hJ��S�L#��)�LQ(Sڊ���1Aݫb9��|�NU�6���!L��a$����*qb�b�fԘ��F�	��k���d�:��ߏ׻�ׂ���Q=�����=Xԋ/���_<	��i�O��q���j���)�>�dca����T3����kZ���T�]-]օ������/��g�z���݆lK��J�V�N�
lP�oT�lN� *�F`����@R���A�v�Ϙ�i�����J�ʳ�)�o\!��?��ܑ%:dgT��Y	ц��Q�-�S�_Q�?��O��	8��i�1e-&�+��'�
��c�?�$���jY���C�� �u�Гa�Ȣ�sI��b�Ob�2!0��H���v��QBD-2�3�?����=��ÿ<oݪ�BY���N�7�3�?Z��~�O/肉��@KIT�A� 0�#��Ǭ^���/�l^�h�`���]n��e|�vp|^��e�	��@���L9��r����	���V�IT���%��ٛe_+��X��U:IO�W5�l�Q����i��'Pcϋ�6�NU������T5�d.�:<w�VU�CD�Sj���a�RpB��e��a":$<���4�����ð�]��*#df�{wÖ�{�^:�=���(�rxt�d�h�Ȫ��z� ����O]��	=�=[�>9���DU�4�cY9���f)���X�?�#C�ٺ_�P�rZ��q��"@ٺϔ��D	�-��3����B6m�c����V�Z���6�g����d���0��ǌ��=]EF�Z��xJ�J�s�]��O{���O,,�u��?��ǃ����j�q��e��^9���A0bUrt��P����۵{��yjBl����X(��0��^�:��x����3000�x1�į!�x06Xz��.vzb�t�5993�ۋ�.6�Qݑ$�����&��
vd����D�s���V�x���&I�����-�TFz�BT+�˗�v���yˮ����?���E2l8���.Y�j�k�o��mXY�q���[�ik�v�3��=V�]j���"Ñ�r��*z�]0͂n�z��{#@�Ђ��`!�弯h�zy^�$�S��ii`��67���6�d�[������f_�L��������?��?���>���]��]����UB��F����� ��.��OoSΜ^r�CIHHB �
,@T�.��u�r��˂���/��������E��Ы$��~r����y��|�}�g�L�����r}c<̙��S�����r��6o�yY�l��l:�`�[��l�!�T �ȸF`��0c�@	A,
.��#k& ;�Z�"�+b5m��G�F�����N�@������F�d��	g�85�KӁa�d�B�h\'a9B��%�1C���@�f	�T���',y���:�.��� Do�j���P��Zm��X!��dYOg
���[��Jf�i�쎹s˅��͛����o���
���T�444e�wq执455Mf'���ǆƷ��O7�O8ᄀt����ɩ)TR�0�L�@��(*N%є�1��B�����0k;O����ϑ~����~r�uՆ6JO�J!?�G����Ŋ��L(;%۫�(��%�i��X�/�t\SkJ���r~�ξŋ4��F������'�=�L0�$`��sC���oO��X�c���`��},��ܲmw9(�s��n�vGF��Q"�U�V�m�1��0&�G���2e������9����YⰍ�tjс��@}���#����|��p�hF7q�0��[�����BA�B�0@F����dQ	�Ih��+��K��9ꘊhw���"IA�K�)�&��J	�!4dwiJnYD�S�pѱRQ����lF��쪰}��|W��#=�����d�-�"�"p��z��W���Z=g%֠��1`�-�;�p�x]R=����3��`�K"�Q^�K�0�0��b&5?��JqlR3��*�nd`��gʀ��E�M	��|���Vp�]U�����r�|��pgnٖ��f�u0Ì$}1�s�@]�!�Pa$©U� ��w��`ao-G��|-$C�E�0U�֭�=��o����KԾñ1ః�_��F:�w�w��P"X*��*	kآh�g|�c�������|�K_�_�T���[�TL;�Σ���pKu3M�A9
���0OL���� 
w���T�W���ZoX\kab��u��+�9�m��*upB���=Q\�%"�>U�JȆ������c;gΜ����@d
Ղ���0U{�n$ݣ�
���`�*X"ί��/�|�Q\�����9����������o��������W�.�<ɣ�����'>�	��G?�Q~��g�J�w�_���Y#�[�Y��{�);Y�ꪫ�����ݻ���#Pi2���s>dY��U	�2���9S܃m|�Pd�\"�YEǌ�j6���H��xOG��9�![�<�HU�l�L!�����D�-�9dI#Ooɍ��xD��Zd��5���Ə�����3�Y�4Qʱ�͠��$D�]�j���M��������7�����D��9S�gc�\�S�u h*߹�:e`�[ዙ��C?��I𹮨<ҌvL���7�aoL�^�gh�]Q�����i94�M��-Z�z��;���͛��U�D�"(�oxy�^|���H3�E����ջx�i���������˹\n�3�� �_��XMA`Ǧ�<��a�zgg[[K��ٛ����];��NW�;�f��Ba������6���`�v|�i����z��,Z�255ŷ�Ä��^{1s��V"+rp�S����~x�%���6l?�7k֬|6���+�̜9��˄�/�����W0�g{`G��z��'��,��Ջ�s���	���""dDj*�����q��z[��G�!��)p'Q&��0E2wnr``@r�T,9xr����u=�`
E�'H���1�a�x�<u�^�@Pa��	�d208�?�8�\1|���H(�,(s���ͪU/خKZ�OI��dU^ߥ��Z5 ���7 �q�AI�.���s^,�1bզ��rkP�u�J���?g���YÑ�z	5`kV�fO��I��NY-JkkFLa�_�J���aw���P��=�5�;�e�>��}����Z��m�8R�������?���SN�흅���s�����,8��S.\�/��۽}l���V���D�y�'�����/�.q׽��V�@�'�Z#v_�y�c�� n��ü:�Y�"��G�Z�����(�
���61h"py�����in?�Y���T�J�D�������
oi�Z[[a@��b��P�*e"�q�����3m�t_v}�4��P�_�2��-����a|�)�1��س�	|
����#O�c��C�|�Cɀq(+(R'$�@�䥯�HBww�S�Ǡy�R1Mq�}������,�e;�,���/�K��#.�H7�.�KA�ʂ�:����f�\�_Aܤ�}QĒ`E������"�l32��,B�S�����q!%}���}V��:�%�u׫��%��i.���ij�J��N���:���k~]0$�˃��BJ�(�t�y�}Z�/�	�FBVd.�B����|���������1)��0�����x�3ojz@4��hT+6z_pg��튈liER�!e.�ä"{˽��}-QR��n;�#�1��U���U�����^|���������/�+���7@~��?�&
���
:�2�]�"����0�?�ُ�~�w�퟿q�_�{���&lh�
#)�sCF��+��x�e�>Ѻ���L�z^AW�}���BU~�Z!�����;̸V�j���r��Qx���*B����_�oܪ�AX�*]�'h-j���/kr섚�jB�sn��k�Y��������g�}{��Έ*{������E�ױ��/D�C�2��� .�=�U�S`�:Q))!̣�đ�����ͧ��fݺ~}� �"ERt�_�ⷾ�-Q�~���g��`G�*\q�o���������/�X)������������ni�;�l�y���g��C��=4��_=8�n��wsJSV�Y�t4V�
�V���cw!i�ŋ�o�����:,�[���3�����=X�X���5E��.1�;�5	�\�������L�/db�"�%��b��Ǥ�te�m�ԇ"7�B�
xc[�W�#}/J"���$�W�C�����(�4����[�4ALI�4�1����ˣw�˃jDO�8�@�?!aZ���]0g�]���/�Wrsa��I�ٺn��ȆP�� ;D"�9�`�����s1 �n/�#K�U�\G�L������U��P@�7�W&�ܲD���A텁jj�M�EcZ0��zg.]�$c�^~��W�l��k�>�L3,��N�m-m�����A5��B��L6��^r饗vΝd��!Z��$8���o߾�ٻ�n� �(ǳ��Ι1l���	�ᦽ{3�ti|
�'�;������m��6+�!��L0����?>x2C����W8�015w�\��`���{P������:�C���Z��� �_�<*��4p<]P5C�%P���䁽��ͳ��T*َ�����~�pR�\,*Fz��7�4g��D�'��x��姽�sQ3,�����^݃�R�"*�����4s\���I�9&��mVo+�.��l[W[:�8���.&�ޖ2�sO�téJ%Q�-�fRˎ��~���V�0<�����Q���X�XK�,������Qhʀ�ZQ�2����%���l�=t蕽���s��'-^l�Ƥ(5g���I�H-]���dr撓^޶�vQY#��v��X�������b�!��`�'��*6Hwe�Y��vU�����g�B(�
M]a�X$+��M��Y�Vx��
���@��Vԕ*U����9�j��z���UEW���Fp�#N��TA�*7I(��¢m���f����ˠ���]UvqTE�g�R���\NV��|YQ�w�#���e+��c��Ҧ��T
BO��xu���������c?�w���}陳�0za��C{�p�	�-ۋ�1�ޕg�i�7�ǟ���^�z\+�|�ݍ�! 8�����Ж�;;gt�.欘`���^�E[*�!�"�!��X��Er|y^{&Px�w4�n����������^g��\!���c�Vs}]�g�u�{��vz:J�2�����&-Y)���	Fm-��ȳe]�eЛa�T,���({!8�j��*,v�_�ɢIV�4�*ܖj���z`��?0���	+6�G�,?�uuvvJ�>�ӏ>r������ vJs��k��Cԍ�T�##{���:{6�B�J�}�=���;��Q�

-�rJ���rS��	c��&Q���\I*��I�酡r��L�|'�t0*dU	�,�:2m��a���E0�,[�Q^K�h��!�j��P5SDDKE�ơ�<c����;B�G�q���L&-�u��B�L*{CI8nޅ��!�҃C�<
G�u=EX)����<�;Z��r|�z�7Y���3Z�`��b5���7U;a=��?�q��UDkY�mZYr�,F�4L��f�'���5�O+	���VT�zXfn��1C��܈�l�E[K��RQ2M�(F�;��1��0�O"�<�01v=(�A�tG>l����J*��_����[������(���|�� D23]_y��O<��Yk�����"ڸ �/V,�'[d_�����J�6Y������l/0p3F ���?��k?�/��/g߱�X� �"*�Ї���Z��2i@�aω�G���K��BRm�!Ul���Gۂ<���$<��������)��V���S�[q(�4�c#֠oꕾ�ڂ����DAQ5]�E�Z��y�s�=���S_}�Մ��=�q�
f�E|�O�ӟ��g�����J�5E��M����h������1�s��v8k��J�=�̇z�̳�{��%YK&��J,u3�3_���|�;J���n���<���|��_�2�	�	�|�)�����P���Եk�]pރ�{�����d�u�#��L7Sǁ�&L d�ל��V�-��!�?���Z�U	<D�� �)jѯj͡��xeJ}ꏒu|�4Ҩ��{�A�	�����������dCR��Z�����FX�(�̙3���݂c���FF��X�E����>/(j��^��!5"2��g��Ђ�Z��Y�
�,��Hw")�9�#���%)��<Eη�ij���x_����t�� �����.'=˼����3Q�c�����e�X,�y����{���K����K��Q�p٬Y���pcXI8:
Ϩ�6bI���/~�7<r�e�-��pٲ���/o����y@L/�u�+W�l^8�B�@{~��܃�vvf�1Pڭ��{��{8��5���OD�ӳ�`jcЄGg믘
�꫔7dF$�dY��dd�JQ� �Ί�֯�J0J�DnlÆX�/�7n|���׭[��с٭r?����$
����U��-[�����Vs�Fe_��͛W������fv��9�
�����X``��S�"	Ns����!�1_��\�t�~�i-Ӊe��5�4C�|o��&�_�v�0y�b	Z�0���;wbAc{�)����F��|��\�^	��4A�D=�;<*L
�ī!E�k�j�G���MU���,"OoqYR�|Z\���j*������0�8\-�wXU���!>:�ŭ�j���i���0S6�z���O$��⟀��5��������&���T$�<C{�Y�X���	o�B�G���`��Iy�������u�:�[aS<��3g�Z�t),$89|�b�
ǭ���i=�v�Z8�m��Ɨ�����Dcg�	��9�D:�M[��@��.{i�䋣E� �W}����1k5���cJl��}\(`9�6AԞt�JÔ^ͮ���=k2�s�"���;��۶m������J%C�8��W�`��	��=2::�Ȩ����t�U�0��ɤ[�����P����T��ٳgϝ;w׮]q��h�";�����;F~x���y��XB)3���4K��2q;<S���/V�kȄa;�'a�xY�m3j�+��s�S�
""ʒl��)�#h	�w���$*��w=���H�pcX��Ǻ�^�H�B9d��I�f )p̝�1U�#b~�a8���
A"<*���X��ɘ8��Y\�W��,pX�S��L(�e���{>S|O��Hp �[k��\C���.���9�,o6�]l�&�nvY�aP�������ZW^v����Ԛ��ո/�$�u��Գ���n���?�y����-[��w�=�s�P�;�䓳Y�x,6�nM�hS�LFuPD���K/}��ǋ>�m��p�E��{\���UY�	\K��.��k_"rW�E����Q�c���|�~�}�s_���_��;B����.~���
�,���Ὸ�U�������G�]>?�/�������g?��{�{Y�\vi0�F�Q.W���n	YH]�ne�H�Kل������@��Ə�ڏPfq��;K���W,���n�����V��s�ۗ��P��zU��'du��'��C/�XB�W ��hj�ؕU+N���˛6�=��X���G�I���>s�7����ud�$=i��~�J`�`cu�*�G����(&�/*���FO5R�)�sʙ��=��7����弜��ߙ�w����!��Jf�6�D��;����{ywt\y�5���{?F�F������_��׾����S��Ư|�d�]�Y*+�V��dL�\Q���ՒJƭL���j�B}���>��2���,>�wa��L}%�@�K!͋�a]�)��`	�m�Je�;[@qvvtp�TKW���������ԋ�2.��i�� ="���EX�c�m�2�ڛ��4���WS�hNczl�lV�"H~��u|,�45]�6 R�0��Z�G�� ��S�)�N���-k�ut�4���Q�L�P�D \���͔�:7�P�*�PF�M�Ev�G����:#oM'le�+�����$D5�n{�q�ڮ�8V�d�f��Bρ*�\�Q$���w�d���e'��k��LL�M��IK�Ƭ�Lƫ�T��kW��B)ͤ�tKX�$������M'0�I�4���� 8�������do/�mgVY�<������&/粠͝
8�H%�#?
�6��=`�au�J�9N ��\�#�V-҃���� )>���9���hj*�R*ٌ��Ҋ �D���UN"A ��f8��cp�41լglf��a��U��I�Q=���̈́Ԝ��!EN �,k�V�#Ɯv=��L����_�$M+RYi��	X��ظ�����j�s��S�5�~�m1M��)p��ID�.�S����S��^��,]��@gR�T�H����d2�Z�P1=q�+d�&E-��pn2�d	Q؃���a_��b
c�c�OR$/�ύ�(Ural	b!@BP�<�#M*�`2,0$�][��d�B2#��f1o�R94=�X��0s�L��׊�)��0��I^0S(�M�>
���G�T��ּ���&�4�@��=-Ll��噮7�~}9v� T�@av���b��Jso�/�Xzu� �d���������d��H�MD���\�l)j�X*;^��}�hg����¥'��,���HSL%���)i���ZI$��^St!�E� Y�zN��R!Wv=�4m���TS�d�ZUÄ�+��]�3���gsW�w�P�YV2�H�8_4�s��h�y58���)&C*X-Uq�i%L2*�;8
�`x�K���I�:jnOv�����"J����r���
�c ��`a��nJ���������۲t����[q�TJ"�A%]Vu���O���zTC�C�����ɮ��]F� X��|��W6�t�I�=]z:�J	�1������Ύ�ע��$��F�bsj��m�����8�G C�u�{�����q~7��?��O~�^D�I�qC�~����[�v�tI��������^u�8!��n!�!�IS]������ �*:9眿�����|�3�va��3�8q�B\�s�.�馛�y�����1��E?��O��ۏ&z�F�\Xx����z׻,S|DK�;�([�WK\k+`�� ��X��0��U�P���HD��˘�ɺ���6�t��B�f}_`�*�	>�?�KQM)���ҁ�a�8"�����n�,tt4��PJh���_.��2�R�� ��z1,Hr�_�u����_�ַ��ž���ii%���l��M��S���4ρ)Ő�/��Շ>�!��_Cֶ/��{o�T����s���[�)�U�s	o��co	~-�+�ھ}�o4���e\)	���D����?�8�bQ��R����3����U�{�U��6K�'*�~��2�peF��\��%D������GbKB�
-(�J(m*�e��'{�>p���q)rO����Sw��~.����یw����{M<҆�r�8�T�רƃ\�8��Z5���]��#���I�#0#�]�K̶}�@xp�7C�����ucWVTD�ĐU������y��_v�%��X�REn����	��E�^��Cd��	�,�;������Ɨ��u]�b=7�j��Pp T�cQ���7��m@��@Pm�95(���j��o����C����G�a��""���	=����j���[��c�+&�j9ZU�* �t�?a>_�R�T*��,Y���������_��q��9�J͝3��e'��{�ŗ���Bi*���3�І�蝣�P�2j x@�U�3�$��ᘑ��:k�#E�jժJ���c�½]*�#�B�����4��ổ|-�J1��@8>�Hpg볩�HO���DK.�X=CK�艤K��d2��2*Åz{{ad�Y����S�T��^��Zc��'l7߉��1�(	�4���+ജt�i�W�>�w�������O��	�,��S7Tww'�m"�UpX�iӪ��}��W�
f��l�AvdPg��M���7��t`` l����[L�d��;�sN;s�ҥsf��S�m�J��f)`,�J�Aq<x�����B$�B�Qt�M����0|�>���^#�w���S(�/!�<��������'�Ȁ4666w��E��Y�=��p����?�s/\��u�u�]���؋�o��6�Hp�b17cƌW����?�z��mO<^"8]����Y�4��})մ<�(4��F`�J�8��!B�u�
F&�������E��ă/�hw�J��Pr�����#M�Z�����z��_���W_z> x؎����;`�MNN��G�ɖ�C}}��=K�Pt��P*uu���i�Z��\���jb�z���
�y1��Q�i���ӕ3U�&U��y��0S!CRQ�d�J)k��0�F��S4
0ƇZ����|W��k���5o�hq�C��~��|l��=.z��g����{Fa�
!�d��'Ҭi���K�M�.�\��gưB0_Mp�3�8��E�����Ϝ9���y���C��z�!ذ\��Z�E��ϱ�ѨF	o@N�lr�7�Q�5������x≡;�����s%|�6x[[|���(�����"�kҪ	=��"��Q�N��`��6l� ��뫯�{�����%��Da�H����X�bŲe�zft�ןހ�<������@G�T�y���yq�nx��%��훜�5�e2	Ϸ7�Q�9��93�6ڻ{`��J�"k����mܸs�Ο?�ܹ��r
�̎;x�axs�٧�8������W�tR��������1��/���5��(��eZ�J|׻���s{?h+��MJ�ր�%X�1�q/^|߃��z�*��h��+�7�q{��_w��41L7Q�������?��/}���!�{� �yR{����D�搌vŲiϞ=�ª8����+T{݉E�	���7�bpW��TH�A�0�����_�p�B���{Gp�����kݞ��X=��j��G��c�;��p�a�B>*Q��˚)֪�؊��$E��W(/�*�EYo�s+�$��2_�qR�8{>�~��߸��/��r�*���{���=��o<��sO[�J��H�{���� A���
8sH��_��-��t�s��y�{�Gq������o��/�����[q�h�Cb2UT3��a~�	��iP���*g[[W�(��s�[�k�"��j��bD���9�*�90 YC�&z����N�$5�5����P:�-��<B=�\�=���zI�3Q�+�=)�v������b8z�܃�[T;C�ni@��13A��@���2t9CE����D�UF�I7$�67ЖUIP# ����:�z#h�}E �?Y�b4��-4ĞyJU��'2���έr�(�I�FO#�$�ek��+���2��*Q�3v�N�"T+r$Ñ*�1�˾j�/I��8��@W�q�ڀW����G�E�4?"� Y5I�K��,������	�┳y'�+���0���7o����G�ż���>�¾�$A6(�Y�L�2A��~��j@]����|�frd�$�ޮ.���ݒb�kA�4�$e`o�@�1�V��,b����8T�)a'��WKqhvM�r������*�X2)��ĒU��0TCLU�'��[��C�VW�&�Dydm�q�E����^��UBS�)��޿go�0�M���+��9�ɦv��'�	��Е�LV���kݍ�2����{ fj����2z�I#���kj�/�(�Ke)!0�z��߃�Ν&T1_���L^�
g�-�<P��QBh�m�� ��I�l�j� ��B����OH,T�{nQ��%9V�|������,�մ�H��4:2��E;�
Ŋ c��В^����lo"]��t��f��݁�*	AM�^�b,i�b.��v*1.I-��X���E�c$��p���.�b��©�}�n:���y�����S�Z� $��l�zRTX0����T"Tt�)�Q�&�p�m�X���d�40��q*��T]�0���� �U��]`!MLe+�|-b�UX8R)n:t�l�v29V,6�d%�E�C�{�m���"l"7B���!����@_�X��ᓈ�T�R�8���9E�D�<�a��	eT��늡�01��+S.-"��	�S<��Ƅ$���
���bc���yYB-WL�����)��JHVU���p.�B��`D��]�p����� ��)j�)���S(��a��0�@��-*۰YʓS�?�721<v%�ݔ���	����ЌL"e(�ϏYa*��S*�|x`D��X����r��O�ZƀGm�_���w-sNEO� �B��q�b	���eX��a��b)�������tBGg���4L�w����.X0w��Y�����{�0[p�m�����8,�@� b�G�	�{�Ё��Vk����-x�AI�,�P��Mfڛ.9���FFm�#A[����*��$�R�w�������,8�ϥ6
E)QNF�U"�ڲ*���q�x��CWD���ʦ5kNc�pٻ.���*T�-K�ޜr�ک��E�\��SO���������W\q������
��O���o�;���ʕ?D���u`4�)YP�(��-;�~��3�z�_��}��eu����>����߾��o\�hѥ�\D$N�=@sD���}��>�D2�f�?`pe�U�W7nzq������D!����0GD���	�	�CC�p[�^���T�h�IH��R�2*��i�Fk���5c*]ke�56��w8y<�5���6�@"�J2�Gf�G�r�q`z���\�g��_��Ϋ��ՙ�J���+/o�(��������
C�M��V��Q����%�����I'���H�/���֜����?��{~��5ן jx��]{-���O?���SD���$�o��������>����s�<��wV3�/����!�񦽲�כ����_��U}�#����.���k\;���B�]�~�?�z��i��F_荿����t���I����Z%o:�P�D��ϛ8����{��'����/��a����!�XD�w����C^)
⸧���5���Z�O�۷|ZP�3{{��?�� �
�̆����W����������5�)E���8=�E�1�R��/�V�9s��	���0����c���'�<k֬G}4W�� ���g-@�P�vΤR)Nq�k׮���K![����_�������D�������%��f۹sg%��6=T9�@̮����*�C��a�'+���쫚P�ː�(���4�֭[g�;���R˗/�
��}{qК�a�r�,��O�X��q�����r��[0{�슇=?���C�凇a�����T��L.��E~w������d	�ژ�ڵe+6�xlr�x)��T�0��0�jT���q��f/�|bIGNfVo�� >Otwü���?�Kk���z�j?�0İw���æ斱�����xY`'Ȋo����y)��[a���]��DFmf��L���Q�5	�"���Ah�L/�x/�4�a�()�՘�	x��x��M��W�(�L� d��%\&zɒ%�$T>���}��:�_xf�����K�'���{aalz�5kV��������޽�P�~x�nE���`��ϟ��Ӄ]a��^x�!.]�0�րP��s�p�$>�Q-m˛!+���\�^"����y�=ؤ�a��H�Dl���/��b��3��p޼y_�N i�� U:::�����.xG��lo0����5kV�w����>�,/�����O~�x3ˏ?�Ӱ��`�D��y������t,m�o�B��{&.���{�}��}����s�����F�g.�ګ�Or2���ARE<bq}E޿���b�7�z�)H[I��ƍ�>�����
L�B�P<�oxx����
�1���m;A�n޼'������v,���3�u��ׯ��_�r���b�L�M"JaK���Y=V*U("����sǎ��bk.�܎�q�FO�d� �[���O8�/\8����+��� ���ꍋ��t^=�X�-^t�E�	a��|�{�������͇=x��?��S𰧜� ������s}p����[ÁR�Il���<���:����w���/,]��Q�
+�[o���������k�=�� ffd����牁|�g=��XS����4����uH�|#��"8�q�'�I�R5_�G��z�s�~�P{5J�����)�~�u�BG�eE��o�h�8=��l���(�����7��,	�����b�LG�@� 0h�x��!e�\�7%�R����k��|7�<����֜���нT��i��p�7~�c{�m���O7�R�7-���Ԁ|�ZD5-����+���b� �}�<�T�hb5�\�	&�`�<C�e�zu98|!��7E~��i|���o��L"��b�Y��H�t�kԇ���F��M���z�}��O�#�����j�S��y6�$�q���>y�R����˗?5[:[��2`!�c�T��e��2f�U���l"��nDJ`b�Zj��L�̭�OLK=8�0*L��IlW�
2@<�כx�Y����c�.xc<�V{Al��g�B$�1��-�ړ� �x�Z��Q�ʆ��J�+{�&B�L�Jkxt+d&a?� ����8&�ɀN�E>�hIW��BH1Sӛ�)�y��2S��/L准�@��
�	����������TGg�q��w1�y��@\�.��|�%�-���h�
�����`Bm�@#��E,��U��0��+CSۄ1��)��ٞ�f�%�,����a�b��x~K�	F�c�-�
	�#�|;7�������+�WC�^ڡ�b臊�F�F����NM��8B)`
46��
yl�챐]��EM�R�Q	����֥���L����U����4�\��øf,��1b<R�z���q�')!�j���KXuO��d�U�s����4���*jLq�1�9w���R}���
�`J�lo�^A��ˎ�+���C��ǒ��D�wqU�����d2�B�_@��N����T�����\wd�Q*�7o>8k��'*����C�j�tg�feҲ�D�ސ�U�p
8m��G*&K�8Qct�a�q�"��h��υk�}�ɮ����%S:e!�,岹���(�mz5��e��M/������*��ɜVqQ��?��3����~0Ֆ�kʱ��K,���"�E�F�vڍL,k��[[�(��1���ɼW�3F6��R�uż�U��ʴX�"��|l�����[A2(��U�*��\BD�h���X3QR	1�C�ay�K���b�����_���I'J� �Wx/xq�Ml��[�4�������P�7'��{Mɽ�v���:�P�*��m�I�g�����Fh�lϘ�35�9S��n�\6�y��� )�p,�����t���x_���x�!C�n׶����f-���&`�(l6����{���Zgu�0/98��iL����3b󍸂���Y��yO&�j�D�
K1%#a��/�D��Q�ts"c6+� %��L+Se'�s��xd���\�V,�e`�A؊��dāϤ2�=�`�ON�����j��2+���D{7�֮�l
�p``YȆ'��/{���M�	U�BYI3�M��:i8IA*����'�J�-�\�tig&S��颜�����"�N����K0]"P���d4�~����~�+_������TҔH����\��g>�s�e˖F��DZ�2m�����jv��7��͝�s��5C�RǋCC����������g?{�	�᫪(S�(�L�)L͜3�[�����|��y�7� �k���~���n>���<�"1��p��n��F���+DIr��0�b9�u����%�:Nn�X�*��>���=���Q�W�m�����	�4�y}�r�E��,���"&�����z���/�类��w_v�*�"����_^p�E-m-.h��t9��n�x�TMI�W�X���5�]��_�y�&�n���q�U���;�+�x�%�=�1����փy��Yk�v4��ߵl	l.h�b��ܞ7�w��=�Z�����8&dI�m��z�|��(,��&���C�ׅ�7{Sk�����f��u�����O��.���Ax��c�ǝ��GG8b�h����9�݊����+�k�𘓎֮�1�`���F$��N�[v�����~ ���]`���r�)s��EԯlL�*�$��pB��u���B�z���tm.g�2���p���֎�����(�/_^�wb5�K`A��yEx���]a!V�499;�t:5/�x��H��
������p�Op���a0/��|kk��'�<92�o�2����r_�*���&%�k�N�k�b*���n��!����cӦMn)hjJ,���9��J���-U*���@�(߱cǶ}C���'̝���1b1'�1$l(�|�
��a�R��7m��dJ��K�σOJ�!�a �&��X���ބШ�M�("6�FL,���5===7�������yǋ���3�wjj�9%��E�1PM8�K�%�	\�3;Ѓ�B^���t]�-��L(�{�W���aw��oJJ�\s͒�+�+Y��U3�~����w��ϲ��+}���JHQ�l�ÃiR��`=E��A	�c<`�8z6����V��a��!�VQ{ӬY�6l� ���	��_|q��������fw�6N<��spf�P���Ю����(\�v9�$�ˁ�L�..RߦӥRi$��坖�.��⤨m߾��dD5���Aƪ��3�_|�խ[���3`ON!�`mϳ*��Wq�'�}��a�d��?}f&L����#�Y����u�w.Xv�瞻�m���'t�)�q�W0�0�Ɏ.��v>�B���,0z�� �0�XI�A8�O��'�Rv۶mZ �"�CE����ߎ����5>�K&������ǽ�#�������k=����S�������#Y�f�����uB���Kچ�87�<
�X��c�6t#s��[ZZ8��D��0�p�[n�fp���I'�������A`>��3�� ����cOU���-�-��0�������0�N��G?��w���>��ӻ;�AV{��e�8�}���?x����cp<'��%
��q�Ɣj�Y���͛7?������v)w�dɒ���G�|��ib�?���/��Oh������&�U��?�0� �ꦎIQ��m�}�V��E̦8�֝�ޡ�I�F���N�ޞ={81CiކZ��\�-L�%�\B�K&�/ŵ+���r�g�����<����o�M.JC7�b��������=s���,��?'?q�
p�$Y�؎����<���ɒ�ѿ�zKՕT��F���MٴZ��#�������~���/�];!
 ���\p�t �`���Bb5
�hٲe����x�-߼�+@0E�5��g�[~�	�������;w��Di� ����ړ	*s׮]�4�p���,�?X��F.�z��;�
��(��cN���j��1O4�{\=�N�8cF=��2RÃ��8�3""E�"I��]M�M����|���.�c�e��.V�w�G� �D���F����(г�{����IQ6��\볟~�*n>���,^�&��I<OHc"V�)�XvմQ������Ga����Ԟ���Yӵy��=^X՘��wU�»"�i�����]�T���gΗh]�J7�����PY�Oq�1�h����s��a�sLS_� 4P-`l�����N�����qU��b�yX��dI����|���
!��H(4��Y��K*�9� ��w���>61!bw*�Rt�td���,/�A�-�k²?+���yA��
{i<4��ʒ�� � XH\ �]�cC�(K��i�0����P�v��Kn�)��=��H`2�*��I�)����.�	����
�h�~�a.zÆ�qz��-!XK$ v��	7�GB�T�L�H�J���B]����A���K�X	OLC�:Ĝ��
+���iC�b��)	�c�<�JRg�,
`#��zj�]q���U1�s9�ET]� �O��Ӭ���~8�x!�#��#ٸ��E]ч��i+��!QUdɋ��6��3�*y'�2=��c��
Dx=m9��%S͝��ԭ[�zMM`�>n'/ �N&M/e�&��m�Į��b���S���b�E<w��,��mJ~Z3��z�YY�}��RG9�o�MVQ#���`���~���0�Z.z��K��
XwZ�-�� lV�� i��s-�Y"�5�Bd0/jSM=��Ä�s�`�~苺Z�='2�'D�r	QQc��6a���	E��tU(xb��"n�s���h�0 �v�� ')�DW�<�������߹�b,9�*���������z �!�����k	5`�z�4�#M�������"^L��&�����9w�"*I-�c{���}}}��)0�5^�*���2���+����I �HS���ݚHw�Z�ap`�9V�𝸭��A���TNTH��%&���h�ǲet+(������:�m%Se/�
N��.��'�GRD���T[\�B��E.��y�r�YQ�{�.:���)��Q�L�ڐD�EN�Y�\�d,��;4%���+��W���q?_Q�	�ZQS�Re�\�=A�1�������J ������ly��ݱ�vw��s` �A�,m޶�.A��M�8�7��?$�����谋������ȹ���b�n3�졃{���C+LLaQq_I"�P�ӆ��D��&mUK���������AЈ��1|KgL���`M�ta�(
U�D�i���}O5�8ta;|��_y�{�}���z��<���T	֞j�ܵ?b�9��d:�ԃ�����Ȫ�;������Kt�c�<���d	+�ϥ�[rl޹W�����0�O�e�Ɩtj`t\�oP�H�������r{�ן˹⚎r��x^�-����`(���z�W��-��sO;��s+6F�����V���ߺ{��ʁ[V@fIV�h:�S"�4�y�(}��7}�c]yښ��	4�jEĢn�§?�iTD��i��-:�YT��K�"Ù�!֞~x�ӝ��x����-�`<��[z��Zon�6��#K�oPQuK���'.ȵb«1�ѐ���A�7�j�A7�V�1����S���4}oL|��F��Fh܄>r����N��%�a�}����FXu��i�Z���eb=nBy]B��-)r<66���n���茁��UvbU s]P�`Ս��8,0��B(��!taM�V���K$:::t�K��&8!�+��~������`h�.1�`�tU#����^-/�_��:�)F%J���D!������<��a�%��4D�$�w�^��+�[u�����q5��cX�Si���P�������zx��spi��b�z'�х�$;[����IS�z�
�@����9���DZ���c(1��+ŔLb(��I̲;�Fה�=�㓘�k�Cc��ѓ?����X����9'x����F�Q;LMk�y������)fa--X�`Ϟ=��:t���idȞ5khn]Kbd=��K8yU?�����V>�� ]bi��遯Ni׮]{l�'��l�.�#ܬ#��ZRX�(h4��%j۹�{+������tO��:�`���0 �>���N����m"pFg%�K,;D
��|9Ų"3�B�n�j6;ɰA�)p$��"��w�D:�B�C�Yf�ʗ�h�����ie�t��
|D�e�]IYx��Tl�j�p�T� �e��v9�v}�C�u̛7��E�M��,L(�dꘊ�X- �6l� �@��ax��"MD�C�ٟu>���S�hó�k �F�SwXZ	z���S�B�LZ�SJ�0�---�S"B��洧����M���L&I@a��%�okDB��zVX�I#I貈���:����H	���ۙ2j�X������ڌu���/� �L���W�;w<��-B����Xv0bA��ȸ�}� �oJe�`�8�0R����w ��� �)��w�2�~*G�X��۾}����
B�ot�}}�@�O&�q>_J&�b��$��[����HVH�q�ƍ��[[[I�Q��o����|�#��L~(�.���~ƅ�5W_�=!��  (�X�3���3"PJ�닉U�|ӦMK�,��!1wr�W�
C�n`��ޚ5k~s�ǻg�!}(�8Djq[�*^ �5��rٽ��}��P�|��SO_|���7s�]wr.G	+Eo9~��aq��}�A[���YU��3�i05��^x���߿e˖3�8#����O~r��bBp�K�(��p`� �+�5ne8����?��ѕW^������r�-p�/��SY�j�����]H@"o��U1�H���`�H�n.}�A�?�j����)����Ň���d?u�T�}�:�p�sTj����j?#e�����3r��,��!��2d��l�)5攣�kyۈ2td�dܐ_�#!�/���Q����0D�]�%Y<7BOT�1�Z��.#����ԍ�s��/5�U�%��$��Sz�X�"���@W�/����1���)B\���Y�ϐ���$¼%~�B�/��ר����j�����|5�P�W;�C��k��!�:&C9V<�P�5ǆ�Zۻ����K%?���k�u�� ��N��	� ��� �	l��X����9*@B >7$�)L=a����'����'�r��Ts&].��,8N9���qdWʮ��t�9�/�6f���5c���>�Z[]Pw�G~Ll=�DQS5�L�H�puY"v �,���45	�`%]�/�h�!F�8���{8 ��a:�~,��貈V>u��U�,��3��`�!w��g�-C�A�J̛7��a�D��Xn��ݻښ�s�\�o߾-/=�֜NaO��*��]r�%�W��;w�z��e��"���ؾm���"LS,�!25q�z]7�Z'�u6�g0�;���5AB<4B��۵��g�mS4� �gl�x���X�?����k2�[��ȡ��ah��m�Cs�S�\��͗���ܹC�y�@�T!�\��9�&��C�f�o�8��"�v��)��J1�$K���c��`~�G�Z�z��mM�M���zy`�=Ͽ0>8��1��("ѳ��H��vr�YJ$`;bo�MR^���r�ۖ6@>����/b�F/c �f�*?��#T\�F^̤���R�ū�`aG�_���1��4�e*��C��矣$̭[���C���xv
��l.�|�U�H�V��U��]�%UVl�ǁ��f�qI��|n�L�Ud�����f`���+��)	����H�` .�x �mplDȕ$E�}�c���)���y^��XϪ@����7�~|��!"��^Ģ��A4��֖�ѡ���=}ҩa�pvp���\�s�M��;���&��c�H�U9tZ�S�[%WV��K��L¸ܼ����=%���T�	�U)9:*�X�LY���.(��K�����PF�8�iiW���H�&�83�lY�H�t(�Q�c��(r_+�-P������8�ڑ�y8�\wc7��nikb"��$+��a������#1��ɊW�0�*y������fS&�0�nkk��ؠk�
��(��WdK4t�x�%��d��������JK����sL��T�2�f�y������㵺,����pP�zo����O��w�u�U+W>��#�����Fn{\�����l��
#����K�vBY��-^t�O<�jJ#�Cx���a��k���8�����r��e�lX�5���XV�U��r�ĥ+M#�b0��U�c�3���*�� �p◿�-y�Ha��Y�������w�/��R(3_�A�U	��#�p��J]���?��>w^�Sk�%�	;�UM�К�e%��s���?�v��]����]~��Hd�����"f�a=b��$u3p]6�|���"l5�~{�O�X~��'O?�������Ql���`�@���u���h��:�b[�a������^z������L��B��O���/�ת�ƱC�G%�y#G�J8�W�4�,D���ţ<n�xco��#O�6�B�S�Z5�5��Dx�~ʸ��d����Y�\)r��{�꣨���*UE^��)b@wrX3�ܺ.1O�$��vd	��S���ar�G�yZ	>�$�����Z�.���X'��T�JP�L-J`�_y�?�����j�f@��E{��X�^�唉�2���<5e�'R.�ބ��3I�rD�����(x&�̅؇h��k���I"��d(D�����q���/E&�܍�7���r�T4v^2�	�b���"�.e���)a���͟?��'��H�L�!�����=0<���F�E�+��B*<bMh���p��ŋ�q�����������}5m=��]���Q]H�-�7(�(1ŝ4����*�l�8�>�9N��̄���ڼy3�ʰ$ZZZ`�����EX<X8U� 3f';2cHȿT.�`�9X��r�����E]4�?�uM�&\���E��+�r���H�<�L���.P��G�QE7u�.��aT�K�:�ݭ���p-9�.ȓ�2!��� � �1�5^���E���4�����'�\F���l��	a��O�k��6�.�,i����WT�ŕ�Yh��_@&�B��M��D�i�-sJ($c$`Ip���_�?�^�W�����=υAv��ÞFE����p��*�3���ι�f	!#	I�AEP�����C;�8 ����v7~��g�  H+(�̂A�!!	�s���ޚ�<��[���MHhm���>J��R����{������h�H��,>a$�ܤ�2'�������Ƚ��S� n�߇KaH�mIK{/*ZC��-�@>9>nd�c��4p�k�2ܫmdZj���`��H���]�7I���'��_��$��I�G�
σ~�v�H>��L�B�ݶ}��ɽ���[ѠL2Yx�\?�wb�7���hT������jD�\��_����j�q�$��[����!!;�/2�w�(�k����/���M�JSA?*�3ݭQRi�@��Z�y�}�Ľ����:XB^��s�>���۷o_�tI'���g�}�����u=�#,�p�"č�M�</�����<�!;HEGc`.Mq�do��"��7f�̼��+[�n�sĒ�Pmq���!n�}��5k�L��<���@2-?����~ZZ�/ux���s���l.' �4����?���D^,4mO�ML�4��3�&riH�}p�/y�pd���V�н-�Ii�\�������?�w,_���SNvB�t��;�l[М��Y3g������?�y/Brvt�Z��� !����I�s΃�?t�m�}�����@cl:�39�v��O<144�O}J��i��o�����/$��{���ҩ�F���ߟ��֡�r#'�̐��L�ɮ/�9�(�$�M�ߊPc�9*^����VF�Y������,��U5>#i�>[ʆ8�qZ`�"3��?,�b�%?��4�4�@O�d�����/ğ{hB��� h��"6y�/I�<Q��P�99��H5X���bё9@�&�������{��L��:�Ӆn%��*��H�E[���uC֤��"-����LU��ᤕy]�%{Os5T��R�PX%!E:$��F�QfZV���T�m12Od��<��ʭ_$�E��� ��PFɲƼ�����*ѕ��F��;@/�g��������{t'F&���v��[���N#���
B9T#s��t��ɒ�55�f�sz/^�w�#N�׮]��}:!L�4mڴI�f��\��'��Wk��+Wё3�ҿcw}p��q ��a�dO@0H��d5�RW�!�'�k�Z�5�b�LC���0�x5)�u����ي5$YF��i� w�E��H�f��:�Z=�%+�F���y�6n���P˚��~M&�JEd�Db>���ή8Ba��xdhY���n��O2�m�f�P��.X0ur�j>���(6��y�	Gܻh�����wn�{穧Κ9]����k���>�������I�Hz�����?餓Y2��iӝw����f=D�J;WV	�����1�ǘ�� ���ƒ����wwJ[)�iG�o//Yr��c�F7oݳ{Ѥ�z���`[
���f*��Dr=by��B�����.�T�ԣ�ﶭH��4���������#5,�US����Z�=p�q��>eʔ�U�+?���3�H/��������Ɓ�*$͏�؈�|�)�G&Y*�D��1#��r�B��Z,$�w�%_���D6�+��?{�Zj2�[����rʸ�U��k����b�,�z����sVޘ�5��=��,{��ٴF�B���d�����=:·v`J�!7���6;�5��^z}ˆm��u�k���W7,^�p����.��m�`@i/�����i��|��#;���͖�8[5Gx��]�i �Ñ@G�:L���|Xv7�rn��V2s�֭�'��ph���jq�w� ��s�жb���p�YX�r�p��Z�l�0d��h��X�l�(`�T���F�kձZ5�h'IjV��ᾢ�5K�����8ύ#�{�B�!Th���UC<0�� ��1�u��N���҅v:�<��e�j�\chP�ZJN÷*`�&��qB��1��6���8);��&�M�*�i��׽��ꎔ��n�3+�B���<Lo������n�w�,��K
Ĥ���;I��q]��ޮә����zH���m/!.�]d��JF�Tޣæ`�7*t�B��V&��)�D,ռ��n�)�������}ރt,d���\��9år��h�@�6d��I�����5����PE;�O q�_�H��H�!l�D��f�,:Ň2�F聇���h@��9d�Fq�HǜCkU�!M5p��bN��u����T�*�̊e���6i�K�K�v4o)�Śﺴܐ�J��ok���qa\�[�(�A�\d�R`碰�`j�[p��N�l�2�.k�B0ëJ1�t��Qh#�6B<*�,�Xrv���Z�����p�l˶��˗,R��ݕ�_�2���б|�\4ޓK�e'�I��,��D¦f�b�����K	/�b��ψ� ���S����?��K�-��"S�J����ݰm��?=_i�_�� �ѬȹVV�Z��9O�\����T�"��و��i?nڱ�,�8Ee5*�#Mσ�4��+��>,|��qKb�28���АW̄��6��0��U|@d�&;���R����&���X���5&'Dڤ��Cx�����DP�j���9�����n���\pA�h#�G���Z�,U��m���רZ�Jj��q  ��IDATG{��/X:k��Onx��E��0@ĉߢ$3�?��`��b�@�y�G���e�\�/����=y��c�o	z؂�D�����g/-�:>��/+\�,LY�EQ��S1�?�3v���g�9/Mb4 ��_����4�Vp�H�9^-���ʓ���F���ǽ�����J�]O(p^ǰ�у�7tC
����_�H�����Y�}ϕ5�S<�,!�*27$�{���H)dYȹm{�">ĒG��� ��c�rƑ���I������XK���s��H��"R�;_8`�'Xb�>��$=�e�9nҁR]S*!��|��IM��xL=������@tL'�3��ה?>�v��^�'�PCp���)����	����� (YҖ�t)�1��b�_k�(I?T�T47v�@�]n��n~v6���wH���r��=)fƪ��c�`/ydy���TR�{�eq�?k�����ab\�S�B��KU��Y���TT���o�;:h�Z�h����z�,Y�:e*��<������Z{^�7�j�E��kHNj��$��h�"Z�]�7U�UQ� ڼ� C^ڨT*�O�Y��DJǣy����pb�;���+��---��[�^��c�wt�}s��"�	B؊�-��vwwϝ;��ӦM���Ν;�=����7n�[�+V�:���]x��N�5:��������TS�s�̙?~��>��gϞ=y��_z�������z�����J�DHj��{�@䫽eTV8D,BT��|��X"�!ICCC Η��={}�(�����ŜHa���Υz�j�*��7Ѡ�'��mQ�%8QMǌ��4����S�N�3w���[׾D�uc|\�gZ��	�\*~��썷��qh���"ႉ���ӝ��Wp�����X�e52����n�,��&O&�X�H%�'����֤�评陬��Σ)�������k׮�9sf��9�;IA��A���,
�"tj���SkC$}���/X O���zL^��wN�"Ꮅ�<4/�K�d3+9� �]�-�i"��-	"v��@�+��OR���
��y�B	�S��j�<�9�C��w��]:Ӆf�����gIQۖ%&�O��7�t��[�_���$Џ��"y8�c����,"�c��Y�.q��Z��0�Z"	i4j����$�(��M����2Ԛa2�����5C)�<gD*�8�"�N� ����u˩s3'�Z,¼Q���Y^��KI�%�	ų���N0cƌ���Ir�ڎ��3��utҨ��+�b�\n�٣[
�g@�&���|DM�y�%+��j3G)WF��������b��U����fv���h���r�+b}zә��=҂�&��l�A�}����7�y��Wz�g�u6�2(�i��P3#�^r��$��U�b�e_�P���&�I3ЋLF|��s���w���o���S�8���#�>��[�n���KI�^t�E1RUIKD�"
����yS !2 T6��-^L[�< 2;�ݳ�>K����)��
{�~��$�n^$;�$��f)����\B����)V��f�hشHսq�洋�"m5}S74Q���E�3�'Bv���%�H���>M��̥�|�+�@N;�4�3&@[GTvIM_��]�Dw,Z�x�����q�9���j�sH���S�	F&]���o?�S�9��O;�7��C�*��W\�~p=]��?����,M��-�f���ߛHp�d�y�',Z���A�q�2:m��sQ��d�����e5�{�3)�a�8�.�I���rA_dcaC����֒��"�2F"�������O~�&#/#n�-?pHRO8�Ļ7*"#P�v0644o�2Ra��tY�4o�����N2��f��K/����#���"��fP�?����D���SN��o~m;V.�?�9(��P�9O�x!> >���~��.�b�4�E{ \��HA������}���f �������N-_��P	e¯���t�2$��(�������җ�Q5}�]ρe/��C�s�r�6��Z�&�k#R�9S�u	������ �-�r�B�T�Q��*�J�+*���$�r�~��s̀�▕\6'aєm"��:�p�M�LM�fyK�H��y������� �G�|�������L̡J���-�{gM��=��wR�uh]��-����zkKKdWk����d�*�)�6l�F�px�!�K��9�ha�\���=�A+��E�y���:'uw����i�4����pe`���$��A� �Z�i3�._���]��T*!u?�� )b��|�Q
2�H�sȥ����KuL�~q����>�`�ϵG��믿^��͚6�+_n-������|�1��=�e���ێ�?ۘܶ�?�p��fͺ��]y8Y��s'���'�vvv���e�Rk�]w޹u��O�;��^������Ee�A:A��ZT��0�۪׍Ln��JW�Y��ǫ��j5��ʗ�ɽJb:?3F�*�c��|�<g���$t�%{ht|�n	U4rb���p1��8���s3p@�V��2�l���2X�l���Ht�&��L<Q����x4�5Ne8���"^ͧ=��"R4��}2���Yb���
���J�p��@�j����gxx�eB<�5��WCE�	�C+[%_��M������H\�l�>���-��R����4��t
Y������ t,X/P	�r1"H��%�.F��,��-�p�;�B[Kˠ-l��� m	��n鞇�Ƙ�d�nϕ�pi�����l|#����ǲ���
=�z0J*�T�	�MYE |��t���a���PQ],_C-���6��PI�lR�du4d^Ģ���C?�Ĕ��#~��cy��V*�ر�����asm߾]xX�����[I���&���[yYkm�z��5C[����4����`��|�2@�;�H��ӬV+�'�B���q�0ؾaCe���۷��[����ӥ)R(	J׈�?#w@V#:sh~�L�2V�FFWe?��Q�D�<8*"f�!n������a�	CYCC�s	�*�WU-J��=�8��@Y��G��S��'N�_�~��-0�E��'O�����Ys���N���N�f���[�1ӵ�|Yj�/ $\��&�-��A=�LZ�F+ྉ�``�.V��Q��sM�X�a����6��nXdn۵;��8kE�_��;�0u֖{	<!����0ޗ�y_qJ^����9.)��o���y��\����|�I�@7sϑr����I���]ht��N�g��j�!k#�LlM�#��*�tP��[�g~y�M���O<��㏿��{�<������:�U���W==]����h�\��d�V�b�� �DM�a;t���~���?���>�!!!7�t����/�0�1��ً�80sP	P$��	Ϛ�q	8'F���������bM�J��X�$*��&f;���t6�l��I:���52�D�$Bad�9)k�]�����h桇�?tN��4̀�Z3�h�����Q/�sV�y�߽�v���_�Gλ�#��@���6Ғ�>��_P���`�G�z�Ghu��t��0E�*<J&a��O?��j�/=�7��ă�8v�3��:�C�T��O�_Q=�, ��Y�AC:�0t9/qҩ����C����"+����UP��x)�6#Ck�אQSrC���y*`�������<�2���t��Y5��`!U�D}�y�B�7�|���&xw�o~�����a��,&�v�B��%����)]��>$�O��O��8�bo<��V�w���)�)uf$�T�o��n�^ʅ9���\��C��T#HM�N&���"�W��1����޿��7}�c�����ꄷ�|��g���M&�����]x�߫��$2dBfh��x�嗻:&� $T�."򧧞��p�0"�F�6���O~�#?��
2y�������wnrQ���֏^��hѢ-[w�y�I�~�Oσ�IR��3�ت�{�w������n�ᬳ�r\,b�9����f�Y8��-�}N�D����$�b�RuL8�T*q_WD�M��Y������)S�D~��/�=��
8�5�?�De�0�tjs|F���%/�E&�M�s��!�R�;h9"��6��铖�������$��zm�����fKv%�5�*N��[��h����O���5�#@�����ա0�\��a�Y$�Ӌ����>�y�斖�v:-�`��1�WM�>}�o8���Aj>�o�\9_�D�"����i� dq��+���X�e!��˙�(�����@����s�n�����ФI��u4�:DjY�������m������.���0�������B1RĞ�[��TĄg=9[�~�G�c,B��7#�N�饵�1s��t]�sR'��V��GWW׌3Pyeٴd��c�4������F�"��,"$�`� 2��E��3g�l��
�=���c�s�����h@S$�,��H����)kbiH��1|� �q�;��#��i#Vfsk��\/ȉ΋;̏�b�nL�V��B�+���␫�{�����؈W%�uNR�'��d���7�^Ij�[�@��di��B�\�f�%I�l���xBec��%���f$�-����e����Q�_�yQ�md�~7�D+� Z~�`f�δ�SpJ�1�unn*I;�gB0��C�$K&�GD 8�N���2�"�HT��v�t�|L�~Kw�&L�W:�6��u�b�K���Hё�q_�Hз����ά������$�'X4�Ŝ9sH�v��I/Q�ʡ9B rm8h �Jeט�Q��O�Eaj�8��!��Y�v"Io�t��D��M�[�Iڰt?q�A�HxX�w�
�b
��[�\M;� ]�+V�x��G�;��֭���h���!`��x�/���_���Q��;!�,N�\��1n�ae_�ō
��%H��G��^���G}4�1�p�ɫ�����}���� ��
�Bؼ�R�8��'���>����t�M��E�M6���ŋ_r�%�I�h�B��O 1,fu�|L��C�&�l.Q;��I��sqQ�����%\��7ŝ�Q)��&ޙx~q�;@kd��� ܲ-�p?ڽX�>Qp����B���w?DvQ>o��#F!*I4�1Ĺ��Ϋ�%���k���/,Y���\�Z�[o���~���vQ�q��#���_���\���X���g�q�/-Y��&3��7<X2�z����Ue�hm.�����C�k����׿��/���Ǹ��7���R�q��,8$L��|v͂B���9�L�����åRQ��={ގ}����m�v����	����FtGz�=H��dT��aU����J@�ƛ~�~`���vU�^{��=��޽�ז.]y�/���_[(����W,_&�$v~����:��?��i����+����?��5?�ӲTh��OY����К��֘mS�hGA�j���SX��xh����(*������
�&�EJM]�j$�Lh@��70�-T}	��t�k+���kϑ���@3%���,و�}���L�7^Dݶ*9��GqG17L�	-��8ʘ̴;22uR�SO�[��PIu�Y-'�ZYWL:y����q��n��g.c�_:}��X���p�Y4���׾u�Uts���&�%�TFG�WMh���&�N#��gR+�>c���-v]וO�������_��0�ޓ�X'�l�a�*�d�b���o��c�0��!��-1�@۬��;�n���\ߐU�\�!��v�۱2-g��w �{�����R��������;�����rkq���(�h�5��᳜4�����b��8�[����$#���q}�^��䐮�R袃�-��:a��݃���oݶ���r{'�������loo�n۹�QϊSDX��\�Mr�7��P�$B��1���Pmt���֪�ޞ� c7�lg��e��T�Z�lݲ%�]����oc(��G�cH��*s�M�ڿs�26\]z��s��|1��<p/���V�c�35��B��V�7���;ц��	�A�5�XFvh#�%&S&Atٞ���n�A�)dj6Gȳ<����xD*���U@z��ȾB �$^�~��ɓi���Ff̘�a��f�2���D�*i�T�X�3�<���,x�wlXw�a��f�6�����K�6�Ȅa.�U9�l��?��-�aq�#��E�2�s,s� W	a�ā�K9Y�r���Z�B���ޅߕa��ش�.�Vn��[�H0ZJezu�:�.S'O	$9c��*RB���Ey۱�N������O>�=�Jh��][GG�-�h��C�^�[�wJ���7KNCG]wI��:�st�@�>-���D(�6�;���&��1�bL�XTL���o�N���h�0;��Ծ�?Կa��ws�N�z�N��I�E++tp�6��}����K��]�\�k_E! W�r����C�l�A2C�"�d�7�fŋ�n�;,	Q�J�cOذk���?_��gH�?z��i/��ȕ�u��r�ktmJE���@�/�����?5}�bh&���&��k��n�B2����6oCt��=,�Y����x�1F���!k�m�rd���x&L�K��ǲ���?!�Q�Y'�e2��8)='�t�N' yx���ˬ ���|n�)"Zb�(L�1���~r�LS�0n�Vn	�Ǽʀ��|r|�MR�h��]����{k5H�nAvw^%�Wm�G�x($É*��R��bĲ	���l:'x.!���A�~���R�������t8�s�Z�u��L��o�L'r��r�(dZ=�#��$*(�G9�QR��sQ#�:�L?xr"���(��0i�|�dd+:��]B��V/s��W־z��r���4�W\��o|��k�.��������"{�������V[�����ѭ��Rd3����ŋ�������H㎞�>��{����a�j�`�v5�^ni�-����u��2�ͼ>c�̝��>r�G���F�7��]�!
	Cζih�J@K
5��H���nJ�(�j$3ɄU��F��i'��SX��KK&�4��D��	8'�(��490n1&�<�;���h�L���_���/8����ǴA0���9�^t�G?a�s%J��hٲe0E�Y_+;7l�@��UU0�f��"�����
�������Q�;^\4� tc8>����������Y�S�P$��tCAb��_m��G�^�l������dɒ�;Gh���H��|�o<�ۻ|����|�~6�m����#_ST?��z+�8��[n����x#�C�`(R���U�V��S�<���:)a���<ayW�$��m���0��p�q��B�*\�on �7�ڡ�z�5�|�3����~7o�<�d��W~��/_���P!�=o�����g���O|����+W�B�P߀�4��h������Yh���݅D�_OEW�Jc�{�O
	�MgDn��4���������Beo����)�����}©t���=����_e����ц\}�	d�r�)4�ϱ(���~��g�<�;��/�я~�O��O7�|C�aq�d�f���L-��'���'���w����qǯIUV�Q|�[W���k������9���i�'�����W^u�U�5vI�����/~񋿺��4o�^�ձ���E�Mw3<o�����[o��駟�v�̦�т�����`1��y-|`�L
T�� A����<�����Gy��EЭ;w���Xn޼9k���?|��cO<�H,U���a���,��%�n_X���O?�?f��V)'�7W�  ^���K��h֬Y��������6,������Z:��3g�%��ݿ�~��-�tq��%��;O���t�?��E��Db@v-Yt)Bw-�����Qh��x����� ��d;��mۢ̞={�N_�`���ӻ:;E!�ĩ��JW���[i���t�Μ�}�v׵�L�B7O��~�zB,�f���m�8N��� �lı,���g�y��Mo��&���}�|��;mJz�FvtͶ@�hj�j�d7�x㆝��v��ji!���U�A�v!F8.^BA=�f�c>�cQ\w�]w���V�Li�i).]����'=�f��'��{���0Mn������	Y�4���vD�u```hd�����NcGX,�/:�&I�p���������Pa�<��"�~Q�3˚6iҤwΟE�[v�J*��m۶�gf��᝱k��1	Q7��@4�p�6�**
��i�A��x%D�ƃl�H�c�B�m�O�B��,��j%29�@0Fb݈0W� �zRk��מ2�
?1?� �����o����@\�c-���f�<����̌�I>��i�F�FI�}���x�;~��?�=��сТՀ%���Mb���`r�&�8��� QFL�=�5� 6<碋.*��н�v˭}}}"�����B4(��k�R8ڱ�,OhK�4�i���N�*Ka����9�gA��
����Q� e�k�n���s��F��E7�D|�>�Y)B��J�@���'EOj`G��Tn�'4�hk��{��/qɬ8��ۺO8ᄹs��ٲa�-[|�b����iqea��M��Uz��Ea�mo��It���D��2I{N�T4ǣ{����0{-ϔ�۠Z$�=v�_'���d5I)��W`��H��
��K�g5�1@t��x�\���(I����I���eq���u���a5C�P�T�^�������^\�����Șd�"�D��>.���r�{��\ ��c���BE���[�[�,$UAt�\.ZL&D�-�l����%u�bs�qT�(r�&	�DkAi��Ǌ�`� ܅��&�x���f��Ĺo�=E�;���������s�쩲�xe�e���P1�n%���!D�����)I���T���a�b0�"�!�q��[�_Υ���E\'�X_εɘ�(��Z�)1���Hg{���ϣ;�c��=����_��Rt�Ɩ�]z���^�������ϋ�`�ڦ�}��8F���y��U�� �g��(����Ɉn|��?��ҋ�\����������ǯ~�4��y:���F�N�=!?[)���n�"��~]%S��Q>$�rI����	^�c�H5�*�E��y�$�$b_��9:�{�Z�����j�U��5Ѵ/�)o��DX����� Eb�	W
<�L�|��V�L�*]�W�"�L���쩈��q�C�$�¤����W˱	MA����;�P?��M��A���|N��0r{'w���<�������l\q�!t{�m��g�n�Ҙ��.��Z��Wn޴���x=�n�١bjr�D)I7i�ۧ�}add�<���+D�-:�4ݸ��������e�|��8����n��^y���ŋ���Cw�j>���������\C:��;���w��$WH'����.��_��?Ns✇�q�-���hP�&�#�nM4|%�RGiі犹�B�TH+�� R1���3:Z��b��/����_�gu5��1Y�����5*�C{V�^���m2��]N�q8���%���+/����=��l�z�$�I�p��y�TGq��^ym}�>�-utuu̞=;_.��6e�,Z���$��JcӖ�������j�:!���,�<IU�D]Ď)Vё�8d�8$.;��:�^]}�Qm-�c}}���<ȗr~D6�ভ�^XKS�6�Y3f�d�I=m����7l�m;����w�{���i��{�l�+�?<�m�����{z���)^��蠫W*t��C��0���>�U��Hx����b��PNAX6ٜ�jd���Ǩ$�ifH��.^Y���G��$�Y�����7�x#����![�e�40�h���#~�eԺOGZ&T�!�̬m[����2w:͒��0θ���)B��G�i�RA����o�z+�P���s�%At��I�7��bN��|u/;wl�d/�,9��u�vf�U����P�v��$�����qJ���Jvt��^��S�秩%�\z���xy�)ee��=����Nar!3�TZ9G��{9Q��'�6c��\� �ԉ�,ϧ��yH�ɣ�0�~5�H�a\���e޴y�f&�ɛd���b�"��VaAv���Jo�$��-�����|G�$H8G"և��q�yutQ*I@���ru����@MRS�$�������˨�]�1VZ8o���g�v���4�'�}���k;
�V��s�'Ԛ��h��LZ��k�xx�S*v�)U��ryԮ&�:{ֻ����Z|�*�Qi���nYtP��7R4p=����d���!���&�E�,&GSd �"-H�
W-\8u���	�R�×u����2��a�HI-�ʀ��|DG��D�����k�+Hk27M��P�J
���S����J~E��!���dr�Rk�����X�F��:i��WN���QF��`��1��}��-;w��I��lwlp 	�_��9|*����$�Ș��Roo�ys�4���� 22Vy�Gt9G>2�L�ƴO��
�ESg��ݪ"ڎ��ĢS(���z-T}��q-�MO��م�Nv�*�X�u��#�~X�[�No��au�B�>g:��ǎd�t�M�U��`�9+��F�E�@�r��w��k�:	��PVg��pޗ�[��
�M�8��"
�H�6�TCSy6b��q���g��.�KA!f����$R��Xe�? u��)����A���4�P��4P���6��fPHK��Q�Nc�� M&$m�YǞ`;@6$�k<]��$P���������4�C'�mqw8+�>��Ȥ�'����(d�p����Z5���M���6��e\���
"�6�i���l6�=�J1ռ��_������躘�S��W7�^h�\�����5�(�@��������^{�ED�|��@�d�a6�ht�s?�o���C'�&�j옘��m�>�|����O�Iu���y͕[�����;����U��w ����߃�����#�6j؂@�v��)H��qÆ/~�n�t�I��=��CC�?���-��=�,�J��o��X4=�.`�٨�G9
]�X,2�$�.ٌAHB:8�J*%�GM��Vl-�/H��`.Дإ�[�Z�`8�]Ļ�D�H�d3Y�/uӍ7��Ծrշ�<�L)�ќ$F� N0�!�7��ɚ72r�.FA��t�]�שʬY�2�כ	i���쬂d�r�-tT_q�K�.E�?r��\�׎��Sg^u�U���gh|��_�I޺m۠�X.�,�!Cd��w��>��={��UFK��ZD7�R!����N����v�˝&����h�_[�8�v�'���K�Q�|�➞G7�8���N�s#���Σ�:�W^���U�uN�v^{��o���/�?t�)S����B�s��m۶�Y��g^"볣�M�Q�T�t�Dֻ�pք K�o�_���W���d	u�tө_(�aU�[�C���߽g���o6M}o��rj;�IٰSeHQ�a&�tWr3�^x�l-���|�;_��[7�;�tO�+���O�B{{,� �Tu�̙,xn���{���G C5�z�!�m��e�� {��×�o�|���۷���?9��_�bW_߳�>{���O�<Yo��PB�`x��9x�:�����Y�Č�덆-��)\�������� pVE��m��#4�{z���T��t5�p�x�1η��!����D��B��B_��,w��ٞ��2mڴv�NJ�[|���\���j�Z~���+DE��&ثLD��>ǑD8#�;�=�����ª�ѥ:���,��IDd�����˷aw�[�˖,�b0FS��B��vl�V��Ix�Q��
c��������q�I%lx��з*�x�<��Q���<=�{f3I��~\���b�g��6�|�F$d��]������xӦM�w�loo+����s{1ˮ34�I�I$0}H��eJ�Tv	s�/���	v��L���[�>���O����m��+W.[��SރnT[7mݴ�^̟?7����09��MO�qo���|�4?|`��6`�A�� 4Q�Y.\H���'_z�%Rb�/f�����������e[c�	1c>s	��W�ӤW�UR�$K4?����$�n���	(~�`S�8dh'7���8��ؘ#I4"�ŝ,S\�lF�r�4w|��sz-�#��d�z]�K�O����5w&��c�=�X��8�K��g2�8�y�c5D�#����e?W�A�x��f�.�����իW����o��v�E���+�[���w{VL��c�&ⲱ2=�3ǩ�<�X;�����AC��L�~�p.�g���s��� �V� ;��(�@t�u	5�Z>�g�F��T~Ʌ�f����JbE�%5KCu#�(%1��'�l(#6ž´�I�%NE�r� @ݚaj�IOKk�Y<)\3��%$6���k�ז��4�URiVŋ�K��c�t}a��M����KU��x�&P��^NҔ�7˽Đ9�Q3�܏/�ˢ�З�Z��A��}}�+��D�sج���]�s��2\SB�I�cؽ1��i�bǑ ���*PG�*b���yL�d�~�N���Y!��q12���Fù��민�JA%+d��l��ح��k�yFײ�R�7��&�H������ltɦlZ�u�)���h9+Jx��a\Kj+3]g�i����I����{��	�9uX5N9���W.�-v�+V\�/]w�u���=�c��Ț�}|p�ʕsH:��{�|N?Ț9U֜ 4U-��� w���&S?G�$�N��!��iaZ��^G\<Q�`�av>�5|���ʹٱ���!�I��8
�n�F�u�g�
�}���Ire�3^}Ԫg�z���(�ݙ�5:���@��E�{+�6o�J�ާ]�B�����@�I{�w�X�Jh���3L�(���N҈#�E7Х��W���[��'��-@O�X���ֆ�ĭ��c?��S��vjgW��Zp�	V%P�l&�8Ge�N#�8\W�!{�'<9T���%�/�ΰ8�䔏A�TU��:EY�oK}��O��������d���B�-P�gۓ;ڬ�����[�d�ξ!5����Y4�͕�+&s�
�q�r��_9���g�\/��$��*�ˑ�f�]�#�|e}_&���<�#cc��G� ���V��e�if�1��ӆ�Z�s�T���vk�ɥ���8�.4c|h��_܄X�[�b��~^VqJ�5�a�"�ձ��o����Ki\#Cc#��ƫw�a虗�
��kd��2���C�d&���m7���ɕ~����#��1<<�y�
�t�W%�+�e�Or����$	 ,���B�WĩOV�d�,e���D�'gң�*�cR'e�	����"��F��k)��*ٟ��]��+��U��c�Y�E`�T:���mS��D��C>��4�e$�m�g�s�������ٿA���Ii
�=ڟ_hM���]~WK)����Cx~��=�-�����u�Q��ǫLǆF�:��hp�`�$D�gϞ��^m�	M�T�gg�/��n�>+��Yw����\��Ʉ��"Jf��;vݹ��дۃۤ9�vf�g��E����V��G��dY�H���W��"PzhYS�n��5�j�Ch	t��vpO����8�$�T.����v��'��w�/��D+k���n�A�AF�I#��v<@V��حm��-�r�#lP�EM�n�~d� ���tEe���PaՅyXr%�*�U�G1��}.bh�~14��oF�+�lk���n�B6��S	�n_��S4�0�2e�ǐ\��7�����l�s�q~>pꄦ)Y��ð3�V��!RN�ڬ��:'�4∴�j���U2Z�%c�����hD�7B�ů�W�����F��Z�d����Í�,X|�60Y����n��B(��z�q���6)�t�Xud�l�:J�����1�l)J����Z����L7���J��'�"�2�Y�fZ�߷%@�%��!�uG{qiȼj��h;��Q*�إu�6���*��W�|���{��/8td`ޙ�����c���b.k��=���HkT�s�I�-��;ދP��32��O�������}���g��t�۱cG��Ɔ��~s�m���c���}}}$�d�Y�m��U����s9:0,�ͨ������]�g��k�`��4}"�C��m�^I�N��]#��(<d�.�cFTT�@2n��!�V�
�H�d%e�|������c�4VZ���E��4�4�c�v=�TZMx�9��b�q�@;�v��Z�20���E��k�˩q���Ơ�[��q3�TJzM$���|����f"))4���~�䈴U�brNW���:���e�&�S���s�$��3N�Q�eLŷA����,-�@Sk��O3� �3d����bxx��E�<Q�#���]a�3y"�
v��b*�D�#4%��	��HD��j!����6M� �K�]*#��q����O\ �=3�c�`I�S�g�g,�i�_�G�9�W]y�����ߺZ�������7�^�H���^����b3ʡ�'�}��_w�{O?�5׊C�n�%<L:����y�l�F�7��nF�I� J6�-[H��H����%��x���uM#o�	_/����ӟ�w�Gc��M^�k���g?��%�6S#���N�+|�+���7�H�h�jK�����{���-eH �4}<%��&lԔ��`�J�A�	)�R�"/��q��ݤP�O�xY>�7l�`�3����wĮ1��Bɐ&�Q�*[
ǶW�G�P��+/�ڽ����3.( I	�E��D7dz�?d�E1G�������E�3�:6�w	$������/g��Q�Gw�u��];�=�ZD{{;A������c�ݻ�~��؟�}��%��	�eo�x��4q��{+
D��Rk�v��/��$���D��{o���;�\~���3����x��i ��1�6��i.�6X^��H܅��q*�L:c��d�c2�+K�)
23\y!�ǂ���P�kx��S�Q\�!),G*���"�`@�5�փʕ�#���֪�G�f�.�0�+:�(��õ�<"9L� �=����'����ȡL�g���$x�82�2V�`ch䜖t���Ҕ
JCQ�$D���u�*�:���(7[�lQ�L���02�`���L��u��CE*��%���Rnݺ�<�	��H��o���&ً������f��"={�}���A T������q�Ui�#7���
�Y�7=�:$r�gH8�bsנ��v)!OI��6��qݗ3Zׄ�&||����VZ����W�
����̙�m��Հ�(��x,b��N�d�9�f&�kmmE�ˣ-��ꏍ��!����\,��]9�	�*ȿ���i���W]��!�qB�y�8:!�4��t�0a@b�����ʉ�=�� �����1D�s28�|.�E�z�U����
·��I8B��]q�r�3���O������H	

rHz�{|�ꫯ�󨳔�wh�Pu����J�m%|���S�=�Q�ڽ{w�����ˋ��]]]����hݻ�LEhs`7I��w�KRDӅ.s�
�s���>!F������Z�lmt&�~b�Z���L���e�����GK%�;�
�']�ǼIb�j,��"���87O3�8'w�Μ�@�"�!��x�1�R�_Vv,|7r#�_lm�mi�@e��R�^� ���uk�N�wv�asg�\�f����;����7n$�LZ�)���p @I�i`~E����a�JD�	TO�6������-账ge��c�=v޼y�=�ʺu�.ZA3y���!=3��;���q�ٚ�*�R�Vd�	O��&�.�(���P��PY:�e�$�I*�N1� E䏩��!-鞂z�B^[5>��h��_I��G! J�i8�6~(>�t�J1%
�/�)s��'�NXV:^���,��m&�A��	�U:]� �	S��SM�47)`�ܬ)֝p������eM'Aa�"�������A8�>E&�TSfO1@�^rĽ���$]��LZ��Ǜ�<���O�*p)>N��f�1��ILI�t5�YJW�18�t�I�C�-w��bdP����Ҥ������~�7���o\��k}�;���w�{葋~�a:"
�}�Z���"��n����y�e����8W
�޵k�����!��p����5����m���G�I#�`�y������3�fvh������[�s�Y�F����EϊoO�6yhl�������:���'����9��^��)T�(!c\]*$�y��_��
m�M^N��Ns��B�/��u���Yi�}��2.J����t�0ƀ�(hjvhqyGs�O���|��y���A��;q����~��/����bT�F�I'�t�������&��E��"	&���𒥮�%_��<�j4�z`�j��`�k/��<�R{)V<F��J^k����3��U�����w�w�O��d���\�5k�ǧ�x�w��3ψBw�٧�tݿ����<��C��0�җ���"RĪ��n&�6zSA����vg�����n��"�@�8�g�����Uo�J�o�(��o�\�﵍#���L`��%_D��ؔ�E�=ٝ�ēU�sN�h���6&ň刌G��N犊��z~��ISE�:VD+j��3���cɗ��'���#h�K�(�}ăH��'�8�9� Q�ɠjUi���)��/r?9tI��/�ff�-64�C�r�N�[�@<�/ˁ6����-�jIA�6d�nP�2��-�������y~[1�a#�L/h����9À�';Hי�DQ��x���-�~47���Z�L��9�-�3N���8��}؊������d�}�l(�1��Qlm�c3�N+�w���e�pҤIB��E�E"`�-}d>����f9^&W�#��e����T
:C�uM��Wפ@KU{���8�&�ߗ�Ya��=�~w�m�:��Ic�>�,�b!��r{�0*�. �(�1zh�\���"st�@7jN�l�(J��wּ�K"س�;�/�TepTc�~�	�H.KJ^7úk�~V'Q�
�\����J�֣F�!��qM�	R�fhլLa��ٚl�}ڻ���$���r��(p룅�<��� ���-�Ȳ��x�!ʩ�����6L1���`��1sTr���ɹ
_��itvO"�J�z�<N�>��V6�j��˵%�fn���"
���]plc3���)��#�!@(RF�8��C�&�888@S���5u��p��RRV���?�7����س���%�H��G>�ARh��\�"�Jv�焮�r�]�������;e���=ӧC�3�y��[��-�)�$&�	Ĩ�(W(Z6�$�MWV��)W}-���m��j��� �Il��k[�gՔ�R���Jml�rI�Ё�s��HWb��h;P�=se44͵�����ad^�Tj��.hkS9{P82�v\���l:m8���A�8sw�"!sY�MVu�G�2mʤ���(��Fc��H���/lܸ���?r��_~u���W���sOӧz��59�:0 Ё$#�[�܀�8��3���ҮY�~=�y����m�j�F72�mpƬ�GuT{1_�=Έ|�28��Bkэ��� ���a�d����h��c�`��B�`����r \98��Ic\r�?�"�Kʁ𡪑�x�&�	O��$��H�
��Kߠ7�0`FY0
$���|8N�|i.ɉ��+d��f�\��~�IͨQZ�.���m��Du�̽#qVJi��sD]"gRLܿp�(�&:a�� �D�ҾpK�# ��'��Һ�-.+7;�����Hr����I�eD�
w!b�Q��+NB�41�f�b«��@aU�D�-`�j]���3���^E�@U�6bH�� �WSp�g�Z¶*"�I�R�aYP8ﵣ��5�O8}Q�q�#|�A ��%Y���h����5�^��R8�{��Ň]�9�=����/��׳�'[ɥ��8�>Zk[J�����/@yUM�5���W{zgut]���ѹ�A.�3 �b�p��m����r{W4! ���u��ϙ=���ξ���=?��L�'k���`d�q�$z�<���O���.����墂�Sb���D�^r�� �~����^D��	�W��Fu����#<񜪑�ՔrTt:�?q3;1\-Ҳ#�~'�p��?�~)�
Z.�\�F6�9mM���p��d�(��"����K}���,��IhR&t]?�1-Z�FE�m�����Po	 0���3e����q��5H���'?��.9��S�������Oh_�җn���z���M�ѫgŒC>����>1�*���������	�a��*PQ���� �$3[(}&.O��-����Ec�z  �P�A��(��Gl�R�7��u"!*�7&�	���XhT�?@�C�3�Qd����kLC���T�jM�P{����ѧ2�]��b>`�BTA�A��.f�����bYI��b��SH�C2�9-6\��ۖ�<�DHO�8�N����p-���EEN>�z9#J�!*��"��Аȳ���s�qHò��4{�v���e������&?~z��+(\-8�������/6#8�x!b�L=���'��a�j������5�=�$��V#Ց�r�?�M�xPIn3J�*�H��\��G�D4O���&\����v 6��w�4�DXR�a��OToook[n�n�/ڸ��\(H�9�~�+��XŪ�t���m8��PJob;����X q���� Ic{K��� ��ՑJ�K��9sH�
�����+�"�l��A�N�f�ۘ����T��8�QR�"�W8�)H�;j�x��5\!�����!��F�l�t��\Z&���
͐��ƵD!p��I=���
��H__�h��tĐI�!����[Xn=����A$�'��i].}IE�wiFGG���Q��#+qdd�6�Z55�#����P*+lG�<����H'�cEAww�Z��?EtNoU�q^~�	f��
���
��&�4��s�HQs-��H��f����Ӱ퐬Q�=�O�>=j6e��L(/pD�	��AM��٣눤	��qX'K4�xG�/^L��� ��	�ӯsh��y�	S���&�b3'3m=}��T�K�,���Syo/�	�.y��]���T����0��D��apG��?�͊����vD��i�)A�W��fҺ7-��E�i��lR�<c/��,�K5mzOx?9�SЕ�lHo
���'�E����+�Q�¹�Ir&5���sF�B�٠�d̹���Q�.Jx|$)m�̛`�&��kip�JL7�_��	U�h����8 �4�$E8��懌�U�R��9���q��jDt� *rm0���w�E�X>o�v�Q��)S�GPs�ޏ\����J�S��J��uoL�>͎�,hY�W��G����R3��aÆ'�7J���gn�ܹ<jqP���6@O�й�͛4Յ���;n'Pq�>�����)u����a�-ʶN�ӟ���L�`X���U+�>���{�G�Ȓ	�8�̀ɏ��	�˄��s�@��B�"�4*R��Ja*�$:��k뀂+5-~a˦4�	m7���b�5�sm	�r,�Pv�l��#uvwUގ�;[�j\w�%M�����/yo'YU��}�����=����3( ��	&BE"�Q4ɫD�O1B0��F��`�v�Q�Hd�Ł�azfz���ګ�~����[�53�o���i��Z�=�9�y�������Ԑ����O��f��T$+#}����s�9�s�:*��!�d�F�6�.�E�%"�O����Gv>�D��G)��.p� ��8��d���=s�o3׮�2�������׿�w���~��B�h*�a{��;w�;����w������O|���X	R��W������F����"s�>Nc^��T�JY�P{V��7�}� l���z4�	��Hs���Z�06
69��O.`��BgT��f3���-��
>w�%�D>��2Pk� 䃤���,J�`�r���5���S'���g���&[�����>��f�XT�xG� ,'����s�O�G�����fQ�駟���'�|��%��D)���}���1�ɍ�҆��|6��Q���,Z��9���������	��R�%O�D4�(�O�-c�B��*I;��������i�"R�������$>��C�5�ޭ7,C�z�N��h
Z$XMcr�52��dvfz���l��������g��*��{4�$0�&|���  �D?���^����$�k�ka����h=�j_�@��;W�(�#r�*��]� ��@:��K�8=7+qH�H�_�E֟bf�z���x��
?$K)	t,[�jJ�Ç��ddD-�&�ٺ$'�"Zt[���{������-/��5�dh3O���:���{�����}y�F��F�ZrnR���t�0�$��=�I��B��]�z�j5�JX�2jN������4��`(��H�H�"�܊A&�G���쮦��m�hEQ��[�M�q6;pꩧ��'e��린�hJ-����]���$�	5np3�ɘ=rc�d�_��H>���k�5�
B���c�>�쓿}�19��o/��|�͙�s�+7��<33s���K_��o~��}�1Bm��&⼖_�'�P�f�R�^�6j+V�Xr�a]t��L��4�l0��\�7J�Ү����w�<Ȍ]���m��{�r�}�_�944TX�/�o��5�VoذAg'��M���k���<����o۶�?��?�B��ם:�j������%2�����NLLq��u�����]w���Ds�Ӣ`՚Uoy�[�+�v~���ҿ����L�v@�gp�t��Fa�3���?/BQ��a��p(JGy\4�K��D~}�S��[.�늢�Vܾ�^��J_!K�c��4?W^�n�����}}}�76=�Bǋ&�I������q�(�f�4W�������D5d9�h�\�25�ݴ�k�m�9Ǉ�_��sc��`�˓���{GFF
&Ω��xe||�Į�K���ȣ�1�<-�~�4C�Q���3ID�Gf������	I��o��,��
0���G�
2�!�fz{� ������&p���ґ¹Øۆ䶗��&#=�q�9A� ��dַ�0�hKu���{9��S�-u��~H�E�A��4R$�"=Z�U�k?��R'���W8a���c�uz���<�*�iT�����4�H��\��P��j_$���
�P)19�`�&ρ�q�{-Q]�Q���9%��"�	�}�p�0IK�`{���uR�G��A���w��J�Ռ���D�Q#�!�YQ�{מc��p�)�|����!��!
]I]q����R-[��$Tt%�Y59F�A!�#��]703�/͉��h����\��[?��m���qj�6�O~���Ëi�(dH˰l�Xz����yM����ʧ޸q�>������>���]��/��PU��~��6o�|��G�d�k�����?N�<��Bb^�(�*�4݄6L��.���Q;��2���ޠ�KqbA.��b�L[!����U��s2\>��'���o~����M�w���a��'A..ޏ�i!��L�m�~@��@�	���IZi��g���;���6l<����Y%с+���{ｵZ�MoxCƴ�8hT*ټ}��?��k������ܳ���?�uU�И�lڴIpM �'	o���C9�;%<�>'RD�Ë��~��K$m�5 �`��#fY��FcnV�����#9�8���V~� =b��M
��X��I�&bh*��dA*�!Zϵ|��,�����v���YnQ��i�}d�4��{���:CJ#_�}"�?uQ����wŊe۷oo��S��N	�׹=3,��/}��7(s�Iz��I:D��!$F(�@`/��A��Kϻz���%�9NTc$�N��ܒhn���l�g5^�=9� ��C��=�@-��0@0��j�J����!A 2�,���4��?MV`���H��=���Vد����)uE[E'�L<;;������sd5r��@�:GpL���K�P�w"^�0u�s����,7���yOj�w�A��G�M�,��6q!*2?�8hh�*3����2�L��wD���He����uF��Xv)�,�֚ڙ+�@4 �}ݤ�����t���\`��XD���2l��"��b��m h�!��BW�K�B�T�4e�2����`��8�J/|���^H(�����7n�HMMM�ܹ�TG������m��n*��ޫ��]&z��U��&�*�8��_�r���,�>�}�R�v��#"�&+[�D���5h7�+�GD�������^�*�^P(`$�˝��N�U������=�@���a4�,|-(�C�~��V0���-���T��~����Yv8�&�����)N��RD# �'o(���(H�!-��e��{���Ҟ�K��}.��� ��=�E��˗�)���V��$��*,Y��0��-XU皂}��PS^H��La�m�,� �R���/1wՊUf?V&�"J���ueQR����-��;�?h����������u�3:F��Ra�w<�;c���N.-<ؾ���%]~JW3��O�O锽u�@a��n�"/�ZwZ��}��?��-4�F�֎�K!3�Y��ܾ�6d@�FM�����U��\��r�X�]��dI�&)|>�:���q,��`I�n��}�Wjg��X��l٢�\�O��c D����v��~����;���P��2I�>��c�~�Go���H���.��ϹKh���\���Ǎ����_��|���\q�G葏}�cw�}�����6OC$3p����JD�E�_��
5�XZ��a2�2�/��ү}��^����G}d&P�?����o8��_�����yR$V��}ő{��_�N� ��<L���~:��N����(�K�f*Q�!�a=;d��؆�;/"������=L�C[ZPoaS%RG�h(�:P�O��e�]�[�H��Mo��+?�fŒ7�AKv��^"fk�e�6]�R���-ײ%]s45�z�}U�7|3���(�#�ђ-�TT�05���k��Z��o.��_?����SO����l%dJ%�:�{q�n��OW�k$�~��#���\����O}���t���gf��(�H�8�V������}�����~�sl��K/�9�)�4)�jM3�kϟ �y�.)*/�p�u�N�4Y�&���Ӕ������T���S�r��=`��$Vc�o�d���8���"�Kпe��d�E��D�&ʲ�jP
�HƲ�B�Q�qUh=Eb�THr�O�k��)#�T��L������իWr��\�S�$����D����դW*��u���;�N��H��X�)C�M6T�
N��c�ڰ�Kd-'�qLI�u�N�-J���b`,�-�i^3�Ѡ��]�e=p�%Cm�0rY�@}U�N�Z���1j�pq�&����5U���6o����vn����'j�
�9ve�{��|z[����F�����
9��s���A�4O��{^�)���"�Gp��,f���)�� 7@�)>ꦲ�>R�}N�E5�VfI�~_�Z���,�O
�� -��'g�m�и=Dl�}�#��g��'ɾ�����r޺��1�>��hv
k�ڶ緍ɺU���4^3=W�I=�W�1��Z�U���
������wd�Ỉ7jZ��#�1_/�1�P�j�lt,;~+@�1�C������ �6BH�vV-�c�F�&�y������&�Wg,CFȌL՛aDƷ˝�'W*��#R�f�JAت7T҇u�w�>����uk����ɂ�M��2G�C�k�|���ߙCt�ӛZ>�*�9��^��W��#C�N_ї��4t91�r��x���N��ۻwo��7_(��Ѝ�MWh'��?q��r3����rE�څ��z$�����mW\��L�����w^B������={�|�_�yٲe#�T�r�20��Y���P�v�\�Շ~��y����{G�gh��eU~�gf˥+V��MoRW�L�����8˖�S�?O�ngiv͉'�u���_�~��c֮]��7�aӦM}���U�f&&�(LUw������w��G�OO�OLl߱�\����
y�Fa��������@+����k�$(�U��V�	E�� n��-��䅏��Q�>�l���d˯�?0>]2+�:b%A��w�Q������&��#��mXC}C��מ���Ϙ�-��e���5I���S̓�ʳ�㵹��^}2}��=��`���y��;��_4��槞��\��|�߾�#����Ç���#?�_�bn|<65%Jt��`��a	�2ѡI�kKV|��0����E�MA3$�:9�.��4�DD9>�4\&'W�u��!ꊚn�����c����1h[1&0��I�
������%i�̦Q̞wX�i6��;U�ݾ��Q����>�,�EJ�S�`&Y��v'�-��h��������`uA�w>��;Y]"����2��/�ƀm*�%m���Gƞ��y�TKB�(��N:sc�F4t��셾%�_8Ԥw�$����/L�+*JɵLR�Ֆ&����'���^2���̇~�������p�Fd	�K��_������_��&�r��\4����?���A5�;�/'���ŭ�W)��s�-�42��WS��<9'��J�}�E����>���ҏ����M���>�t�"�8"I����%w}q���2lv[m�Y�fͧ?������?����x������Ǟ~��뮻���_p����C!��~�`\������}�$I^�*��D*mN������퐹HO���:��%�-ю�	�����wǆ�[n˰P��ƍ7޸�g���X�o_��������#.�b����i�9ϐ���`�'qo��u�r�1�{K#�(��o4�v��XȂq%o��W���SO=�/��/o��;�P|�t�W~�_m�ַo�q�'Ǧ�z�W���O_����~�Y�!2l��j��
���ŋ���~�����i�h䧟~��ɼ�o�`�R�Wz��k��,9 Y���N\Y2�Vx�<w����2��d�L/Hk�@Ǫ1^*��LFj����J
%b~,�y&�S,��) �3<W'��R8�.�4]f���̈́�Aa*��x��D�w||�m+R��"����$l���i���N����0z5����'�,�2}��t���%�4bf����t��-�JW�
�yK鷺��N�BC�7�x��hZ�Bv	�M&��tR�iΡ���	,Z��:�~2��f+"��z����#�#̃l֪e�OE�Ȩz��8��l���wԉk*�BN�{��ޮ�AgI��ϣ����9��Iܾ����g�����F��͉tYC�<#�g*)k�U��HOOO_]:q5�Z��>݁46�"W#b�茊�P�~ ��w1ʰ)�BoА\NZz�'���{l�gmpI�m�9�4�����2�T�r�������I{��6���y'��2P�vPe>�Rv�U%m��D���k��8e��>�B��	�i�)��h]#	3O{�%+���24	4~��MO�k�-	�L��!�p��	.5�Lo`ڦ�v��2�����-�h3��=�c�%��޹f��Dj�0<<L/+���+W��Q����g�UʅBA,_��fż	�^�}jjj~~~vv���\�$�~�x������ڵk��pI�-�^"��jf^j��BAT��J\���躩2���x���A�@'^]�2�M�ů!�	�Bwԓ�^j�E�^X�78���]AR<7��2<|?�E͂(���2�5����DUQ�&F�627�U*M�1��۷�����hZ�X��[v;r��E.a��FO��0�~H�t��~'	jU��\�钴8\�}i<QNS%�^��(J�����T��҅�Br+�0D�F��o���I��t�DtU��t/hH�f�:�tfUf�Ġ͑%����x\m#v�J;��� 
C8�	���.Yj���}I�cJ8di�,pV�v[k�H�I��ޗ��"��4� I�6&ق�1����.N#���d����k;��>n灎֋��vj��t��D���`�HP��-+U'?��/\{�q h��'���{�;�Ʌ�t̵6ZZ�!�1'LBr�l�ux��cX�j�����O ��Eq���ܽ��ǉQ���s��e�k1)�
�D�5=Q��#ǈC�mj��sѲ��rMK��mo�̿^������Oz��k���?x�1Ǒ��$C���7�t���X��r����Y��K��Q�5��a%;=�,G�)�s$�B�S���m�G��v�9r�$��n��|��SqTT�J��"{�unZ��S2rD�cd$΁Zvݱ���ޟ�t��=��H��z�d@.s���K�[*���^�Dɗ��lI�����(;sFQ�~:$�D,ל|��c6>��7��;����U�o=TPx���_u����F��WΎ巽�<���~<uy����[Y���}�k�}�SW�~b� V�?t��#�Rh��l�op�|"�.I���b(M��͂,ŭf�A�@!K�4`k�%���$iɌ����d�rEmI���@�0���z΍��`��M�T*%>0�,E�sw�ȰAC0�������j'e�mR�Sd��3�+3���M���T���8��f��#\�/$�"�Q�������I����N���cZ������	]�{z���������5�1�Z��P
T�%a@_��M/�Z^`��X�M�֝[�%K�̈b6�ئ�0�O,��7�\fC.��*D���0r=v��a��q�Ty!�	*���:�
�:B֤�@�L��[5�)7�Eŕ�QH_�ȪD����]�����+��<�d���z�IɣYo$\FӞ�
Y�T�\����`�	t~���Fӻ~��g�5���#˓��Z�LK���|f����{������kpp[���j/����WWu�cd�U�l�JR,��W��r�I���cM=���o�G��(�:�$k�fʡ211A��Lֈ�!�'@>4��0,��M4�N� -rHp�F�H�&�As~>���z~���^eu}~+�[ /�~�M��$G�$$���;��o��f3��'�(�U�,-��G�]Y�|vZY�d�7�OR�GvI�gZS$u#T��7��ɬ8t���܇�ua~6k���ds�p433?���]Z/��.�z�*����AS���3x�^2;0�Ԗf���Y�$�x�}��G'��Q���p���z詇~K�mCA�d�U+�'ͪ:Z��\VS�s�Ry��)�L���"��I�n�|��$�t�7�XV���C6u4:���H�*�j�Q}�9�CBm���fM���fE�����q�7F��|�ɦ��$Gat�|���P���e+�M�M�N\����3���`&�"�J��׊�4C���N���$~�6Zv������{v���>z���r�?\t	i�m�?�Ѓ���}���M�tn�2��,�Q��R�):dͺ�b�D����@�k�|����mT�g�鬬i�oy��9�u�ƽ^�淪�C���C�a��[��3�S������~_S7�k��a��˅�oX^�����~�ɛ6?Q�\+�X��ؽw�^��y����!!g�J���E|��Çg N�G(��Xr�+4n�����;Z�ϗk͹rmպ��b~玽(s*�����$�l�2tkn(��odp���v�o�\�[RV�Ğn����aXo%��K��ٞ7�e]X:0::�!�/Ӧ���Z�-#�P M.���߿|x��ݻg3�Q���az�` ��ݑ�3���ON��[|��
��޺e[~졙�+����x�@���*&�J֍F�o�6t,�����cu9�W��v�n~�;.VMT��ued2�����=���wu��%�q�{������'��$+a\S.JP5Pz�}���VBɓ�9�����?��G����`����;�����F���}����~�����_LR���m%B���<�ꫯ>�ܷچ��aS� Mw �Td�}䡇^y����o�y���f��E�_At@G���0hw�IV�w��'�6
���2�D�s%܉�M�%Y�i[���J��QY�c� ��T�6�`s;jI��b5#Y�n��������VN?�[o���,��$��FA�w�~�1��7����>v�?�w���=tU��y����XfR
4շ��{|�lBR��<o�d��c�ukA���ږ�}�΁��:�Ph5tvġt�=��r�M��l��}�����Go��yP5b���C�I=���~�K����쥾V��ҥ��ͻ������\1ڂj�d���U����,Ձh�̙vn��������'���_v����'0�H���w\r�%R�{����֭[e�����Z�h����X�2Q���f)��$��ƲI�v�|oO�%)�$�"����Q���l���DzD���6�yZ���ׁQmn�Gm��#�/s9���[�-cп7n����oz�+_i�L�G���/��rC6\7�LCbD��i�a�@��Qєi"�#q�q�GF�e���W�����~&#��Ƴ�s�w*�&:�n߶m|����]�4Kx6Ȥ+r#��ر��c6LOO�[�i8�����kך�v �T����7A��������Ē��E�l�v[��,�(���'�/t*��-[�,��X�|9��&�����0�d�*UD��,Z�B�-��y
�;��1�IH����-���Z����D��Ў���:��� qoOcϊ��;�qD��>ZR�+|��L�W��y�C�-�iV��(H�ɟN@Q�N�nU��$���>�C|c�W�{U��,���vC���*�Ѡ{7FG�!����y#c��%�K�ly�n��`�'��p��ȇٳgY�u���V�FϒM���|	>_C��Q����v�*T�e|b 7�S���I!������&m������iUܤ]R���n�tE���>K�a�'�O��ʱ@���줒��6*mZu���HZ�N�]J�i�E&��Z�| �i1�Az:&���#I\��!�*�3�0S7���)�`_�b�6<Do�Mл�(��]�!����F�3�Ff/���˪`G�����bI$o����f� 8����4�����Z���y\X� y��U�VѨ"�\̷�e "��	^�^�p��J@�kG�FOO�4��`��
��Դ<Km���g�����ɐ�;m?����g��[�nr�.�(a�u�X�I�Km�Ps^Y��L�����* �1@a��{���l�۠�
�8�/dFܞ�^o���E����|�,���M~d&��\YN"�̉L+H��ѧg��{�U�}�"rlDZ�|����3U�l����Ji�OW�b�iU��@��"cut�:q�y�Tj�2g��ǲ�_�����\�@V����gF���h�4'�0����KI2��Ǫ�0~:C8/���򓓓	�{� ����l�-�Ů)eaʋ�Lm\�g�Ve�g��B�t�6�("W!�8
�<���~�k��+ل�0������/��:7����݉�8���![H���`hK���=�~���"QN}�kV�7�t�����&z����w�i��\�A�F�}Z'��,�g�ίs�9g��]i:8����t@BH�\ �����:�&�0!Zb��m�?1՝%q�w��n�����-e����q<t�G�Y$tD�ӻ�Y�_J���	�.�^���/�&%�]�:�#E5z������w�+����4���ӟf����u��4�ܮ�E^�����̿]�[�d]Փ���f酟��'Dm�P $�1���DXGJ��>������>���fݦ]�A�/����%_���:�[��>��.ʈ���,�;���9��Ѧ��p�,]lKG$	e�t�>��G\�z� ��
�݊��Z8xȍ�D��`���-������Ձ��|� 8>��t�j?��� ��Bݚ�y�X:i'��Oӣ����9"[Zb��-�fg2%�e��ƒc��qt7����/}�?�=p�]�2'���`�v�n�����ɰE��������N��dK�	��XtӢ�o��#ʭ���W;�z�3$Gj��"Qe5W�߲u;�#�\)�bCW�QfY4hZS�.Uز])�`��|Ws�AbД'��b��Dv�^ˢ뗱�?pU�^��-?��ĥђ�#+Z&�b��j������kW�A8���܊=���aO��h����&�E�#����d:�.���B��,[��l���>T��{h<��3d����,��B�M]�r�th�_��jèP�9�&|2��l@��ؾ�I�H6Ѿ3�6�*0f�γ�1Q�s�S�a�Ϙ��|x�6E!��T��X4ႉ4�
���
�J�X�b3V�(�1��ruo�^�4F���l�2�`����]���*0�B�*�ʌ]O=ߘ+�kZa�K��YXuSc{��<BӉ�����R����b�꣏<��Q�sU���3zz�=�ѳ7;��/��� 3��$CkE���L���	|�Mh��F?��tO1t�P��A�[Urj�j�<h�J๞[j�҄������Kr�0M-@�Œ3�h����M����VM	�rb�r��dLُ$<fU�̄���$-����YKKUL܍
�d���$@���8�L��d4��m�P]�+ka����'�i~��i�uC�P,T*%��a[o"�B��n)Q!cŖCpm��S�ɳ���zr-)�3�F"��� ��(���f�Z߷x�.��-���Q�D?���f=�r�Ⱥ5t���%K�̆��#MO�y�T&��f�v-�yC��uT�M#1g�	o����������:B�༨4�^/R� &�<�O���\���L�L��<��&R�f'����	�!Z0����(�2�TW ���n�l�F�%wӦ�%k�И�m�F�|�����:�*4�_�\��p%�Ĵ8vF�ݾc�s���\�l�خ�g�{n�ƍ�\����:�wbll�2_�Z���0�(�ZL[r}��L�%n�r��m{��,6i�[^�tiLj;��7핋��Z��@V�����e+s��ˮ�k0����Q+(h�vO��n�d��$q�U"c5MM�[�K'��l��\�t�f�ݷ,�,��$�����]��ؗ��1�V.fw�[����P�P�n�6�Q���9�d�F]��r�N��cՔ��^:8ܷwf��Zb�^F��=;1^�!�.kg�(VLY�Z�Л�λ1y]��D�l�Qj���>�z�6>U��׭��� N-��ŮX���%Nd�����_�i�o��3~����tAS�9zԑG�.=��y�5nx�j�0���;o~�2�{T��B��?���~�������|��8�h<3q�X�-4'��z�G}�{.���o8�����L�~��O_�k>u�g׬>��7�ŉ4�[�Ro{녿��=��UdK��l���t8��k�|�C�����a��%�v8�|Иl�n��w�(�\�����v��0-"�"�O�E�T��]�E9��w���R����s�>ᨣ��������y�y�4!&}Ҵ~���)��MM6e���u���z��������:��[o�`��R���׮������־�-o	9K�ԣ�?��k���{�y��'�z��N���ǵ׾�s�8�Ҋ�FKǺ�E2b���﯋�_��}��.AN:�9�sމ�/:���� |�e�k�H����wr�	A��s�/
�ӀA�,8��
�p���r%Y�"8G�'�(Q'J�J$����Z��m�hc�0y���#.�1/�.�jh~La>���	���$^,�OE����U��D�9Z��g�(���!~���wdg�񾱡T�E�n���lw�f�ѠZ�Jx#��R��_"�쀎�5��¬`{�`=�����i�����I�N�8�\a�hd�1����[-_,�%���\��-D���Sj�W�g�̐��`�E�D1_\�hQ�2{zz����o���;~�&�,����H��������u�|�ɱ���scS'����)U'��`�~��ٌ&���R�a"/ag��_��ח���?�M����^��B�Z�V,I�6�ڴ��;���g���&�*ɰ"iYĝ���U��V�r>*�ʎ�>%�H���0O��>� uit*��&��n])f�{�:1i���#p�{����gl|6}��,�J�[���{
���?�3��,a>�ئ�-m���萟�^��w���D�X ��*#MF����ǀ�=<0��w��&>�iM�=�1�H�� \��"�X6z������3]��N�;�ȋ� ����u�ֹ>2oY���h�u9(��1Q�UwϞ=�-7dr<�9J����'DF�a��@{�-�A��ZA|����j��w��1�pi$C��� �k�!1'�)8��GcW���'''�{�h@��e�:��޴��rCZ:l�}C��m�1d�dI���Y6C@�g"d9b�A[��Og�C�]�JHNҪ<���Ҷm��s��47z倞
�G2���G����$���ŋi'�%U���B�m�
���p�xn�-����gggQ�A*d�W�|u���&Dc�¨�)JW�t$Vl�Z2ZI�8�ld8mӡ������Q4Q�������?�c�Eg��u�����ݥ2�Eb���V�\Y/M�\�Y��R�YL�68�w�^�iO=��������c��r&����D�L/رe��ݻG�bs��B�y���s�=G�w�֭��W]uU.� ,���$-��=�,K[7�
"m9��m��
�͛7?���BEH�p��{D~)� ��"M/��d�ۗ�o���S�Or�b�
�"��/���/#$�R��2?G2C�D��b�b�|�!���{�M��Z���֓-�����Ν㫖/9�S�<�L���]{�g�&*�Jƒ����+��2�L�F|�h(6KE
�H�C��Ȉ;3S�����-[�����f��(�L����z�-��$�@�,�����=4�믿���] �����˗�1q�Yg�w�=��'�|\��@'��Q�"0I7�iӦ����6R��kD�(�5e�t�����wш����'�x\4Dξͧ>��K/�t�qG^v�eo<����~u�g�Q��������h�,���@d�b�F�QHc��W�v�������ml�}<����Z	:�=�,VJنCIEi_���赝̘��T����g_dP����_RJ��i������Q�!�P�$�O<���{���/��:8t/�G�z�]wm��zv3�6[MUv��ҵ��ۏnܸ���~7I��H/=N{��u�7y䑀��P�r��'�+_y��}�m�{�+7�������zɫ�JIm������K����"K��ؑ s�%�GD�U7p-���Md[�jg��K�&"v�x�������%���EX�!3����nF4��4,B��ĽO�A,�|�6�H:���& ���&�k�&+JR#���0m�����%�>�v�b��s��[]VLR� 7�.�MOBI�Mz_�������	�E��j�󣍉�)G2	�S�t�dW ̀U+����b���d����bD�U%���:�i�Y����2ˈ�ɈL1ͤ3T/|�pr���CV��)��O�(<^�f�E��
2R�f_�ρ�v�8��E��M�c$�^�Fr���<�æ׺����u� QP48�S��ٹ�a���d���I��(��sE��Y5�{ݲ�h�1�n�وQ%�ߺ'?@G~'d��at�}�U[�I'�b�R���۝�8A7��?�V~@Ƅ�M���y�
��':��Z֤eId0Ţ�J���]<<b;Y��f�'p�0���vl9�%"%�E��+o
8w3q�m��.
�:A�"fVe��@"��T6�DvK�F��Z ������r)��z���Ԣ��I�P��91�}����:c+�A��qI7�zT�a�zl�ʠ�j�ZuYeU�/�.�Qݎ�7{I�5#$�Β�-���|:#/�i��ffI����[tFŌg��R�r���)ph��҈fd�:��C#�=A�%B+;4�~�7q��܈��%&���Y�/�=�m��V$���W��.��B�\���jQh�d����Hj�"ي�/�Y��ޔ�+Ũ���J�'S+�JT޳�9[�{�����d��"��5�b����[z;.7�W�x���Iamnzzצ-��63�ش
����v[��Co6��E�Fo�����L�:z��E���Aí ǫ�ur&ݍ�K�#՝��g��w��=$�QD6��8��������$��ĕ%� `��Ҭ�����c{{a�哧7�-�����hh��4�%5������~+����x�V�Pь��x�(�MMXNPt��X	v��H���� �R�,�ׁ��V���
����W��rKj�l�|��|t��+�TXM|�:SoƁ�Dz.S��{=��W����ǚ���ѮX����o���]�v)S�,�T�*��iEW�$��LO	�����G!'j�@�COn~�g�;���U����4#C{�v�Q�d�~��`ƙ���w��1Vz��V�1Wk�������e�W��g�r��~�r�g&��^�v5}Tsvnnl�䇴�tU� ��m+��S�,g�*^87ET.�Ӿh:eMGH�"m<�{���ޑ�~:Mv��^�~�k_�Ν;I�m�FwD����׽�կ�'���ƞ�m۟����oh�`T�.��@{���۽�c���>���￿XԶmsMKY:4�l�i~z�傷��C��z� t�H�Y=c,X�x颾���V3�tjl~�+��>��+'�y2�TùJ��Śʹ��˥6?����d�s4B�-Z����mϏ�]~ŕo��Ð�dI�Ǒ$$�f6�������Q�nQ���=-+V��J�mR6	=�����5�<�ۘ� 2�h
t�%�&,I�7�w�-;�v��'�����zR���굂�X���e��r����br�����A��ɿ����>����}����eQ(�\ϲL)n���̔0z��/8���������������Yh:���]c�Wc(���N6�q�)�����$6a
��A���?;��*S�,|��6�~�|Ϧ�+N�pʃw�fbvj��!pp%������Iq���v�׿a&aV3b?��;w��3��W_u�ɧ�@W'��Ր��Z���������_�ʿ��Wv6
�(Bb��i�4U�h�/��/�0��;4����[Bǻ��/ņ�S*��`/�'��o?���>؁���׊E��H�w8|;�r`oJ��,d�:o��J�~mr<�5�0�4����~��dƥ����iL���"�*`�D�Yd�E��E�u�H��B�}��O���'������"#g����u,Ce�cٷM�ΈJ�f*���F�f8 T��PP�R��8�� �P�kZ��N����gÑ�D|y,��? ���r��0G�T�FfC�����D9�O�2��AA�)�*���� ��S�a���w��ڌ�)��@O������h׮]��Bn�}���<[*����###���4~_D&L?0��ٖ4�UtR��!-�ȸ7�[!eM0x<���#���?^�tٲeF6'�&=������	-�X�>�E^c��pzjb˖-��X0[����N��1Qv��0��P;�'v�*��V�u"�e(���$+��WL�>| l��pm;���:��9����>Y����W����1Ū��J�l��
.��V`ʵ2*�*MN�P�sY`N6!]Y�V�3�;��O��m�N޳�3�b�NMMF��i�J�QR�|Ǐy�~�<ݒA^�-�aU,}ff�oy�W2=6ق�h;��<�q��P!O���X�%�?���� k�^I�α�quMH�z��kc&��"����V��x��^�5�+Q�%���;4?��H�H5�v��ɽ���Ԕ]��f�ď�&_!�GqDX-�����$�/��F�3B7\�I[�Bo�5��7�2��$��e�)�Q1��R� � �!3(?0@�j��5��S3�4��!aػw�����w��(DQ�i���6y���q�z �N�պX �PZ�ia�K�YS� �URSX����$Fb`�Cl�}-D�@�F����5G�y��?-����S4�fۏ��T&I;��h��;�<�D	�G=CCh'��4u?��-���5��LQEG���Br888Hkz�]w�r�-��y�~�������3������+�����R3����I����	���hࡪ~��@~8�п��ġF#'u�m�5���M����.
8BA�/b7ܝ(�EO�Z!׶�<$͓i$��i��L��#7�x�%K����yGI��hY�m�l{�}��5�7o޾};`يA�Y{|�dH�*M��f�<�W��UGy$}�۬!ab�1,�W��=F~ݽ��KȮ�D�$=��h2wn�h��K�c�֭4E_�J�?�}� 6���}u��EMrH��!E��7���\�t[�u���SN�����@�qa$<mY�1��2a#��E�._�8��؞�]I�}��^Gviq2rN���̟	���O�����9Ȏ�;�@,#ɀO��D5��<�P���'h���/��G?BSh6�$]�]��-n�h�
#�������t>�2PL�8� _̕USJ!IhQMyaSS��Q���x����s����~����}�� KAmHSt�g��&�$~�'l˦ǁ�}�
��IZc�6l���?�䓶a�#d<�\r	��z��<i\����d{)E���\"�!_p�����ԁ߲�Tw������^v���%ӑL� ��N��$�=Jb:B�^�2�����:d�(@=��ͭ���atW%b�,��w���H�M	���@����I���������p��EH;P�O:�ց��d�2�qN;��:�I2�M�.�h�S
�cd�L�� �s�EX�&(�WW�B>G:�Eꀼ:B�6���4���8�U(ԛ�Dݡ�V2VF�l0��빚j�^Sްz���&�
%nrr#���r�)���P�G���AI4�ȷ�7�u'�p��85�7��B�:�f��ހJbт���	�y ���x���-V����"��D!���H6��8'�$qt!���|�"��`gI%��Gw��h�]��ܤ9;338<ԓ/��Gߠ���̜�,��<��&��mR��WӔ��M�A����r�έVݛ���h�tUX2���V_�,?;S�6a�E� X*m�v��&�Q"���H���0ݺ�dL�V=/�?{�0+=	��@tW!N(¦�j��	e^I37ܔ�I��R��|MpAHQ"7�u�2�\�Y�ކ�ŨA�~�4@�����[Gѓ�� H���Hh輲��5e�S��Ua&�e���Ld�� `e[VA�3iUg3�����*A�� �d�h9�9�b�M��f��3W��d �����^S��#��qՂ)e傓��}��x�A�9mTK���~���e0q~7ɉe5�7L\O,�ɚ����<�Z"sn]�ZCN1o[{t���J?�]�vT�ؒ����8���/�m-U�f�-K�Za�Ƥ 0�n��8��Dr(%�nja\K"��:J/��}78P���jJ�� G�<��L����9���Z�d䚪�j�t;:�W�&$��j�r����C����i-5e\�U#lyQɔC�TٛMhH��Z�Ƥ��ʈmG�?hZ�~� ����=�S����Tk�!G윘������e�Ug�39��%�vv�L�{�c�`�cr�K��J��t�1Ja���q���&�̱����(�}M�� Nxrw �l��"��TmQ�e�4�Uk�EB��V��ڛ�e���gq�r�ҪJIK�h��&�>���o�_�d7������-�Y\L�d3�+�4��I����«�z�Ĵ���,3�ɟ-ϗ�HI��L6���0n��ae�9�B0t�4��
j�LpQ�������l	�V�3��+�b��	3z�d"�%�jJ�'E)�P{�8��\|�a� ц���Ť�v�[�ny�[�~���e+�����oN>���?!PGN��X�����ݻ�ǝ���C!G+Hx~+�#2��S*�t�ťf}l|�[�[�aK����Z�"x2>hM����9F��{I��0	�2���~�t����s�30	rAdű�jS[�?!�+ٮU�B!I6�窐WQ��0�Z�b�yP�s�e�-�MO?E�30�Y�f��QF/��_S�.
��D��� mY:��w2�N畀W{���?�������_��'g;:���V1ؐ�H
�ǟ��l:#��d���|%�B�pPUc6���t�݈��A1̹�0p����B�
��"��?=:g������빾>��L��E)��;o��u���ڋ� *��L!��쀆w��Kn�R��ä����uh��[����/$��.�v�=krm����s��o��s��74~��綏�^}�[�i�C���m�5jd�e+ד���C3[w������ȀC���ޙ�_�['�v��?���������|��+��կ��p�&Y��f�rl��(��fW�q$O�="Z����ϋ;���Wv��#_/;_Kj�Ȋ�Ю�]@B�L��Pi���+�H!�!�2�P���ʄW����Ȟ��'�'�,r�Ҡ�ȱH�;�]D��;�˂���/��:��C�^����*�����.^��,�N���E��RM�d����cvr��N�7{/�m ���b�� 6�C����	ð%�BV�g�ƌ�2\!������#�6mj�0�I:�I�� zVr&���*�m�r�_z�Hjug��^�$����5J��(��1J�!Y}}�BJi0�7o޽k��"�9�r�Y��I8	�ۜ�Ʌ�ڵk�\�C�E�S��M.g�E��u���n4::Z�.��C�rp�w��<)톿�N��@~���c���ۋ��$J�fs��U� p���SRHi�D}��32!@"ԨV�V�Q�B�q|��/�,�G�~��RQ;���k��Jdf:��*�"�6d�I$tM���|�*q\�'_<�Y��tg��ꮇ�����"E̹2���1����c�7@FWR��E� �ϧ����:j�B6MF�pj1�,kzz�X�
�eB#�G�ʒ����a����Һ�}633���gL�qq/��u�E�`o�ܙE��S��&�Z����B/�o�>Y�0I̒���;-D�"����	���YaO��mz^G����d��앙J�����LrE��x�l�S��:���D���z������XB��-����=�SiS���<��#�z`y�j"��������k�"Tậā�����=I��i���D�>�%̌��)8s�.����.ٵ7n����ȁ�oB��+===��x��`˖-�Z�>߶�=0�̓|���XQ�4 ���F���8a8Q^��Q�2m�#���R��dF�$[���}��4���#�}�M�!g������~I���Cs|z��� ����K���#�:$�`���K�Ɇ*/Z�h�����T��$�&d@��4�9C�Չ��0"�������>�&��UC���we���C"D�*b�Wdhr��4�H��,6v�c*_K,YЄ4��O���!�J��֭[��E��;���O~��SN[�z�ڵ��G����'~�A��;�v!ŧfE��I��ܱ,z�����ъ�{���3^�j�E�C�<f�Ν-����xrfv�޽�VAx���
7�``�]G	:Q]�A�/[L_J�}{�5F�Dq��Z�"�7|�Ke
�g�}v���P)��U@���7�x�E�`�q&�y�g�z�͂�ִ�K.���.���!���Ӕ_y商fx�jp"�k�c��".��-Ca�-��V�xAG��G}�ݿ"��z���@'=>4nڧ����������.[�r��g�-1|qԕN-CA����B�Qu�Ձtgh'��b4|u�'�]�����)�;�_�O [Ne �&3�����5���OD;e�?G�׭���ۛ?��h���>��SO=�d�n6Ãd�\d3Yr��.c �� ���[�&��ԧ�����򕯬�P6I[줓N"������������rXVI���䗒?�Sk?�G�2<��/�~o^x�"���B��~
/9����ł�&�h����H�C6�4R��ȵ�K$xuB����T�Ÿx �=�b$`B�4Eǚa�a�p-b� ��أ����x\�f����VH�m���ă9sN\X-"ҁ�aS�@ I0��Tj���->4s�#ji�D�d����D��u�<$:}�q�げ0}�3Fy"8p5�k��O0$��ܢ'���h�����Yd�rT���A��sr�hP�܅�Ls�xN�y"�.��X|(;ԣ��#$�
E���Y�}~��\��OB\���?T�<�`�1"��H��R%,1#��d}��0U��J2��y-/��ba(�+$��6J�=���t�6�P��lo`7��j�Rk0c�fg�<�Y��6tǶff��;����·��=����9���|���L�4_I"��ȭ�����q�&Z}ƚ���t6y�Pն�Bn��YH�r��8��%��@7z���V���Dr�5[���l�ȭ 0",(YQ�i��VY2Ty= e�3�>cX��Q�9�c�^���SIjr�Y������Z�*'�b)e��C��!
�䈡	r�� 4аtZ�b�@D��Ҩ���f�^K��P���5�xn�U�3Cn)��_�QW0tE1K�[m���҂�����Pp/n&_ @��L5P�Q��HS��k�}�P�u����5�f�&^m�����j����b���V��7�J�1�bQ`	چ/3��*�l�$�/��s%{FVcY0?����t�~`a7�Ɓ"�mY�YZ`��<�>��}r��x��G�Y����c&�e�>J�2@�@f�PBQ��:v�6���$ΐ����ĕ�YG��|mZ/s��CW@���}���ϔ�j��Ș{��{�Q`��0H_�t�!;�l�gy�N��2W%��J���	ڊ�A��po�T�55���|蒋}�N@>nBcho4���"�r���+p[v����Dmy�`������ᑑ����fl�;dDN�N�A�C�b�;��``�:��S$�5՘�j�ϳ�NE��!�s:a-� b24^ļd�i�qߋ�`+�#A��J�t�Ak�p,L�I��U���� /�S7 ��8Xa�q�k[,�;Y1�Z�^r��ɽ�a��=�m��O�!�,,[����*uzri&?�{�D}�2��`�ɐ��.��S���r.���Z|���fI��AT+OѶrd��ľ����b�A�&2Wf�Y�q�keFȈ������*���@�X��b���tT؊&��B����*X�����R�;N�1$�lE/��gn�Mf�����+EES��|�R�юX4��v��<��M��F����s9gp��R���p`��-T�Zunt&��Z��q��"
��~]7� ��w��m`o�p��4qS�$Qrh�l�z<#/g�V��b,g[��m��!�Em���Ņ�`�w�����&`�U����p����z�z�D�l�  �"�u�Qj&0B���&��hP��L@EE�Af��硺�k>�����[眮F@M��s�=Oq��}�^{��{��l���ԩ{M	<�2K�@������?�")�z��;３C~f�����X08$huH�\����IN�_huB?TM���ڵǑ��X$9��n3�R8$�6�O8�=6c�\�l�&y�a�,�֮]��m:��7�5�h�l�(Z�1Z����b~�k_���[��c$�K'q��g�bY���Ԝ)2I9�vhU�z�bŬ�&-�oi��T.����!'Vi���Gr"w�_�s�V;_e\�-m��q�ڠܹ��e79��*D���
g�9�~�u�}��m�����y�u7�v��g����N0eGi�$�c,]���)��j������00	<i�@�jǮ]OO43k$L�dɲ��bջ�o����$��+�f��O^��iبCA3Y,��őP��t���\y�|Ҭ������U�΍�?�u_p�����>Y§���	x���q�wW!��(oQS�"W�z/��#���o��F�"(�3aD'��M'�F��b'���L�/Lǐ�'"L���q��:%�r�u�RdT^:iҧ��[�Mf��G�;��9405��)v�D;g��"�h�7<�ә8k��� �HX�I"?�X�[@B
�vh!��M���(Q��t�0���$��a<������F$C(�+����(r��N�$H@&�r@�(�ݫG�O�Z/E#�R`Vy��E[F0JJ=�Ǘ��ϺrZ�+NF��|NU��W�<d���t"�H+�����$9� ��r9�:�K� ��*�f��P(LW+�ɘ����Hjڝ9����b���g),yZ��'�>�|2��Ѻ���i�gd1��,�\��u����~d��Omg�Z�1��ij�|�F�ґc�b[�z5��s;�6Y8���>� �]�^[�jբ��9�ʣ��)C�p!2n�}���?t����:'}H��\��G�>�`���&t��	�h���u�Q���	�]qu nX�-bUr.9��9h&�QIr���V/_��1=�t�&s|�Ns�^���눹�܏�si_Xc`�)a�;Q��Sæ��Es��0�S����(Z���|��H��.M2��~�K؆j-�v[�t���� %/�K��`:�D�mN�w�ZJ�
��@M�Ι�<�D������l8��n1������7��+%RȦT&Ba??�zN�ͩ�)���Ĥ����{��`���cy�³ߘ�zdd$u �jx\�n��������w�dtf����خ�4�m۶ѭ]��w��j�����\���319FvgX� ��b�7G��t�M�F�D�U�fR�lS�˲�a�3i�e��g���ƍ/��-_s�={�b+=52��	�}}huc�9 >�E�*��-[F3�`���:1"#��Y��k&��b��L»�Y�HY�p)x�y�����s������=�;����k�� �����@��)������W��K��Ӄ`@j4�ZkE!�
(�ZTfr# �b۝n4�U��>ej�t,� Z`�_Z�W�M�'�u��	��6v�i@��'��ȇ�Dx�V��#�;�m��0 �LRt���T��L���WQ;�9$��ڵZ�v4�rB�T4irh� �Ԯ�y0�UԹ)�ou��F%J'\ �?��ʓ���l�S!�\����De]�:�tIz
I���:�]�[�qN�弖q~�]�Ӛ�ߖ9�&�����Gڻw��ǯoUߌ����z�1�n��O>yڙ/��|�>A���k�>��s�I{�RdB�W�Q�8��&�-�b�z衇�x��N9�D8�p��qlV�D��}���,X�U3$��"�=Z�|�\�r 7����������5k�d��eމ��a�h���V�Vb<��]Kg[Qo���9�����2���i�E��J>iKt<1iku|]!��vq�����KSP;V�h#yȪi�ٺkZ)~�	�1��ƍs��O��S^|I0Z����g�̐V�\��\��?�䓧���.: ���B?M��ѳF9���j�u\YFخ��o��}�C�q���vMuWΤòvY���ޘp���^p��DIT��U�v���x�Jϸdذ�L����\@�)>`͑ӧ/eS�c��^�.[���"�4@�4���+͐���5D�A�g�BR5ߋ�C�	N�2�Z����������Î�)������v�`|B�a/����B�")-3yi�X�^�D�\�b&�rrsrK��"+���b��dj2f��q�f�8�؍�1�SZJ�<�� �t�B�\�\/��O�j�q��8�*�V��Àv���q��G2�d�\��"�6H4�~�C��ɾ��ق��&�Bk&�L��@U�㦟-�Ka�D�xx�H�%�#�L��9t�l�$��5���j[@�^w<��D�L�[p��]�Ȕ���(��N��o~��� }s�Z#����l}��4�,�YpT�a!��I��XSg�rb�4�0��UE8��BA� Lb���/ۺ�u�K��P�{�f���版l��4��C��,o�mT�B����N�&Y�r)��XB�4�T���@;D��fF����3�<���O��^ܵ�k�.���*e��>��/~���i��`�����?�q��%�_��j���'�(�����ҥK�Y=����d_��h�q_��ilf�p�E-!_k��[o��J�����g`i,��9�-�����ZΡ�ӳ|�1�����U�Q�Z�Ͼuu�n��Am��E_{>�	݋�F��Kf��+>슔����w-{��^7|�)V�@O�N�������ک]O�B��h<-go~�ٽ�}ꩧ�3��i5�Y_�'�h�c3�LnTN�O�b�d;�#�}W���bS�^B�6��b�	�X�"x��$�i��C7��t�f1�������g0Əkj���E�g��W3�Y"D������O���J�l ��M�aG�����U�\��Z�4�@�^�E�h�T��|����`ת8�M�MOM�&�������U�o��܁�	Ӷzz��m:]];��w�#a�y7��$��%������~�dD�@ŋ�{zȎ�~��prB,NȰ��T#e�]画�Q$^\��tII����x�+��2;~�{p0�U�>x?�݃�ټ�����Z84T�:H�r%�8p`zt�Δ�ݻN;�4���^�K�C۶��wp��p�@B���dJj��D��l-^�����_�i�r��/^�Q�8�h:y�+W��\7��Ue���A�Nko�0p�4iܒo��ɞ���%�m���|~݋Ԙf��2)��t^�Z;	G�z��p��ƽi�D���0�TSv��&Cv#h�H1cF��U=��t�LE�hʸR���s��t�����C��+,T�Q��k�ZR�WY���O�F!I
�A�p@P'u@Fd��3�E�] �)B�(��*2��^�M�Ԣ� �4]�=�ܐ2��ע�����=
���G���ћ���)3�Hh��EE�v�ƱaX&3W��P=U��QT,I��$IĹ�[,GJ�t���	�2i�QVSu{�0�X�)U��)
�T���53��� �d$n�̅=�42U�-s��D��LK3�9zM��?������'��d��v4)XY�Bˌ�j��F5(朴��J���%dl�^��-�Zi�D�ut�&��Y�k_s��~����z��N&S���I��k �"u�f��_�Y���?�|I�B�ͺ����<�lf�M�d2���Fÿ��O��_�;�.�L1�w��������Hmr������w��ERy�0'��k����ޱ֔6GB+���@���ڵJ�:�l�����kv,7�.��7T��9��޵�^Q��!M!����Ԉk�^r�i?�����G~��-_�����#M�Fa�4��T=3ճ_�ҟ���;r���V��`�J�N�)��YR���_ϔ����nX{�	�R鶟��aA���Xd'�x�Yg��������rX��Լ���#��2�� ����\��Ä�^p���vK���H�iY^��6�s̞Eyb[��Qx��<�HB���c�`�[��8�%]BbS��"��26h�n��$�`�b�k�����U'�!7���l�<��jI��仒6I���t
�;t'J�2����	\����	d,�L�#�;	���`Y����:."(vQp��{̚0|?ж��KM�`����e2�@9��-�Z!�硇i(�
2�
E%qi�`2�]�����)O�Oƽ��/'�W�3q�<4%��������LS���\�lr1Me�ﳽR�L����Q����$+0�����2��]˖-��gƧaa83��(�������Y��F���G��(t��]��;v�M�d� %!8�ܩ��X�x�nY2�!ý�<�[�Wi#nSKW\"a��$iAo)�[X�kL�$��q�j�{�!_�K�ޮ_�vݺu��}���LNЭ��$Ct[�nuq���/[��f���?���NV�[�,�u�N>��''6n���'��s���p��U�Vх�:	������Ek֬��@~cӦM[�l9�c��ٓ�=$ͨ!׶|j�%��|���U�2�m�V��Мӑ�PLE!=�E��Yt��m\C5�2m��aPZ�d�Э>��5��������X��B��ݷ`�J{�8���zs92ܧ����d���T�bNS�	]%�-԰�n1���BC.��"Bjq�Vt!�@T;�)t�CRE!S�p�G�?݅� ����iD�8�*�W�(���
��2z����.X�c`��X�_���9��p겈��&I��[CA5ݾ�^Og{t�Ug{{���pO#ݢ�D�H��n}�I���O?�t����u�L~��B��S���~���"M^�rc��X9��B���+�N>===QF[r�X�}�|�r |���io��{h�,ذaÒ�{�0Jio߾�.4D��ԏ�^'��1�d(�;�TZ��AZ���i�-\���1��S�i��V�O=U�v��;w�l�j@����J�5���"��Ɖe����X����H��lNk4�B���:vO��H��h��?��	���� f	jVU�JgG�W!�$��8�;92u��۱�q��O���-�X!	��QK�����T2)��3(�����g�B97�vr��S�A�};zkU�_�W��pJ@Of��v�9� L��c��u�}erH]��m�dby�����X_rxZ:�f6�ٶ�ۉG�K���E]��O����,��7���R�8HIٶ�Y*��G�lV��#�1�5�Ne�c���Q\���Z��d����{��>z٥����_���}��E7D�� �LfD�R��Khw��]�B#n�$�%�(\�{X�#�'�f�iT��	|	Ԕ��"� LKi�K�=a�l�M�v�4dKj[�j�����w%�b�P"7vR��`Y�$w�DÖCU�-[�\���igev��V=�-֌2�l3����~��Iv}�;����}��vp�	��X��������/��O|�s�9~ņ8Hɾ���|�LZc��=��Gh _|����У�뮻���C:��B�����r���_�|܂e��$eUW6��9;�����w�j��|�4�5]��6g�L͈aOQQx&CV	j�#mK�sa!腄iHk+�PQ���		��c�$_+eN����Ч��j��$�C�[{R���$;xڲ}9���.I���zeRLtboJ*�N�Cg*d|E��R�;�0���Ud2�������������ݤk�	�pA�1�T���P-��p��|�
�KD,�0��@��ii�v>!�z%+�b ٧4hD�W8\�BIG���zB��D��aT`�F�H��W���de��	-��,0H�eq�Ե8�Q$iP�H�=�r�c�?��z��C�#%��di��4��<n���G���J.ˑ9�h<�ؖ`�	�ū^D~�l%��c�c�5i������șJ�W~�jZt�)/}}>8�`�}WwMC˒�Ef��e^�h�<�twl<��B���ts��Bw-��J9|�&:��A�(&5�SZ���U��=:mC��qDg(�L�L��
��J�sǶboa�`� �� ��� [C�֕�2=��,)�(�9@U޴����o_{������������{����䝿��,���f�=7�~{�����_�߯uu-^w�h�z�c�����П�����V������%�-*->�a�,����C�#��k��;KOu��f�
tfš]	��jÃ��M[��A����$��U�yzRN��,90y(�%��Xm&Z>�Gn������bs��ի�A��Y����'�>V���,7�׍�/4u�OO�\ob�RKj���Bh#�/"����=v��z0p�[�=�y�O�Y�*���]��[<3��� �C.��0�HH ��)�KT}�e�c1�"U-3iM��;���:l_�Y�'�,�J�? �Y<\}
QЌC��0S�Ůf"�,�$ʡ ��"�UU䣬) ���L1�|�M��LWg���LCA+$���$G����Z�D�)xm�SS�O=�x��C�k�T�� 84&���^m�M0�pAoo�Z4*����ܵa�K�V��FdDX&=8:��&����ѩ@k7���.��HrA8a� ��ʻ)�=��󌮮�)t�T"`�w�ߨ��ڽ�ܲ�:{�g�3eO?��S����Kґe�o����ms���W��75�6j��(�䥍h7��`�(KȠ��d�>�w���u=]�.���@�+��i�ke�ֶ�;22��rwTff���4�&CϠm.��v7J�Q�%�	�K�o�����"���-|Z�3v�ÑkOmw�t����XE]�`DS����lL4�%�g�
dWf1M�"��ݔ�7l{�㓸�@/�Di�P�e�f<I_ D��1XijY$b�����)��x�[1���G�'CRl��$��
y �j�Mq��ؼ}Y�Gֿbء�Y�D�4�fI߱	0Ҽmd���R�a�\C���Z�KJ:V�Ԥ��cn#�`B�nwTK�`��Q2�|�C�������-n��e�^M#c��оIJ{�T����L�Ȱs��#xd�$�2��7�ܸ�%�ϻ���}�o��~]s5�������X>55���L'A�e�1V-��C� ��^�qIN�:�qDd�dߐ{�@�	�F��������鴓�-��âUB��?��o?��O�jt�5���(E��50V7<�w:�fR�iG��;�~�E]�`"W�hi��+���⋯��o�������㔀�L�,��fh(x4���n�"���<hB!{��Y/�V�̓q� R��@�4ؤO.Co�ԧ�n�=�����}c2Ю�0z`d_F�1��J��CZ�^Bޯq�6vۅ�|蒉у/�tr���jh!�	AgIk@д^{��n~�+O9��?:�7�t-�d���5+�^z���_�B��kH��d��[��;n��I��_㍯z�+T�u��v���w_��.R43��yA���r�NL�;_��ˮ�S�����.g{��Z2�8�4Q���R��hHX����	\��q4��,��]]ňu	9X��ݪ����q����Հ�F���FQ��|2�:��V	wʯ�+���s �:�?ц�[+m���P���)�妕��r$]�lin6�Z���;Q�H&/ʮ V��{��ܴf1�K�3
�Z(�GO�F(��aRW��y��н[v.��
�2�(5B�Jt�9L�qB�S���?5|e�uT*�_
dM�ǭ[4P�|�RYf������C��=�H�$pWh
�0�.]���3k�s�()w��Y���Fr@AF�n�k-�ȍ�R}ӦMK�>�>߷�)Ҿ�Z��'] {IV>�[���O�Y�rٲe����ٳG�o�iΫ�*=2ݎ=����4y,3�u?:��\��{��#�c�����;x����8](��/�J��CJmZ K�.=j�y&;�����hr�{��]rɊZ8@�5]��Mڽ�����q5��P���]��7����F%��N=���v�^z#���b�ƍ��D�'s�6�lf���2����T*������?44!�����_��4ɽ�ދ~����u�I'ɔ��%�J�<:��=!*T]fn��ҷ �;x��^/�>`�*�QL~o>��
 Nؽ{7}ҵ��$���R�Ni1�ـ�k��i�S�5��r�>�}��E�n:t(��1���y�
��e���h[�r���L���7�$Y���$��;R��Z��&��d�Vϸ�F�O� Q�Y2N�e����+ǯ��Ã�g�a�E�@w����4\�!�Y�a<_@�WGVӟ)#7�X�$� #��\�Oy@���u�Z�`�%A��t������6�{�F���C�䒦3w�q�W�>��he�������E�-�����3t�0lA�p1�"�
�����Nz�Wu��J�A�<�,+v�2T:�ۑ�M�	69'r�,���'7�Zݻ}'"Ц�s�N��b�gHC�H���~8��
i�l�oX<��h.�ch�ә{
0�����ZX�\��]yo5İ���)��d��l����aY�.Z�]ܑ��i�I��$�ٖ�"�9�xfq��6���N��MF�66��%'�v"	1tf�<dG���dB�/j�ao�Hđ9ƹ�F�������� iqo�F]��v��Ӑ�rmP֫5�A1Uy�Zj!�5$�Pkb�خè�d���֒�nk�r�.]��|�i��e�r��ᘌ�:R��6��Z2��Hja9�J��{D�;�����	����t���x�VZ&de�.��/�ܸq�֭[,�U�,��o>y�_��_4��ɐ���CJs{�$6аh����&P���I00��q`S�p�	��~�����OJ�:�n��X�%��~��ɐ���aBƽ
iו�k����mTb���=���l��hg�p� ���s/r�e�v�4���a�V!� $ʑڪ�,��V|i�e�4���܇�f�U��a�ĵZ��b.v�����fQƦ�5p�v��#a~�����=�u�֑�m�s���D��7�n�x�?x�K^���H��4��A��'c��K/;��si���'���.z�'��+�r���Z�K'M�a�X�v�G?��z=�[�_rȥ���?�����kI�v�Ӻ���(���n��648��u�]w�9�bM.�R��`0�]�<EB3�;���7��?"�Fv�U���g,����g?��o��og�}���r���͙YP��2=S����M�����S�)���/�b�5I�$�B��@r!v���d.K~"3�� �����:?�),��$G���<�-�	��_��ɸ�	�2�i��T5�<��+���w9��
��	��w�k. �$@Z$�������������k����jR�=��ӽ��#ra�5��ˏ���t���RD���A*�?����fRA&��׼����743�Ţ`hA��*�IӯX�p�1L�f,_�����kJ�'��p��C�����D�iZ�z�K�����'Ъ��݃�[��fMh�<0�E�E[��zt$��h�0�7�f�E��n��=Yi�0�^K��ђ�rn�TL�T���oh���5ݢ{����޾m��Af�����/_��yg������TU��j�\��:�@ʐ4� �r�F~����POFQQI{��+���ݶD�4���j��R�rCå GGw˶V�Y{�@%�����h�Pޙ9��s�qZ~��ڹ��!ñc���,��0G���qݛ=8�tw�}O&�KZF�BDs��؁bU�FB:Nw�Y,�'��LOҺ]�pa���L�*���Mᘮ/+�:WE{���&>4�w��b#L'��n��$�)�Dv�Gyw�@LE+XN�GI��O7G��g�졳��z;�J��1�b	���TXIj��q0�V�����t�Vr@��i�H5�3�������v�v_m�2�����6�"��$nHЄ(@R��Q�@g�M4�d�H]K)h����"��2��h&�" *R�#HAF�ࣅ����h7��6�� �+�m.�O����OU=����	�4��P
hM���$V"�&�,�74��YB��r���?�L��*�o��4�o��={tzVPӤQ�N�\�͛V�Z���/�ii5K���R�eg�Fqp���:��pCM��An������&�ڱcǼ���=jM�46=5�����ڼ��]3�>TEA�(j��r�/Q��i��3���jj��48u5g�f������]����[��f�������t�P�vY�ϖs��9R������hju젾r�4�ȧg�Z���Ę���)Ǫ��\���q��H����7�j���JW��5�Z����͐�K摩�]ŠҨ��@�	��l5�eKMKR��X(��kZz��1j;h6�QH��Ix�ĹU4(�j��m�"���K`�ߥ��O#��{��V���?�uB3"���3���m<pt�8Ӳ�S�^�
ȩh�韤eb�٠8}E\E)E�r�0�cɑ!/Jښ�tۀ��&�q�}�����8Iq�e)i�7[���摄)�t�٥�$��$�#d�R�X�rC1lR�����:�2Y��Q�� Ƚe(�Ra�o�	��W>|ҒMTچM�-R�eE)Q�U�#�:X�j!�$y ��Z>&�+��[�X�l<N���Y��j�P,�r�	�<����g�q&�$!�4?�?q�e�^zi4�VVT"A:��r�L��@d*9�h^C��~XF1���M��Ti�5@I��tgә/ϒ��~�C_��/� D��^u��7�E���6�W�i01u0ِ[����@)�*���6MN�9�QHZ��f����@����B�4P�%
�>��#������Ę!�G2���-� ��/���'m��ko&n���d��Y��9K+Nμ�{�(V y�B�Γ�*J"i:������n���V�V�������W��miq5rLx��:Y� ����g��9����c�����q���Ϻ�ƛ������%��,jy?s�'����z�3�2JN��[�z�k_�Z��I��C����z�R��C�{��p�~�C�=���%эl�x$��Mr~v��-���J���}�e�]�2�$ ���JPX���G�oÆ۶�M������7\~��яё�|�+��|��_��_n� �6�a*l^q��7��ξ������j<�;ӥ��X��^����H|��W��v��>!�� V���C�Om��$Ƒܴr��K6I?���AYю�ʰ
]�s)\��ecI��˻�<㌳2���-|<ȳ�������>�upp����P�fA�h��t�P�=oٲe?����̩���VG\�^u�Uo�N$
�* �������>��O_vٟG঄.�;��S�"�3$r�o���3D�Y~ ��W�s�>����Č��r�-����{���\�s�uy�a���N����$g,
P+�v�0�]0o���'�-���{��5�jժ��ov�@C�6���իD�D�}�ӷ�v�1�:G�pΘ#�_޶m��z�5\pʆ׬Y�m�����?�� z�����]�rY�{��޽���r�Q�5�򊳑��DK���Ы�_�l�<i�ŋ��M<Q����dɒBw�zϼ�|>�Ԏ���s�j���t⾲�<aU33�e�2�G#����o�lٲ`hCy��rV�\��ln�d�]WA�9�+tG}��h(M��SO=u��w�qt�Yg�E7E�F�:��W�����{��G<22r�y�<x���xhh�9�3�8c�}�B���@�� �|m��.�\�X��x��q�n��y��~r|��0$�� �;r�LOO�	i!��+33ؕ7���it�&GpkILSq�?���'&�!�ʜ梧Pwm��C���o�z뭷g��St�@[��HN��bGG-�>@A��X�+��=���A���F�9��@f���W�������B�GCe"u|3��������tť���J������7oޯv�ٷo�7[��J3W�����Wf'''�@ζN��F���g��%������ �ojM�Znl!�G}��7���E��+�y	�������~v�]B�d�ڰ�ɳ��ީ�����jPJ�GnٓUuJ��Am�JF>YP@�jj��r	JC�g:!h9�vѢE��w=�0�YN�ؙ�R_7�Q���q�*�	̕$<�V�tj�%ZϺm�=62�s��ҷ�����DG�d@�/b�jM$��(a޼B�ܔ�sc�s���R�,v�5�����6�_g2���̒z M��	�(>�JC�7�����R=��U],v��%O�9͚����ysrv��sNy�N��3'읶[��9��H�����2����J���V��G:��/�}�ـ�T�ѩI)3I�M� �а�S��%�2�Q���w�f��)����p�#��]��(pm(��+��3Ś��I�4�#��������TE���������x��@{ϳ�l�-	9&�Na$�����4$E�	���o����T���1[i#`DkH=� �~�a�ug4��E]d&��P��g?��/~�3���n��af����R**
�aox�EA ��IhN?��yy����������-T�\PzP��[A��p��\�2�ʍX�Dr��"��d}�L|ͅџ�/�(	`F���7����kG4t�J�����:����	�?��o|���t��~s���\�&�/�@�|�1��m2�y#�#h#��$?��������*�vдC�Zf���!<<2r�t��S�0r�5/"7:3��D��Md품+��/����$E)
g�$w��oؽ}�������=-����x�W|�^�7o\�L �	�:/
Mr*⪥e߹���v����7]�%�c��}�7��+>��U�8��V�ttq~����B8�	W��i���m����v�x��%X�dc�J�(��<��s������]�m,Q��S	6��'
g����)2�?;�XV!���]�!�i>iE�M'��� �����t��
�?�;N��b�������:%�W�`�ΝN>�Y��w��~��l57S�T|�[�xӛ^�aA�Q�>��%�������7�|�4�0A:%������ȤQ�����*:]��W_w��hFI�я]��/��?|���KGν��a"�L|�O>4ь��>~ť�C�b����o����>|�s͗4C{�w���;�\Ϟ�;�JE���;����_��G?z�*��]��#K��Vʱp�p�^�?��i��0uu����BA�^3���Qr��cQo.�OE���ʓ�<�f؎=�h���oteA^"�ֳ�jz�t���{��ڤej��2+���m�:ן82
Ղ5��f�g�f����:E~����4�6��blvL.�D�p�H�?_���%#?K��Ń�\/����X��k���:Ʃ\�$
B ܑ@�H��	 �h�hOҠ�~�K���Ã��W,��HLM���&/4g���щ]�ϋMWчw�����R�6�jQ���G-������HQ�i�����t���R6��`_/@��d��E�hox�ŮU�W ��\�r�p��҄:Zl(�Z�&^6�fF��<K{�ɮ���R�6B�@��! ������/����6��3�O~6�gx�!T]w�𢑕]#K��ѯT*���`���h���?1�t��`�p_�`�ރ�Ic���!�6�����vl�,�t�R#MR���6���F����s�6y	�!S�@��
WB�?�3�bV�G¶5b�Q=���8���JgH�P'Ş7�花P\��S(�EƜ�ctw�Ca�ܻ٘-M�3�F'�r9�Tf�
�b
?*i�B�M���1z9�gdDdF�h��(�>��2S뫢���4i35k�jcv���7P�*�ݧ�'Hl5�\�� �����^R���H�LL�]��dRN����>U!���'�`s)�<�-D>`�)���\��5	��r孮�a�����h
�yG8�}�Y�E6�d�*|+�^��Ur�MM�|5l�z*�`�#���4�N�[@c�(%�@oY��TB�&gA�à��=�m�zE�k��)�*��"GH�5r��Q��P1
Sw��[��C�R�b��Ct'�/��8�4��Xq�h���w�������9�?�+��Tv\�#��&R�}�3!0�$
��Z�$~���o��i����۳"�o��FR3��|����i� I3��Urs�CAb�G��n�.�ހ�P˘�*V\�"�Rcl*M�=�3�f��"NI|�NJOCQC�OSS��H����׭��)�}ɸ�����h\�33�f�|�Q_�h�Xě D��d/��=T���fW)��]"��$9�X��p��\Y1����$"��`,�{t�+B'si����U��pf%�L >�DA]��z��@��#w�%)6M��4L��,�G��鑞��ƽ)҃x̀$!�oʥ���ۊ�sa�#FBݠ� �1K���	:����!��H���r2�Բ+���
�.��T_����KhB��$���=����[ZB��JAU.h�P�cCW$�t�g�˞��<T)�e��E�P�"�}&nZ��%SD�3d�G��H���S�8l�D#踩:;����D�֝����t�i�I�!��oyr�;^�M'N�:-��s����Xd��B �qv��@���&�?UhЏ4X�YF� ��`ڒZ�{��n��OZ�
�Y2��t��ݒ!Di�����٬����z�H�{l���蒦�c���|�{��[��v
귉�#������,|��Z��rn�����z���_����|�3���O��m۶S���duc�a3���3P���|�V�W��U�f�-�ԧ>����o�޽�ׯ'c�U�z�����i��M�2���Hw��y����%/B�<�~���#�ǹA�ΫS�;��߼�o�n�4%�Qj��moQt���w��g��SI�%K:t�����Ƕn�:pܪvXW����A��(�ѯ�����;���C�<m������oy�[�b���{W�^��j޴$�?���_|��Ǯy�>����쁁|�y��X������55��\}���ܽ����$�~���8o��v�u���/}�c�y��I8(Zd�&�s<�lH�Hg��[����))r]��޴iSY���w�y�������ɇ�?|}{��[j��_g��K6n�8]-�1۷on^��'���?������'�m����n�t&��C��[;xh������wܱ��4�B�Z$�t�w��Cht�]�n�喣�h���6l؀�?c!NOO�e�8;w��{���t�;�f�����ǘy�M�3>$�a0w���������?Z�v�w��jϞ=����g�r��Etk�r��͛V__-�͛7����ӳj�*��=�tuu�^��==�o��lG�Vշ���4·z����Ou�Q�����i��SSS4�n�H�:�V���1���0%;�Ri4k��eZ����=zO+�����W��ʆfܵ&���{�f7o�[���]H,)����E�-���//������1�}Q,OX����I�����%��H���W;z���ӷ���X�����@�nv�2]���%zz��-ȓ�U�����9�L�.���еU��c޼yV�0Z.ӨvܹbŊ�K��)�'D�����Zq����2y��'��}H�{:��N<QL�N���ĝ�z8� y �>x�y?YC�6#���}�Z����sϥ3�u�Y4�3�>�����-t����?���CȲ��i	�X�Z�ڗ��܃B{)'��s�j�+�{�dɔ�3l YL��4��,�.⺯��M~nYD��.�pj���/0�]��͢e�s�9<���(���߱s��̞��¶y��^��.�L�-�uu=��#/>��������vD3h��G�M��{|ƛ�:/�V����e��E�Yʞ�V����ٳ\�diމ�I5!c4��&�[������{�(�K+m� �'�DJ�aG�����2��d鴴��S�4T,T�>��� �0�$�q�d�fؼw�����-[N��4e����:w���˖Eb���� i��;wӫ���[5`�F�D@�D��'�D�����ۻh�mO�*t|i)�,[7脿~�a�S
�jNT����T=��H�1p.���Y*3-�NQ�*lQ:�y�Պn%����Ҳ7Z9���}גY� n�]�3��{�Hϱ�;T&�T�UV��o���5jO�sZ�ri�?�Ȟ;���|.4HVJZHW�7O�\/z����fT�ª��dG�)e�DJ���I{�+�� ���r&;s�>�h;�3��8�C�^p�V��
}�:��Kڷ��*�I��H���%|/��@%zδE���~�ot?%�+5`�|!�T�� �w��-������>��s�cN�%1�ﱙ��G��O��C�qg#�gx<ㄇeБ����#J�D������_���������W�5�)����[�2�ľ��On��W�Z�O (d��Dq��JQ a���?o�B.Y�Vo��D��%���)���o~}���e�l��5�5�0Nt�A�6n.Zp�W��s�y�{���/}��.�nٹ7�\�V">�@�3^�r��X1t��W��ص{�꣗{Mȅ��P48J����9��XQ�ɞ��b�,��"���LK�H����Z*j3�};wW�f3� �J�^q\o��蘖
��c�P��l�ON�)(�h@V_�V�5�3�Cc�c�������w4^�Dھ{�~�wt�[���q��Yb�f��qf�i1*��!��ev�=XN�����M6t���٤�5SwN�\�����ܿ������#d33Ȁ�(#�/��;;b��|��A��*,�&��n��������у�amr2�����"�7�GGGw�N|����+��8�ԓ�� 5<�հ��\�15rܷ0��z�ڈ2g��;��1���c_<�hӶ�v��e�
�K�ǣ���X�0l��Os,t���L�2Q�EF��$'���6�&)<�5��S�)�/��j���i���N�&��Qo�ɹ�ObF��4M�$v��&͗zI��4%�v�d��;�j���gC+�e�d�Qrz�^ݳ����"H�,4�	Z`�W�)¯*�J�V��c���� �DSH�6�8�4�����"�/����l6
�c�d��5�(��(�;��:�9��h'�ju��}�ȗ�ݱ�8<TP
tw�:��0Ƿ�O��R���u�Ż51Y��� �ܬvwg;ə9ɒ��8�Q���gj���X}ݺ���
	���k�,F,�H�y}�8|̲(���ݝ�?X��%]ǜ|��7�lsO����%E�*z�fiͱ{T�ѓ��d�#♁l]a'��k�胷$L�ЃL��_ʔ\����eYE��r��������9 v"P#��>�gIQ��Q�����܊���ËF���޺u+��3SȤ��^��$I�Y�f�ċB�ZMKk�s��Pr�93��}�7U��ۻn�Zr>qY�a߹�GG��K��e�h�3?Qې����~������:G��W2�)vq�ߚ�8�5 Q'2=��Yqd,!���P������U���Z%��#K3 z5�.Q!���n�&�<z
��(p倂� {F�?A�S�� mA�M|�iOrN�G�a?$��ӔE�'��1f7p2h��`�J�J�|����^:�g쉱������F�`Z8NQ'͐�}���>5>�l�Qih�(>�Ø�H�G����V*����X��N�=%������Tj"p<�Q`������z3�i-U��9#���B��R4á���"N��<a��2V��4T�T�E�x�� �ę�ڙ�#_�[��B*�,�6�d�ti�V���"!���1Hύ}'�u�9^���d�@��72T�Z�B�s���j�ұ�Rq�tJ�:$��u�e�ψq�5�:U:ڇ�W�U���p�o���h;ؖM�V̦�t�$v����΃��w�(����k#�J��η�X�ɧ�����|vm�5��s#�����ٹ�3�h�1��^/8_��~&V3Ӭ�(d�s��,��}����|�5���-��ǁLC�)UU�X�. ͚+��k���w��7����r�y�	�O�^�z���?��ϧ��}}]��[�y��r����-[��|�VS�3v�3t�����3<�?�Ӷ�0*����)�:�,�	X69���h-'�͇����E��\�n�d�F���y��!2���+�-a[b�t9�߹s'���x�i�a�B�M8�"�/�6m*����?���ڏi���@��=�=���͛z�(=��3��5z�t]�yrC>���}��׿^�=IUޢa�J6�h��]Bl�*���<���ǷC?)���V����>��x�y�8��ĝw�p�� �d\��eF��p����x����݃Z�ۇ��ubj��)�s�Et�������T�J��TLOO�'�Ӭ&i���K���А�dv��x
������.D�7ki�dF�ٵ���mTS�VD0��:�c:3Y��������Y���Y"��w��E���(===尿{�~�[�*�Ʉ�@Mf��>x�]��[ɶ�-n���ջ{{��V ��b۶mw�Jq2A�%� NM�T��E�/�[!�-r���k6l�0�|9��f���F_�gտp!���3ȴ��O?}��ե`�ʖ-[h�cG�'h>�+�E�=m͚5)�)m߾���
���,hh.W�X1od$����e�
�\�B�V-R�oU�������#Ðs")%=wwgm� i�"�'�t-Y�r�ZBԳh�D�W��̔�,��z�R-_���L�����MK��-���'�m#_ˬ4�٨�Ӏn��E��5��{���� S����CSd��VZ�Æ��R	�w�JJ�&#xێC�}��4���2=%��Uǟ@g�r�C�ɼy�hziA��&4���1�#z�X�>z-]��0�":qki6<��neE�x�sS��M��pQ�.�d$l�i �N��1h$�?��8ցn�S�ȤEBohS�*z����?��{��E�M ��;v =L`�k�н�쾓�ycIX:���_����������>�919�I�9�����s ���$��jnQfɓ��4��Lb���R��h�К�%J�(���l�G!g��: �d�=�I*)���f�7��!8�B�,�qqtt���	5�0&G�R�f=�L{�[2�`c�^�0�V���/})���O<L+y���y�R�I�x�+O8�E$����v�I�q��_��(@�2�W��7o��D2v��	�"�F���FK[�t���ŋ-2ؤ�� �-ȍ~�����s�gY��O�e�a�~�#�~��ʑI��5�ζ�Z|�3)�Q�:8���ܣ�|d�!"��ϑ�Ѓ�=c�-�qJ;�=�oE;i���:��Ka�,I��nɳ��3t�|s^K�A
��^Rp=[n��}��:r�uwʳ/�����{��y\/8_K�љ6�Yդ&��hy�U߾�⋳(;a��[�;�D]�rf�Y�E��i���~�=����o���G��_t�nQ�\��jZ�����=��g?���t`��<���n�ٟ~��TK�=�!�4�ߤ��#���#+Y�0ȃe��pL����=��v2�W._�D��&��M�b�:�B2D:�źe7b·d��Ŗ�~`և?�W��ß��U�tT�x�0�TO��N��O<�����a �����d1�5�$����\mj��ղR����H�Xpb�W��+�1vp���o�Ч��ο�N~��-[ј���x�5Wox���%�W3'KdKGk2�(	���L�6OV��PhB�:��h� �+�S	�g�L��
y�dpK�$��C�Z�a F9�~'���^���If�{���U��Qƀ�@���C�riz#�Q�2�J�d�k��B��$��(j4����A���X��UHǽ ��wcS��,���&�mN�'{Uk�#P��M�`	"nI���b�2����`L?5K�5�U�|��UZp钆��L��RlDa�{xt�8�{�N��j___��j�� �����y���	9ͦ9�bD� 
��v͈�~�f�sL�I�{��
.&�� C�.d������R�`u��,6J]E#�g�B)+#��Ț�i<���b���P.��_���+qb*�i���q��r��f��Q(��<o�P�w��y��fM�?�^7�9�fM��ř�v����T���iZ����� ���\�Z-�z�p�`��f�Ʃ-��hzD�=�'Y&�i���U`BK*5B��Y�5�I�u�T�8"�ii"0�r�����v�g|b���N�Q]�������Ϗ#��JC���*|]�c��kc�q{�n���/tǨ���z��w@�T����i���� t�E�MWo�wZW��j�ֳ����=cC���B���B��{���pl\���8T��ڵ�Lީ4S�@�fh� �c�{�����]#$�.����ʨ�(u�.zQ�	d� v�ߓk-��LMB�	2���(U��HU�\*���_��E��+��������@p�W��F�r%�P��ϤA��%:�Fx嚣�j@�u����d�tN�P�4�������h�pr����[��[X�d���c+�'�V�\P�V�j+�~�4GHi���t���Rҹ�؇����ҹ��Q�-Co0I~�VW��	�ڤ�X�!;�DL6��h\�{��T���7Sՙ��f�j��=���0 fq
�q�)0@SR� �R4�tZF��\�$T5�4�B�-WA�<r�Ԓ	�����[�l�(�e���6m�V�?�a��S��#?�2T+#>�;^�d�N^z�UAQ.cU���:@�(QQs�3ܶ��vk��JV�U3��8�J��kfm��%5ڹ9Uuw��tT���nr�F�gȗ4-k���ݑ�m&K5n�u���UԷ��2�	�P��3M�g����v~�vs��K&>�|��=���td�䰒�����a̛V�B�Bpsg�3y:�M̗�bS��)2��Z�2W����X���t�^���`�wZ�;�M'����3܌N�Ub`H׈� -J��y�N<�7=a��O.�;;Ł�Wu���O���V��0�U=��q���ڥ��̞j�$��#Z�$KK��rzv�꿙�%^��V���C���D�s��.Y�T�У[6n�����͓����h6\��<��7���O�Eq�˻�ۼy��w=�(���r�)�5���Z�д7�x#m����e��c�}K��s������yr���+�&J���~��+W�9y�8F8�k����珑��J0/-�U�{�w�Vo �B���/D-Gӳm���"#OB�K.IPVm��K����ܺu��ŋ�^�/����D��ۅ��u��]w�È�����Jr9'h�[���?����ɧ>�O��r2��wҔ�w+V�Dx�7��uo	��*Iɶ3<�g�ؒe�ҿ��b��0 pI/�Bq���@�1�;snF�g��.�mY�"����-�>��w��*:|R&K�T*������8�:�L�(X�kɥ���mD \��J�iG�3���Wɸ#��	�nA�K%� "�,tͨ�hk5���h`j*���i�l�����y9g�������7YV�駟�+��
Μ��Cie��iɕ9���mU���<��`^#��e��0� �#CxI�.]j[��I��:+�%��� `�F��S����7�ƾ}�d�ujjjff�h�t��W�^-���wKi��D�m�ߋ6��K�dK%�-:�Z*YX�fYN�cӘ+:�οlٲ���JX4r�M`i��	E��L�[~�Ծ�6�ι��gjt Gǖ��]�2ȁ)���t����-}Vj��L��bB$��\A>�����hZ���Z t|1*"�� �
A�3S���ug���n�9�����{��U^g������3*��$�$�� T���Tcl��>�׿���q��5ql���$��1��i��ޛh�iF�ۙSw���r��HB�N���9�Μ�g��[��ֻʻ`pr6GV&&&����L��5Dcamppp��*�J�a��+�v�/�]���]��'�xb��W���%,��R��ee��`�����$i�gU=�Z��|���=�q���E�hV���PT�i�p�Yc4f����?96NĘ)�)�����1F0j���O=y=|>79���re��FQ0�W����G}���|�+Gy䖊�{�����CI����I�G<gR��)ZTq���Ə�u��T��u���0�=�\�X����m���9�"nrp^�6�HM� ��Q�q��ŭ(� CH�P��V)[�d3_�hfܱ�o@�a�c:C���oyi�d�&��|�e˖�jȝj>gRV/���!�*5���w%��4�{����- ��S��V.{�g,X�N>9Q�9j�R8~��(�F��9 ��4v���׎�T;�Ǿ���?�+���X��^�<�-� �g^�R�ÃO����-H��d�w��o�B4�7�&Ә8k���u����9�{m�HV���!���Ò�*��襕����1��%�>?�A'o�9���jh��Ւ?&5��)Z��_o8�%4�$�U  ��IDAT�@)�t��}������s�{/���n����|��|��P����ӡ�i6Vk�"��>D�e���������쓟������{�]�&ؼ{'�x�#��Wgv"��0�{?�u�io_�f�˔nP��P>�X�?������/��rV���QF�$H��E3�;�8���#}}݉�h���2�"�X�����u3���V*�ãJ2�cM�
v8	�Ï8��'��m��}!����XX�{X��PW�>b�D�ֵj�EsYT��L*Ck_��U�#�G�^��䨷���t�H�~|�>r�9�:��?�g��%���_��_��?���s6�~��p#A\��/|���{̽�曯�d���]uJ�T�Diԭ���2�<J*C�-�*E�8]STY�ͶZG� �*��U���=8
�:�Z��j���+�UM��k��M����e���)9�N��
l� ����8��`�!a�@�/�IL�
�����:������ K��l۶����q���j؅�[�,��BH׋�U��~���ATL}�z{��=��×,������8|E?֖�a����Ju�'��<�@N+ [)��@L*��D�M���������bI1�Ҧ+YMg�z:��{�j��oXF��'���7%aB���"� 	�YC��v�J�(%r1�$r�f'+���)�k�����V�cd靖���r��Cǽ��VZ*��훚����6��mm�e �S�����R���G&�݋u&�G@�JD�ٙ�;��v��juL��)Yٶ��A%�[�l93��$a�_f��+
�<qŋ���?%&����j��=Tj���I�S�/���@ƽ�!ԁ�}/�`N)����}+w�Z쳴l��Ԝ�(NN��2�R�;S�'�&�fK�S�ˇ���&\71�	�V���q�s�U%4ø:>V��d�$-Źl*�ޯ���2 @ ݝ�����շ�F�����Xs�J��_���ѣ`���3< p����˺z�%�n����O�G2F5���R��[�A("r�F����Fۯ^�45ʑ)�PO�u��%��q.�5��#ag|�}�N��Zz;���EU�����:E:i�K5��1��>��fe�U�V��i�� �K,��!�D�Ƹ\��=<18����{Iς�"�<��%�e�6���G�z�<��?_ӹ瞻f�ap�3C�i�L|�C&�f��`_2�C�o2r��hX�Z�"��ucJ���,��v#�{��"��� Is�^E/��n��5;6���CX((D>[ ���6�Ry�2��f[s�3��ٔ	#�Iq-	 �au��"��QT�ؖSm+e1	K�jQ����V)
{��?H�F5-�qa�S�� �o}�i�-zy�n@;[��])����s�7�Ƿ���s��===�{��kk���I�d��)s9r`�4U������yx���AL�*�bb<�r���}��}�g�ctd���xPC�m#ݥf$���a9@��*�;7�$iV��|��s�
9���-���7��������$x��a���<>!g8W�OI��:�+������5�/�1�V��̙��I���`����t����68��]� ��|�L����$R2/ٛ�	v0��p�2�y��/�j�m�����}"���-��i�Ha�/EU�
��y��F�~c:8D��"��c��A�R�ܡ���g��}����|4n��Fè�ah�D~�}�ƍ?��w��w���TGG��0dU�*��Ϧ�Uh�f0P?���q��?����t�7(ί�/�����G��_o|��z衙��SO=նl�u���*��E�`!�^7��PQ]�߸�_�jՃ>��>��Zݵuq�%�\���a�c��q�q�b�GQr�³���7�w�yi�z�H&6����x�m��;���j�)|̝زy�-[6�s�7�:u#Q�L>�g�f���`��V,ӈ�����.���W_}�Wb'�8��~��_s�17�tc�dl�[�|���逸^xө�za �l��N���W��$������?@��Ub�Bv�:���2���"�$�'eE�M�K�M.'�ȏ��f.Պd�YA�B=�1b�k��j�D��#��Y�wo�㥓�{ġ9"%��K0҅�'�>7�P�vG#ߣX���E�I<86@�m�Y���O�j�6�U��C�b�~�m�EC�9��c�4��`�]$sWn�g6�D
�*�N�L� �D
�"���tF*�qV�ͧ���N���a�d��b~�������s�7o��\�l�2D�r0nޅ�����L�k��Vc�uς��+W&��ꫯn۶&�n�(�̀�d����Y�%�b23�3L��*@��M�c�R����;1C2�f^�3���� �!�����Hڭ�cݶ� ��`-x&�T�3�6�PT����:+ed�� S)%)\�NS�<�0X��⋃�o���Ō]�*�L��G`�C�>�4N��`N�	WI �J�tgG�-W
�	XQ6E� ����������>;��c>=1ch+�����_�p�,7L
t*˯Ql�:�o�e�:��,2�ōL6\A�9�%��ݻ������-+��x*��\�JS��9ɲ�\J���gx699�u� o�O�v�Z��0�%�I[!���7��L>ul�Mǫ���O?�yig�����;��ҋ���8� �K�T��:�Lc[�TRPx�A�[#4c�X�k��R�����˽�	X��: �:	Z�y�̇ܕ����kL�\��_���:w�&�5j�ɶ"�'�88��tǩ�&�pc�s*ؙ:�-fJS0 ������#s1V��MR~���ΑFɠ8?��eEr�y�j�
C��b�
��ᜯ�ź`��|d
�Bqu�-����6����/6���^���yI�V�g~�|�ؼ����}�[����#��qx�r�)��%����Z7y��l�|���D3��ޙ
�>������0`�ת>=�q?=��p�����K7����ه�igh=�A���z�a-Ox`� 1:AcM5�(���mڲ�u�`B=��#jb��"���SC����h+�H���r�����zp���}ժ֜v[?�ԓ:4���n������n����W�Y�Z�2XPJ(��U���_���"�i������3G�eYp\{�꒛=��S��;�[�M�~]�*C`#���u�9r�?�|��?6݌mJ��*"�]*�J���O� � ��9��KH^���3�� �P#Q��\]$�&)2�Xd���9}���}��֯ـ$%2�0n�R6Q���{�D�.}�������N�����W�zͷ����On|�%�p�N����ss�ի���t��dG�<��n,�����a�z�����=�p5
�`�:坊@f>qB$DN�`+�B�/ec&���a3F�H�k$�qJ!�^%D���tlđP^�n";E�ũ�R�](1w���]V��P�@�4lmCx�g�@�A�lMVĖn�#�"����V���eSYؼa�И�S��#��*X�T]�c��v��T�`"�p�8���qm{;��k=�p���"�-U�ZL�1�OW�i�65�uJ��C�M�k���K�D}����X�G_BK7"��T$�q}�n�D!5fP�j��!�:�������(N�d҉����	Ƈ�۷�X٣�`��V���O��U�����G���}�]61���#)�g6o+�7e��5ɻ�}11*k��?�|[[����O=�ch`=�g:ǝ�j�m��*F�ҹ�aTw���w�>�m�%��w��'�tҫϾ��#�(��
��-4����3B����k-"�q-1�H��ҫ+3�bV�z����[H'̮� V��F�SK$�0K{'���EvndfăY�T!&�+�^���Ո%B}��M�X
'L��C�@�樞�Ԕ=;F�U�<�B~ibb�r,�-p݊*�]�3����.�D��XUXП���z��oɶ��j������y�i'����`^�L����-��.�r3�m�S<����U��:����a	�qѿc�'4A8�¶�� t�b,�¿�Խp^M�� f��`� o���xN1�Ōlshzz�Z��i��lW7�(�V컠l|��Ł��`j"emp���pk^짳��U�?�\����y���_��+���#�B����lu�;s�瞰B4Φ����G?���tu����kS�l%7�f���K�7(��&=0j_�i?<�z%��3�a3K�+x�y%%�����!f~*)�;��|��7�
�����?W*?�����Gq�e��䛞yӦM�C�_|��+�e����7�Pu�c�t�E��<(�z������x��iút�����m9��������m�B�ǩt��\��A[ h�$�>�2W�Q�%�Pm�� z(�/a��g�S���6ۀ7Z�+NO���exl��/�N����]��]o?�%�-T+XC��Q�@����
�L�2:�����jqi6(�u����{P�W�f�o�e�1+;::LS�=J׭���k�z�F��½�bg���}��d�+�:G�JD�� '��Vp>�Dm�d�%c��r�P5%�;��2zԘ�}ܒ�QG@Up�B�%�-�쑸���`(��_�uwFM:
H���TA�����\'�Qjh����$1�_HXYS��b���ٛ2���SP�:%��cGd#��bٹ��M���=��l>�M�w�h&�s�w�lk!d��&�NG���ٌ|~�h�"|9����$�
�dΟ�/y��1hk�ǟcqx�ܗ��* v]5xFIR�d����=�Q(����pX+nD~qR�JuݺuFς|�W	�c�|�t�Ml��$|4~��q"�l%�^w��7�3�N�d��y� ��+�iö-@g�-���������m��v�ig��)�|Q�?l�y2���e��V�/��(�1�B�,��j)5[�v(�_ّ�_ad�PA��6�$� �:A�D��f�gҸM��q��/���\s͒%K.~���k��L1f�E�fQ�D'p��k.��u�4�4͙�͵̶S��^u�W����3���5k֨>E���]�v]}��p�+����4C\}�5_��o�����}���5�������03�j~���i��)�E-M_s]p�r��x�^��oL�?���(hdbڻ��VD����"e�~�5!�n�42G��R���kP<'���#&�Q	��uE���Q؉��y�Q�ҋ�/��ߖ�D�
V�H��x��9��(_�#I�m�!�2td�O���	vV�+�ț ��B殉inUĞc����*�Z�l�(�F�;
���b��[� �
���Bˁ�_�4X]I.���EEJB�6���Ɉ��^��V-b�!�ϑL"��ډU�V���PN���xHUp��:���n���r�
9�=?�m��`�\F-�M�����r�[7�`7sD��h��z�)�D�8U���17v����啸���
;��e��S:9b%�d��k5<�1���Q����*�������~������J-W�`B}-c�V9�Z+6fff����`ah"<u�H0���X-!s�"��.�J�J�_�ì98	��|�I��8���W�}ߪH�����c�m�;w�r�
��Z�øaÆGy��������nk�E0Z�J���	�)u`�X�~q��p]�,Ea�@A~������AxS	* Q�=� -V=���g�6Ʈ�j� �S��}XE�X7�M�N��? F;�J����ݻ#�2�(2�����(�,mmmp�0�y=�������|��8�y($U�G��]��[aaoijʡ��]]�_�6r`N�!����I�6sju�B@P��ú��F����\�t)I�l��"����U �۶n��nٲ~r̟#��ה�|M�*D����ڍ��d$��˺`��L&��-���X~��*ܭ��#cc�*@9�t$�e���cP� >!�鋼��əD�L� �MM0 p_ݶ�g�0l�T��!=F�%�ȿhn^�?����� ���G�@�p�:�ʗ��"K^ �#%�	��wi���
#E��Ճ;���|���G�-b�>�Ѝ;���� �/��[��w=��Ec~L1 ZA���Ma+��9�p��:�J�Xb��4���Q9��$F\�ז���9�M��@�®ȕeۭ�&n��m![����Ӷ�������1kxc����)�E��W�`j��!᳃合���͌��\������M4��#�����#M���Y��;�i��wַ���o��5_�⵰�ba\���g�o~��sV�:��P(zc-Qh�����៾���/|�qU���v���z�{/Xܛe��V����mo��~��_�rhh��_;�H	�*���A�K���k��ˀ�4l��r���a�
aq����L�x@nX����X�u��f=���{�W�����e��[\Vvņ�����B�?�zˆ��|ه?������'���<&|+:���GE�SP��&(E;Uu1���ُ�v*y�d�@�}�.�a�C)2S&�`�H�֟�������?��/���7�4����~�_������7ޘ����^��O~��o|��o����'ȼ�
�X��ڢ��N:�{����?p!���Sa#��?��<���'�>��A�x��{��1ʙLD��D��"�R�$j�-�NA5ӽ&\#c܄��ڼ�b����+B{4�,�	UtʁVF�mB>��dlG� �r��U{��ktP�d�I*r��1@��d&�n�PY��	}��j�B^��mf!�Ǝ�Rq�̔��J[{آ�by��G/ �ozb�m�EX�R�<�pFL� ��1�b#C�Òdկ�����65
6[�@�
���j.��j�=9Qj~�f뒩0޺���R���YfDw�R�l�p(�ɒk���\0FXXo8/dZױ�[Ɇ#"�H�sn�sbFu�!x�瞦
��Ffx�B�~n�v0iP�۵��3/a��
�L[G��H
�R��`D�p=�"^���Ǎm񂎩R�3��L���3�l�
�R������:����2N�0</�39ee��0���W���e�9!��RdlEˇP|d��MQ
�ːel�%�,� >)�f�n"��TL� ��˴���lR�B��{``�2;	@��.tt�"�?�
N7;<3����2��|��ٝ���"��¢V���n�*��75>g���]r�-�ڄ��kA�.`3F����+�S3�g�\���w%��Ό2���VShb>��yky�Z�:�`ԓ����'^xf�Q����c����uֺ���"W��xB��1�4F�?����6�sj,���1,=�U����D �
XEBBU��we����9��^0t_�KcQ���׮^������-{@ir0�R���b�nʄ��O�
���K
�5爞�֝x�֭[�������`[�nf�;vm��n[�t�,ab��V�/_nW<G
9�R񬫉��J˥�*ԥ�ʀ�e�����ղ��&����x>$�ZS���\���-�Y���c�U����-[wn)J��C���R_���v�<�c.�������W\��/]�eϯ���[�Sg�qV��ß~�Ż�������=�3�[�؅B+wfnr�X�cR��;K�Z۫� ����A���*n=�ϥsYd�t��q���o�^Q�[I�� ��(r�ЎcY����'��������Q��	@K`���j��+�z{��Z���S#9J�ntC�MU��W�C.W梚��Yz�yo9��w�2 �rƐ}l�X�"�حa6p�G�z�Ǣ���Ξ�b��%��ix9���#�8+�ѫ�+X�N�$f<�?��rr���-�u�ؿ�7t ����;@p#2J�s��t��:��;�ՙ(v<c�r�/|X�R��NF_�y�o*)��TL�!?HJBu�@�޸��V�k>���(c9D����8$R��6W	c���b�(����F��=�+H����it.�H��l�q���bZB^)�Qlh��	'Q��~R�#EY�\S�	�\	ּ��J4m��)�)�=������b�6�B<��a�@D�.l���%�v�(aN��2j.��$����l\B�d�=&��l�#�F+���7�_����Z� ��V������_w�u��o ԡJ��G���_ 0�5��+W����Q�u=��������ۯ���/_u��GP�v�M7݄`F���b���SN�ⳟ��m���~:Xe��4ݰ��X7����c7j� ]p`��|�~i�4���>A�.�|k��9������=&7{�`�Z���1�^[��F���td8+���M������㏟z�`"d�K� �US	Q*-�����s��_A�krnn�x�xm5(3�D�Y˨~IE �nݺ���io�孷�~�/�6� �iP\_�����S#�%p�������^z�7^�)��xHt,�0���پ�����	��/�A�k�?��5MfF/�w@6��m�Y�/�0'��'���Ko���F�l�+����  ��RKWj4Y�Z������9���Mi�q!j��Q��2�'�;M�kU���S	avL��RE�/���L:O��f4zy	�L��U�������Z3۪蕄h���u���r�QTUt%�I�Tjˤ�H�X�d���sl�J��q�C��t��k�Eoe��{.�m/"S�cd9�r	W�gf�+u�
)�`cWgs)s�E7h�:�P�������)~���mb�[�J1Ceb4;333�c�mq��ʘ��м����Sֶ�;��jIO:�K�M�J�s6�߫�Y"
j3F���$N=���ed��`����r�7�4���"��>���Bg��q�\sF�����Z�g*&_��p��q���ou�Cԥ8�0���"�
	Ì:��zbv?q�
<<<|��'/^��cp@&�����/�JOJ���u���C/7�Vc���s���!rWV�Jȁi!K�e�#���	����^~.�H)�7?�����ڵk��v����u��|��w�J\����uW)p�"��^I�7q��p�	�-��i`��V*m�;��u~jꨋ1UM����L�������69��4�0@b�T�%�b>OXG�e��U��WrP�����_z�O[|��e� �zѢE���s�>���xvN�1)	P*���P(p�,�������٧�z�^���{���/.�O����9�W�����uï0��v�{���F����/7Z��ϓ�A��QJ6yqc�؅�4
�����d�sɡ�]��ze6�N-Y�$��Ub�}��8M��ĥ`��;22��9hE��§� -����U�4��8ۜ-x�hy������Q�����2��T-����O~z��?�qT��������}��t;E����~�я~L�mt.�_�N{��ͅ|���bx��7�������� �ѩ�ɮ�?���v�-`0�� �;��n��N�S��H��82	�
<QOo�7��͋.����*�������d��_�z�{.ͰXj���O��(E�An�Q���V����l*���}�	9���9޻a�xk�
���ؼ4��k��Wa���bFI%� -� �;�4B�x2��x�s�J��6����9��ƴ�580p�I�c�Iף=+�{��|)s�|b[4Hv���y�^o8�%Gr�@�b0?u��]0X����;�5�*.����r�B_�d���aɦL�)������~�cw�y �L������7:A'�2��A�dU/��_��?�y��w�}�n�69"B!���E��n����a�����U4�2�����c>��I!����M�,Wf`�	���e����F�4V���7�Ȇ!)�qgm�V��{�Ȭ��b>����s3[��|�	'�A�6�egVҴk������АQ@���\OIQ��Q̡1���%QSe�_�-UVB�Ԣ��5�z���&q�O}�������'I7Գ�>��_��q⻒Glٱ{`h&�e�q%�Q
��7��o����������s�]�l�Vv�ʅO=���݋��	�i>X�:�'1��q�ss��j�yje�c1Ձ�I,t�J��E��|~��W���_:����Q����sK���e�2F�O(ӆ��ց�`��AU�l!E���9�Lp��D-����{:��rJ��Hְ�tZ�]t���2��h�g����h�R���v�NK�lq�B��I"u�X����~3�UܶS�c�O0sY��SGf�T��Q@�.�Fd%���kձ�,�aHu�A(i�3;P��juKE�q�63�˚/��aP���="�܂ě);MX�9�Cns
M���Պ�)��) ��-\k�Q�������,Er��S��*�]��ª��X滁A�� ��t���&�v��1�����tZ	��ZN�t���\gv|�Z��}`ŢY����	s $@:AX4*g��j�a�2��?���?�uilq~��@����,N"j��i���FS�#KI��#V�/|ɐ�+�<X�N�:�հ��W
a~E�+�kk.B�- �Jun���H�@�N�a��vڵ��HZ`jU;r,G��K�Bש�$3c�J%ƀ���L���zVQ�x'�^	�s����`=ի��=�vzax����/�>�c#����)[�ly��"ב��a�(zaeN���6k�$��
C��-�ذ-=��h�ZE�Wa�*Y[5u_��S<F�����=�<�j�L5�lɆ7w'����;�����=ѹ�99t}bbb۫ؠ�s�0J3��S۶)�3�0�)�)�Ѷ�e�:"c U�BM$Yd&��buvxP�KJ}����p��J�6�0�=�s�Qՙ��X�<�K��YPs��#��[��ּ�Fz"���Zw�*�Ɋ�f}�eM���u�o�:fwrp�=}�lfL{ָ)F��1-��S����^���[ȷ�ɳ��7n,��0˾����>��2�����'�r�%Q��4���ֶ�L*4�!��6]�S3�G�����4�"ixt�h#C�]�x�QG�4}dbR�T�kR�cv^�����H����|wt���:�J�2N<Aġ(�PN+V���R��x�Oի5�zrRM`6�z�jd-e���t{;,\y\���d�S?�rME�Hc8%�P�fFq&�R$��0	��,���0}��rm�}�0�8h���c��|��b�rO�����4nrJ�q��8�p%��ϝz�Q����}9;C�ݻ��8�-CB]˨;h�(������F��K}���k�:����iyN��}��5M��?��W|���&Y���R*��s�ݺ�}�ʫ�򕯤%�`p
�.%9�ЇJ��E$��Y�T0�����{�U�h��������|�_�2�M1��R+h�v��d�����ҷl���<�̾�j}�2�[eR� �-��g�r���o.I��b�CI�fttD��BE��_��obt!�d��fR�����}�s_���¹��K��췾�-t!��tڔk]]]_��g���Z,�&k��x���$y#Ƭ���k�2`�Я`0��n��V��)�`_��p��},�p�Tp�gk�a���v{�y6�tb�[:e��a��!T%��_��_��߁���a�E:UC�v�u7ӂ[슐���<��8Tş��e���|v�p���^�F����l����GW�tDN�2� �N��K��Ig֯_�-C�@D���8��9���Έ}W]t�Ƌ/v=��v�������\0T=/mXt�!��վ��o~�o���]S1h@��U$�)��J�(�<����5�nT#����k�qV�~�_��)z(%��P��i��"��$���Kb�w���W��}j�d���Yk�U�Z@�:��8�@e��^��vGGG�a�
��Rbɓt̗�%;�ݺu������4,gN��mʍ�|L4�k0ѣũ+V�/^8�+���ח�n-�tnxx���~���B�Z�-�_}��0�ZCC�jO�q	��T�ڒ:Pe��J�J�\���p�+~@������5�O�|�`6!?��8<][>�nj)fi�3�XI�(���62O$^8�{�~_�<�֨rH�|��%�po@ƶ��B���u*�1Z�H8=] �c�U��N�e�q�ܕ�,,4Y�1TdtXf�ʢԈ��5�/�pV��2��g�X��$����]��� �x��7��U%i< ���dp����[���7�9[� ����"��1fY�l���9U��>-B�H%���q�t����j�*��]16�Z�H0��z�r�ŮY�G�1���۶m-ah=��}���+�A�\���c��#�X���
�B�-��Q���`���w�ܩZ6H�Ly���I�6�
��T�U#��DÄÙK�
	��1�Ay��`�s��0,p�)���1.��_)�2�,��|zhh襗^�g��V��'�����ڵkW2=_�etoy�`�F-uH����J�+������˗i]�;v�������<����T�*��J*.C���>�,q�x���^�d:��w���yu;�g���<�O�R��b�O���_~v�ˠ�V�]O4::�hѢ�}��n��~����n�"�4���)
�T�e	"���cx�|�����-������7߼f͚������[oc�3�M�)�F���G���[�*8�_�l�����W�\��ÏO`��-[*�K%7�ga��f.L7F2W4�qAA�B�|r���"w�1�~��s��pW��33ŒF�78l�����@�w�A�1"<&���!^�B ���&�߁���!��F[Q(�z�3�8��=���oL0�4���_���w���GM(��#��7��� $�^6�?���}��߿���Bn\p���9|�Ǟ����9����|���	�W~��~��߸�:�K/��4�a� �|0/.��һﾛ뢱@�N�~����dtt����}��כvD��O�����n<���*1�ƾv�- $�}��3�a�����]�$hU�p����[�P� w�l�Wkָ����#i����v� ��M(i�#�	|���������_�zÆSJ�r!�}��GO9���|�;��.xR�ky���ۿ��z�'��N��SO>w��'���~�;�y�/�49Y� ���pXK����n��P�����P3��e݈@�K$��b�|�RC�"+yղL���'��Yt;��Q)�K
�(�#�H{D�$�� �^U��Kd,R�T��O�4��U+��x	����9�UX�F������C��̦��6+�J�?T��";��y#G��j-����p�*vU �K1}��*�ɫj�z-mf"�e�JdC7�p����1jDb���[��f���X �S�|=
��Iرi(��CU�i�J{��UCh ZeL�Q���O��n�c�j˸S�ޅ��j������Z��Ô�b(H)|�e����X��ׇM=m�Ĕ�mT�m�t=��K�$L���f��+!����W΀eTT�ʊ%������������� *u�RȤ�]����y {��JS��{�~�%S�������[��](K4�Cߋ�0�=C���5��a�G�Hi�r:q���bם��5T����N���y�'�>=>3��Oı�ۛ���&ż�ahs�%!S5B�e %�k��ll�)��幾��d+j�2�Y%ck���R�T�5
e.r�-� �����$�E����X'�����T 3VG�ne�~TY'���Ɋne4�1��H�l�!�qu��Q�w�H��(&���e���*�SVރ����عA.U*�����B"�HU��t��	�p�ԤP��}zbL%+kh26t1,#e녰-�^(9���ɝ�ȋdQ�0��6��BU�NLO��a%[,qdDn9Q���&��0�a.�.��|����	v-�cB"�@v))�$[�%`[�u��B]R�n���,~��Ҕ%cW���T�eR5�Т��K�$w�
�*�It۾��0©0S�{�ۊcN����R	�Z�4O�(�ґ�����Z�FgS�P#�Sic��"E��/����F���VW����d�r�TK���Յ�����+))Eɂ�	�"jl���U!j�e�`4RP8��L���X�T*3c#����n9�� ��E�l�N���	0_�d���
�^q����nݺu��v��},vg���[,Yrm`��[�"�jo�'��jYW(����,b+MK$t��&}$:Kw�&��ޡ�G?_���#~!��Mۂ�٥��HN}ժUq&700�c� ����E��`q��nf��&�?t?=�.����Ԋ���e���%F�b��sr�֝m��i�~��fS��� zђ�ޗ�|vd������U��C���5'L�ro�]�S���~�i#���f�ʕ��>���eZ��l�F����:����Ζ���D��a�c����zL��Fv<&R<Ѩ��rI��)�|��ȇ�-�JUR�ׯ;���K;R������^�^09:::ז�׮]���:��z.���+/�NÒ��ؤ�]��Edx����09�7�3��읫��銁��ȗ���NU���Yg��|����3���L�8��v��n2�֢-59�X�x��?��I�7�rn��]��K��?���.��}�����_�|���������z��M�N8q6Z������u��2�v(������#{���~�0�sUTXA��i�֠�.���Lƺ��{�>�M�z��dZDe������O}�N��O�ٛ6l��T��嗷l>�S]Y�p҉��lq|f�w0Y��{�R&�+�q������/�|`��5k�JA�|`��	�0)Ȃ�gD�.�V�7�0v%0������&��h�ז㛭��W�c\l���f�˭ԤʠLH�����J���u�^x,��}�׭;�7�φNp�	'|�����ؽ��}��u"����
'̹v�Z/�d���'�p�~��?������'Ǳ��y�!�7�d|D�ʺN0���B�Ԏ(KձOe:i�� ��Ҏ���)R����(��r}8UKNgr+d�Z�a�߶u�]`C�B�� \��Zx���:�y,Z����4�,��r�)¸��=Fx�F��l[�V,/�{L��P&f%��e���Z @�8j��2���it���K�)����F��i`�9�v�a�`Ġ;M�d޼^;���k�e@ �0P�*�X�~�2f�ã��w��:\Z�|����1`Z�N�d��ȡ�;5U]�i����Io�l����+��b������N̋h�(`\b_E�ω���*��Q�6w(��WuC��jiP�"m���FFF�{�����a�^-�:WLҹt9��L�����z��[Ƙ,�����ҥKs����<N	�v��{�X�n}{{{��3�Jm�5��=�^�`�y�O|���˨pNc��Z*OLLd�P��l�B�$�X���}}}`�cV�e2��!t<LL��+	��Ӗ��c�2v貱�K�� �|����s*����T�h:�F1�|�'Ga�t=��øY)��<�'�L�¶�K�
y�����o�l�v�!��1,���s�"\+[�1&V�����n�3�w���S��oL�I,K21~�+X?�.I��*,������=�!��7�w�����j��J\Aq�1�Y�-�'�� �'#*�f=��&w�����V��
ʳ2��%�Ivp<ҋA2Ѵ��P�~q4����ҫ�LS5]ԓ�f��ݐ�Ҙ�:>�Gv�xcT�`بs@K�������c˃�{�.(CI��ͥx�c1)�BX�I����&#� r6��Gh�������N��������I8`fbf��
���&>*O�l;{.�X��?�'��>�l	kj`��A��R}ӦM9���ES,v�b���9x"-F�$��%�ɋ��MM`mY`��2CCCv��k��K��оx���Lerrҫձ����(�x�8�!���Kp5Q�WP���ar/����tb��R����:j�
0a���
�2===��/��2X��l��c�}��G|>���˗-���?mS�?�w/���]x�QGUJXkz�ᇿ��+0qo}�[�X�l�a�}�v6p[)a-6N�����XV�Ĥ�	Ç1\�?�ba����������s:92���	����w����a�?��s�?�} 4Z/u��ٍ��4��YB�������×\|�I'����b�oe��-������t��*7��/��
ǜ�ʰ`s���nM�~�������;������?�|��a
	�mt��UW]��ff֬Y#薘��G��1�G��DUÞ�) ��m<;ܻ6��wo���ᑫ���3�五�㹆.��;�_��_��'?y�7~�OJ5���}�k�l慁w�y�ǯ��k���`�L|�wƘ�������th�S�>���iA�$��i/�-�U��4i�E�Xe��Z2q���h�qG��_9���W��خ�Uk�wqlXV��AеD"Ԍ��W��d�����;���G?�x����������Y�}������d�IP�d�����֡_o8��1�s&@B�Z�A"����X �FDqbY�����K	\	#*FC*�Q#
�GO�/��J������$*h��H+��B7 �W�`���}���J�H���f,�+���C[��X��Z�<��- �Ǵ^�Iؙ ��F�}����2���դ@$v�L�����#<3Pd$4uL�*�}�66x�o76��zy3�l"�,9v����$T�TT�h�aľ��E�7�P���6v�LՇ��`:�U��,*�� ����8��	��[p� ;�u$DL� IA�aWI�1���2�&��Cr{� �>��KQwI9j�&/�'z(0���nIF  �ήʰS��I~�l���j���(��n�6�,h�ejI�x��k)ӄt�8Uǈ��fW}�/�G���k�m�tKn�x�F�-�6eLˏ5EJ�F[���,��d��]�G(4�dR���,����pld�Ƕ���ܒ�l+AT�YF�'�|�7 ��!� �# 1t�֥�X�+��YП]�����n8ޓ���#�����%�fd�
�{J3��Ӆ�RI���� `�벥{N2[+�p���S����X�J���5�*�q����f��܀͖�!�Q����`��TմnVa��A1�u7,a#Tx����C��i91u93j��ZRu�_t5��5�h����r�Dj�J�%A"u�j�Z
`��cN\��R�m9����*Ȫd�1Q�@�Z���B?��Q%ҩ��22��Ŧ��pq��.Q��&��4M�bMN�%a����[�S%F$EIY�f� ��a����ϧ*�R�XE��:�iV`u��Z�3��b-3[T�^ֽ�S����k)�Q2�bfC$�U�v$Α4����6������i�m�OB�i��;ǧ�,�*V�P�(����ku�6�j�0�.�H~��w� ز�c �n��RC��U�⢶���c�yhl
l%k��]�:��g�ڵ�[o޾w����Z�tiW������E$������?�O<>>�}i=g����m33�~�<����j�߉�(u��S��k92L&O�PZ0#0Ɂ�>,Xnq�S��ryf��Ksq�����^�j��cV��<����z�G��T�;��u,��3��1��w|Z25?g'����d��]�D�G.�D������xS\�є�-�9�*$���7�����J�@�s�j�'���E����u�������� �5;�ccc���"�î�pj�?�-���dP*�0b"��쳰��`�%b�T|����{O;�Wv�q{幗`�7�L�b? q�Ͷ=3]��w�l8�5p��3��<���c�m����@U�X��j�E�42\h�`�b�6�`�º\teږ���p��u@ݺ��O�3�x뙅��TS�{��D����'���[ 5MO�����"*� ����飀��E"�����vq�+��˹gy�*r[)�L��ewvv����R�8��!Ҏz9�+�3vR$CGw�a�e�o���v��	(k �������i$�!�����6��!��.��˛"]��w�V*�0mP@�nVYK��r�CO?O�?��{VVu#71� �&H����N�с���bпj��JJ2�q�Z���W�d���>��] �tÔkԩ"�k|�[�t]{��g^�$;w��_܄�-�n���Z�h�g}I��L9K�04$������<���?�B�O�2&�G
*�ԧ���u:ir��MRxѬ ��=�E3#W�GqԨ) ی�i-1���E��Ͷd^����!l	��Ԉ��ҧ`�
���렀�����\�$�����'�� �kVE����#Ʋw�e��ǿ���(&��p�X�ؕT*�JDP/��@4�	�)4�?/z���>���C�2���Ԭϑ�O#�~ߏ��m4o��2D��ʼ��сͅ��Bjz�S6jvy��_�F�r��0��,t��ecE]����&kn�
��U[n�-ʷ��� ��$B7Tm
�ȡF��=�7��}��yҌ����9������1�B��⣀�ѸvR��������������H��|�d�B���A�'��TF�QLFivVU+e��b(�c"�L��n�U 	aNi��La��6[��|�%dǓ�_{$�aphN�ʹ-X�`ph솎�.���Y�h��z�۰2G�+�}�^d=�@�m�*��O<���g�9�������B̆柯b&�jj�}��#M�a�wѳS'���W5V��=q��p�q�m���@�w�Y�c��z���۷����Y��3O�����_|qb �����	�֭|���������-�YP�V�x�a�J����;��bM���{l�[���ԃRe�b�|�S�e1��COZ)@`6�	Ǎ�*�+��Ñp�A���H�"�.>�Nue(*�B��y�z�{I�<vvv�`��U�vd��F�1><K(Bn��4k���� �{3a��f��YIҒO�N	a!�+��
O�1�P'J3�`,zf#�E���\�<a@��x_G�"��*����gm��N�g��FQ;b�Ք�V��qk͞3 ��E~@�
�]�F��j��le�`��`B�J�P�/���'��k׮ݻw�a�d5�*QP���v�
��k�BZ����.o��뮻���矺���bŊ�N;cӦMO�x�ц��T�rq��a����ѱu��ݻw�<j9H&,�nw��7�F�&c�B���s�$F����ѭ����N.ը�6k�ТE��Zijj
`!O�nF��cf�a��~��r9��bժ�M�T]�P������!7;D��XK�q�L�b?��?dk�7�C�����W����ټy�\��Ni	�&=:::>>n`'E�湴�����wg����b[ü�;`6-)�R�g����#���A�����Nxs�]�>��c��=�sT��2��[R�����q�⨡��I0��� �������o~�W_}u��^X�G�Z]�㨩�������W��́�u*-�B��檑�a��;�y�����������+W���:Q�S℡g���|�Wy�4б}x�4H���~H�l
���LVk;;��!�'Jy,�l+{e�%n:h�\H}�)�[Tu��C:Q�KE����$x�W}����y˻υaI4o�6�4���.K�Ν;aؗ.]��O���[�i��2����L�(C�K
��B,S�R|��C�j2-�P-�ݛn���8Ձox����>�(m�;K~��z�v�?���o��{_��[��hbFn̚�%~"�xr�S@�������O}�������/��T-	���NX燾�"�;��3N;���/�����%�\�qc�����=t��'5�$��4��������,߲hl>�\�2������>����#:�ƹ���&�~��Z�yY.L�F '2��[���w�_dW�|��?����Y1n��:>؂M�H1�{�`����G�O�'�=9�Ӫ�r�	Qw���#��б���!!y�Ǟ�@�����!�A
F���8bՔ+!׏Ҵ ��c$<���,l0a�d���00d�
l� ��1*S9�L��+��!o[�� �!F�i��0[�\�p���VJH���h���a�j`jh�n4��-j���|"�^�r�W��ww-Ȥ�3���ֹ�KUw_U�%���Ҏ!�ț��ܾ���稣�"B�6qL�S�8��U��U34�p���� |��o������K��;���y v�L[�q}Ӷ6lذu�0XuW�f������Dn�^p*���V.z;����OD�A��/�v���k�]c�U����N]|Ċ�SOMONςn�ȁ �2Ƭ.���I�����F��|�B����G���?�<��� �������Pq����ξ�,ջK+^ܼY�}�\̘��9>`1i
�e)Hb?
���$M��`L��c����]DI����,u��aM�����ˀO����a]8�����8
�-�; Y�es�������x�})�&Y�B/pх�j�
�@s:0O��䡑�2g���֓�(O�ؼ.��:��I��$S?��0���\rD+�F�X��t˅<�`��}�[�Yu-[���݀C�J�#�8b��k=v��"
G�g���g�}ʒ%K�l��� �P���Z '�de�~T�5P�Θ]َ��70��� FC�Hikx��p'U���n��wDZ&�Xc� �&���i�2�ٔ�Ij��U�\!�U�Z��̀�2L�k�<k�R3�Ӿ�`l�����^p�1�#S�~�ol����L�w�F��Ф]�ٶv;��w���W\�bŃ<���p�Ks�ܱ�,�$F%�V�rP�h(�$'��R���˾�
%A`V��,� (�)u���W�?��ܮ���ּ�ΜsNFB $LI AE��Zp� (�U�K�jh�^m{��Z��Vk�"��2
"�2H�<O'9'g�{�y���{ߵWvNr�����E����5|����;�~@�$ymL�Di��DǶ�Z������6X-���Y��i���y��!�H��4�'\�^�Yj�d����4-?�չ���9~ȑJM��]q@P��o�Ҳ�1�Su� �e�`����I�T�,7�A-�{��#ߢ'��R�l� w]���# x�%���J�e�gU�Lo$�3�c��]�F��̛4I�� Ftr?����,L[	"�<��8/�Rop�s���ʢV`�0�<�|�Y�Y������l��h͚5�O\F�9�"h)���.A>V�-'&5���n��,��X�?~�Ɵ=�j���K-Z�bEG�w��\�	fS�(l�L�Q0ӳ��\G���u!&�������tN�	$͍LEm/K��$Z �rd١ � ]9{��˖��S�S)���'7��w���@8{!m<�_��[n�;�nEA�oy�I8����ܜ���בJ�[~�:��M��_�r�)��b2�8�Z��T�q�UFn�<�������LyZխ��L�I�!�F$�J�F� j6#10
6�'�>��5��У]]�dΏ3���ř��ni+�W�Y��,�|����N�P�����2bәD��DϜ��l�M��ӟ��5�nժU�p_����}��9�]w�G���(���X�����ч>~�Y� �)n�Mt�/��3��G,�is4��c���$⹌֬�����~R�tg��9n;m�̬��y�;R��1Ҕ�h�G�񨡦c�1���K��젳
;�d��M&��H�Ѧ|_��a����<�~��z����cd�#��@T�-h��;&EY����\U����TOꆛ|S���VQ�J�X���i����r�<�@"ˋRi���v{æ�2/�v^��JM:kx����X�Ĝd��||�!>	��\--I�Os�a���[�Ea?��i��Ǌ�w�@�� ����/j%SS3��'}�%�a��L��3���3czf��׼6�u��=�L��(Λ7���]�v��Mg3�Q��p��zz���d��_�s�Β��d,w��t�-[����'˕��e���Ҡ��Ұ�عi۶m���CCC]NM�JPߘ��\��ˤl\.'Q�?�Ӑ�]ծ��� _⠲� ������AtgXNmQA���-���J`S�U�z�diW���;uW���*�.w��(�YyB{-/Ү��?M��̋Nn�Y�h�i���.�\�<�f����w�9��[%Ӈ\t�gw>�z��o�>��e(RX�2���-%��c���x(�);j�p����099F��+���ј��Hb�\��E�5ˉ�.X�735E�l�2zL:9�$��D�#8L��j�b�dz�A_sZ2d1#+R��y %��0beg��.���'��#C/�-�Jl�$��K=�Hr������s�*�i�%#����H�h�~i3ff��/�Z
�jpgm�$��OkC�=ۤ�\�;�1]��U�_��'�E�
U����x_������L+gtlV�� X($A/{�h��9%��i�=@��sÓ�=%�&#&3���a܊u�ʜ7M��� ��$�9���&#O��~�J?�������u�֑J��4+Zz2�v��C���E�o��-3pLK�����G���pZ�
��SQ�&C/zDɐ���J7:5�,%SN_��z�9E;z�����ҝ�k�q@�a����j�l�o������3�O��k�f���W����l���&�r�&*�sR5c{�CiT���AG�'��,Ѩ��h����$7L����r���$%_�B�_~�����&�����5�\s��W�t�?MOM��(eU^�c2k)��9�����f-�R�t��Q��E!�a�)�N
$Q�mك�]���Czŕo���;�	����ϭ��@c4H���;~��2������I/�����f���M߱��C��Z��!�5��Y���j�:b7���XC�NrY�Kbɒ�*��Q�Kh�b�h#�+Ud{K���8�@˛ l6���<|�l���&D�)�8c��L�6��A�B�K�6^I} ����� 5Ш�#3����,,PBlkjI�X^`qyd�. Z��r��B��%F�� 9�W��h�A�4A S��f@C������;7���A�J7h#C|��7Ks0����i�-ֵ&������tbH̫@�(��;b{�d��m2�3�IL�E�U[~��zw�P�2Ar��8"���knW���1O\041�l�N�90̦��MOdZi��4'{kj�>�9]���Y�N�$i�i�E�hVk���Lě���ů&�[3��I�MyПNL���d4�8����wu;���m���Qj�s�QX�u�(4�v���Z[������齛6m�t�@�ɴ~�+��;�ص�{hp�������;�n�j��7<<���M;&'^q�˖�:��������O>��k��v�i�D��_���V/�?�ҁ�����u�N̴��u�]7�?����7Հ���:���<�#��5`Xf:٨zD4�*�c�wC�q��366���C6t�2��`F���
,5}��#�H� �]j}�l�d>�d��̿dX0w4[�M7e+�f*��Tt$�i���7$�����ƙCC�/3�ΐ�@S5�3�:�hr�����-���44f��d�8�9*�bC1!���l�L���엽dŊ��S�y���<s����.�t��3~������<c5�(f�}��wwe�E/z�3�ܿ{�=� 2Y@�5��X�>�_Y0�/�C�]�u5ӈ�����s�zU��ܝ�Y�A��t�	�Y�M��J� sОzA��	B�y
N
�p$�3�t�Fnݭ1Fk����'u�i5�F����֜w�u��>4�n�ګ�|3��}����z��ɂ�_�{�VNׯ_?�c�4�~�q��_Z��)_o4�||<JR�&�����d�CWR��3=��Z`�ΑtF8�����i�Y	��MՆU	�8���]NS%T!?u��M�-_���o:6�/�1�ǑU�Z~�d���9Pr���FD����؇ SD�5��luX�3�X�L��iX��Ca`�\�yu0DE)��"vΫ(o�-w����Z9�"UuP4k��AˬZ �#�6/Cg0@7��/�f�i-�d+O�^�EbB���,NU��a��%�EsT�"У8%�2�[�ܹ��xT����Y��Etm�a�:*��4�T]B�`��;7l��X���|��Y3]�|ux�Խ"�D�Q�Z��9"#Ҭ���Twvl�غe�|=c�C�y��Yk�X������Ź�7+6=9t��"}�J :`�o[��18?��K혾wd�S?���㞃�����Uif�aY������WB�lǎ��w��Uj��L����n������������I���0Cdhɼ��&�:v-KR̴f��{t��KW�b	�d��ah��� ]y떝?����'�`Fc��Q����T��Az�0S�W�A�UI��*H�v�x�U7}������;'NX�;9��vY�M�X���a��Q�׹:�r�ʟ��]g��|�yZ��N��ZՍ5�f!v4��jT�
�N�g%�ηn��.�˟�}�K_z��o��k>@�a���9�.�Z}���Yy��������?���2�$���a���8����=���(�We������9�ZG����X����2��y;L">)�i��cD?�S���]H�[^ֆ��;�y�=��kZ�WݑH9�u�uiS-΍��%�#���O�?M�4k�[��8K�iT��L(�2Ny��fZe��z�H�Za������>�A;4�|��Z婌�	;9�:+���`x����d�@��?�]�55o��i�|*NiͰ����R�*�3ڰ�/c�%��X�h�f b�kI��C2���f)�)���%��)!��C�ox���$��`�"��t������-B/xE� ���k�>�m�lw�7*�G��̓���HJ�/��y�,YB�ݷo�޽{�6����6>>.�Q����x�K=��,�/��%s�F8T!y<�N���)i=��dC�d˒�;�&�P���&G�V�n%�ɠJuJz�,B^��Qg�u�t�B8r>lň�1:.M�!"�$�:~ˏ��0
�qoo/�W���#;~ÓO.]���1����D���E����'���9J���z7��q��`��	���W� �A�R�39��x!ԍ�	%�­�O6˅38��I�+r�t�9&�'�$mЃ�q�ƆSA��Y���/dѕ���-[��}���ͻv�Z�u}ݺu$��GD�K.LpL1�!�:�R�b�I����?��IO�{勱��A4��L��#�Y����f��ؼ�6Y���F�;
bAH�'O���MQ(�i@M֗$�K�C�ݡ�t϶v���Q>�jgu���Jid�eށd~8瘅�����V���iP���N0,^���a�έu���].�)��8�&y�B4u�TABo:{b��0��(�´h��'�vO����,^#J�/U���L���L�H�%�)�B?��+�y5��Y���s�qI/�T�`F��*���:�̬��������#I%�Y���{�9��SS�	�)�h��,��D@/��S�RQ�U]�8C�u+	]ӵ��J�<J�J�n������������VA�囔cY�y���E!?�&�O�d����Fo�U	�$��:����O?�����aR��F��r�Dq��J�m)Ê8�b?��q�6��8�Z�K;T+�@.O;�r�q�GV�}�>*���Ѩ�}��4P����A@2i�|��պ{�}�uW+$�IР��i̜s�9�^z��ߎ�%o�R�:���#��^_k��ι0�}Z}�<
��p�r�-e;-�S�r��Z�����1�c��o��"q��(�l��t�uXǸUQ�be�-�@<o4���Q���*lg�۴LJ�4�,s�Xk�q}�)��<�t��Q����QHo�If�Ʀ��[��%(o���&������L�E��g�>Ҙ�$Ox�m����T�.Us��"T��1fE���#C��^V3���ǡ)�����a�ʰ�t�8�r�M�c)��9"�&9���0 �y
\t2L��9@�f���N���<�Ϳ|l�S��}p�@߀�:f�Z��z�+��/�hŹ��}ZʡN4p|Y6C�c�e��4�����ɩ�z���@��t�d�,��x3rϬ(��8�I_S^W��h�x��4�FԌ� ��D��t�Ӆ=��E�ܑ�R�����ےX0y�.�{�z�z���80���������~/�V����v�oܰ��'׮]�z@]'�s�و��d+K���c҉��,���'���}�E�C�Y�k��۾�t�^����N=������{�0w4۳<-D��qD��4Q���q���r,��id���"�^���_�`=Ҷ*�2�U��MuJ=}��U$1h6] �'iNۘDIĖj5�-c�����WX E�Uɲum��X�ni��&�ײ���5'	++�鏑����v�����G:9'�qA-O:Ӻ1nN̵%iv�䕡3���Wl{|��ܳ΢���{��͉	"k�6����{~r�/��U4�=]CÃ��l����sN;�e/[1�����>15�k{�Aj4DXb�.ƭp���Ɓ�&w��a\��MRD����&�p*�"(�L�m�5vzUJF�����3�29�i(3˛���CN��� ����8'�_@����{lӶ;�m"������0M�=��/�c��'z��m��xMU��O�p*�w�1y��i�;�jF3>)�+J�t�E3�ʋz�������1`Md*I݁$�2��\;!݊VU����J3�v�=L$>���}6�H����dc
�Qt�ޮ.ރrq�$�6�ԺH>ɐ"1����Ȉ�p	��g&�v�B|����"�ò��:^��04����4�2�
t��i�^��x����ݮ�MzRT/�Z���1��;�|��hS �%���QҌZZJNrr"M혴%G���h%0�I�9���qL^"�Xw�[$ou}2�����P���Ѯ����K��FC}��i����F)��'�Gj$�+pI�>���FN��y��p�!�ةn:]5��4�ϱ���_Z�*b�m��
9�A\���;��X��J����8��	]�����ٖ���<�9����t��_v�>�������<q�k/��޷o�1S�u��Jb�6�$�� �}^M7�th׋-�fҬU,`�z��i�f��iӧ��qd@�&U &�����~���^x�g�]/%sK���#}u�5����y�{ߋ�#�S�5t��h�8� KB,K[�"N>����{��a�VJ1r��-7�B[A�9�=X7t�[�R�/dj���˄������Y����#�6�b�1�G�z���Z�8�@��s�~��;֯z���YhZ��P'k�I���\q�R�F3+W,~���_���W�K���n�j��?���k֬"A��[� jw���峎<~K}�Yq�2�s�C��C�+���ov��β����ã��E�)&�}��������̄?�T\��y�gsDo��1u��������h�R�󕷩���Y*u����#��y�ܑ0���Øֺ0Mg��"H/h�r�c2�P��V�A�{N�$3PD��M�L ЏM8���<��(�+� ��tm�}��a���6��V�R�S�;i��"����6M�����OI��g��z���U��H0�f�T�k2�7�JKp�蛂}g&�$�N��7W�N�n<�A�%� �V&ƙP?i�]�$��a?]��"�%�Yo�-Z�p����i�D��0 ����ك���� �oe(�Z��NMM����?�xO���� =��O�۴iS��-5KFZk@r�$U�V�x��.5f�Rs��	CW�~f1`i���6q���'I6���MS�t�/�0�qL��Dg�$�.0Tr��ۦ�����i��k'�t�g��E.۪��J�#��̯�J�>G���X�e���&��;���픺z(�ꤱ��̌�I�;���[�r�'�8ϫ��5��/�U/�v� Uq�B#�3rI�Hm/�����r3e,�"ɨ�Š���k��$D� *��L� |n��4aZ�87����3,CAt*"&ٿ���Fr��*3!JL���|�4L&''�z2i@��K�G8��I+r�s�ȳ�!�f��5K�]���s+�45��
�����#�vA�V���`69��3-L��Fa.M�_�$8�7��~.�GI��8J��@�0�rG�����m,ݒ���d�N�2Y$i"���6��u�=�Y��D���4�7/UY#R�(��$���]�s��_��Z$�0H�p`E4I<� �M�w�v����[y�lO���4��2E�2?�ŷ@'����48�����*_ڛB��8Ro�ڿ���M�PC���7�|����UW�8��|���^��G}ꩧ�ܹ3K�]�mZD�(<)�R� �a(}R��u�=Ҫ�u��/~�.<�E/zի_���|G3�<L�J�?��/|�yj���oҢ@gr�h�E�j��`���A���7��o>����ۿ��'?�dH�o~�{���տ7o^=�Q�,�0'�>���O@Ͳ��2�J_B"w��N�i�2�{�*M�戔0r�|.��������;�+_�ʛ��Q>t��=�l��]]�DW^y�w�����ߺ�KiY҉�$"�>66��w�����F�G	�������o����}R��2�:G"�kG
�0�I!2/Y�h��2G�f���jz��:g�3�Yq�)�p+�R�P��E|��ʔU�y'�>ѹa�o2�̌ɛ���y�g.���%:_H�E��8	zg�,E�\I�Yh�a�d�o���h�%yB2Էh_���ox�e3�-]�����w�{����Q3��V�[�h�'s�~FФ�/;ypp�?��ޱ22�rF"��%�\r��w�9�27���.y�7�h�. ��B�*����Z�bŮm�1k�����]�U�.mY�������������tv)��T��6l�0o��v|�B����h�E?��qI�ꐥ[�@Je{�
1G��0�3�քNK"R��*]վ��X�q�,޼sܦ��`qe����P�M-��ҡ����:id��,�j��'q�l�a�^9~�	�?�����T��P�5�j�
{)~+$���蔕'�ӣ�����ߨ�����$ly��>������_<��Y�{wHg9m�b��PR,c�Y��R��3�<��S��W�n�޷L�^z��C����d���ɃSz�����ׯ۽{7yP/���N[0�70�s�����u����rmz�uO�[�ĺ���٫�X�t饗���+V�9唍���qm_�v����e'���S�Ӧa�8���9�<Kc%V,f��0H���de���a'���\A�_a�+Sܭ�N5Z伥 C�1�����M:o���\x�^����K�7m� �Gzl�����!%+�A�r�hT���A
g~\�M_�= �<�euej	�떩�qB��p�L��@��2>m	�e�M\�F2�Ȥ��(k��-�%A�׃;:3~�Rɀ�$Uo,����?x�`���5�ԫ��S����{�~�;�}���뮇׭���{|��5�`7b�pw�H��b4,�w��O�7�3�&&P�j�o�:"��+ϙ
�UM�w�U�k>61�����kg����d#u�����0O�<M����.���h��6�������t�6o�k�^q��h�q�i+hf�o�F��q������кH���N�D	-�ٰ^׹~@�L�-񙴓��$g,N�87�Ŧ��f�	`?�X��{���h�-Z}�=}Ѝ�LCM�Oh\U(&����Ubht�;��)-��$�蟈k��n�Ѭ5�1�{���lr�9��h(�Ҥ�3i\-������c`C�Sn�"�p�ւr�s��ԡ��X��X�H�PMZE-�L�sM��q���N���.���(��/��ZH�:�MPeM���O��1�	)�H0��?b3�;��L-��m b���ӓ9�i�m�E�%��xb� -?#Y�a��L��,��R! �5��c6OPk/%�LzJ*�����a�B�𾪷�mx�`o/�#�"8�C�`Z���(�V+Z�9z�w���'��6ׇy�
�匡����;0�K�Sjb3%��:�����wۋ_�ʍ럜�_�p���u����O_��\Ӝ�VYWx+��L�J�M���̆�U���m,�<J̊&��/��������}�?��N�si�<cr^=���?��+�x}D͖oU�j)�@)�b�y�O}�[��ٿ��_~���B��όU�W����D��"B��K�M_ ٔ6�U;�v����#���ڱ��U�@Վ�U�2>E�a[6���d�h�n6+U����wlذ��������~�{>@'2�*�8Wk�X��^&�eDox���?���~��o��Mo6��N����O?}�&-6P�H���(n��F��Ѱe�T��,�#�N������=~K}�gL�M�����M�z��_}��-�H$�*�ƍ7^�>����/��W�������Z� ��舀�c��ӟ��W��߼�k��n[vX��a�e���LE��$`/ɋg|����
��E��N�`��#A@��Ƕ����,*�fLd�ka�ַ����|�;�������,���$�u@lM�4-Z��~�j�i�|	�#5�8�fӳ�s���_��d�/�Zͫ���?$����O|�O�͐��,۵cǙ�w�`�� {G�#�<�dɒ�[���5�$��� 0�H�����v�,�5�V������
�������ek���7r��;v��u~&9K������(ܡ�!)H�T\�A�l�
2H�Vss�Xt���Kp4�X��`�Q�/���B@d$ ����(1veJ�@�����霪#m�� <�)�6j�f�k�FqY/G&8����կ������'=ȼ^SIF��P��45����pŇ�DLA�ڵ+�Խ]LҚ�ݍ.���a��<�T���Y;�p��vN���=	K)��u�G�Io�D%o m��I$btt��n�+I&���5����H�����:+�԰��]|�Ӗ�Ƭ��7�b_k�Éؔz@��������RB�Z*�d���z��n�SД��|�rX��ʕ+{�zz�!�B4�4)��Hr�sh6i:H �q���4R��̨vC���ʒ��X�W�ۉ[�ϣ�0��W3oGC��3�<d��� T 7{�U1�3	ڷ3��h��=Hޒ���iz�>NN��%"#�vw�R�_�;���*��nU���$�����O�v���N2�a�q��I9-��z �A��O y�H-
���i�T2�ʤ��Q��M50���G%��������r���e��$��I�y�IDF��;i�H2zEA�,��:�yzo6m��7���}V�ռ����JgB~?���v�ow^i��8�����]E��[�%�ٹ��u\�a���p%��.s�J+�}��)�����v �,Ky�SI��f*@s�n2tjv��잢��c���Xq���s�p��?����wQj��F����?��8�A�3N:㿨p��a�W�U��Rb 2@>����b�|ժUY�����җ�&G4fo������/s�Y���Tl�v���_�X)�pW:��6lx�%W�qǝ���I�{��즛���ǳG�0��#"�%�A:��tV�!ZE�+颴:Jo��s�Z�t��vc'�#�#�H�9��昐m�_��__���?��ϟ>�j"]�7/���f�Q���O~�k�Y��<�ID�|�+_���KD2�nv�IQh�l��Ciw�$my|}n�yd�+�{�-��x��z�#i�� ��3d
<��z��q��$(FNH�i��o��+��|�{_�6�-�h4#���b3���m͖���]F���ܐr!u�ͩ���\�b��4���|��/ٺ���NWA�8�mn�E��v����%�2S�q�$y��?��O$-�[o�%Ң4O�8%3�ԕg����=9�B�r�k��|��_����mn w"���c��������go����Eq�Ś���=R[֣�<��w����_s��7}϶L-B��{?��/}�����I˗]z՛��G>�ɖ��_��?���y�f������߮~��o���Q�ݶ5Jz�f�V����7��-o��[�Z�`�+�l�T�ƀ·(~ٙ���eG�^��axeh&�=X�P�SSk�V���@���=wf|rll��ð���*F�����5S5��KS�fl��-\�5�·�k�+sЩWsC�n5��-���bb Jm��͹)�,���>��*��oݮ��gȓ��(&�D�v�>�o��Դ ����I��`�iy^���0�*Ur�b��L�2&w����#��[����_mؽ���ޡa{��������o�:�����G��ٺ�@��}��ᅚ6��k�b�d�ޡ��V�fڰ[�,���I'������j�Hs�r�/��E���#��������`��&�I�L6\��j���n��t��+d%�&t�Ν�?$b����lt�SKNL:q��"��}�,�#���41s���~K���t��^�
C���o�rR͠{%+D�h�c.�i�5�i�U,;���XV�<��@n�o�V��w�s{��]s�)}�5�W�/|ɋ�/Z�g݆ԛ j�\�ӻ���̬�Jm��OL�Z��K����ʽ:) ���[��i�j&�<�Qx�D7 �s�s�*�^��9F�yP�K�v&�Ì�Q���=g��%��V��(ٶc�$W�Z��Y��qJ��K�0:?I0Y뺩M��{6"#��z��Y��8���FŘ�jM��=~1]��̉���Qz�MU	��5ж��-	7�H&�ݶ#@Q �Q38Kc��銔l�����`E���F�J$`-<��y�	���S�c?(��� ��	's�<���Tr��G����8cF\�x��xFa�ll-
�(�}���5ܵ[f���-C�R3���� �,M��F:0.�KyEX���,+�6�����hphA�����P�gF *�M�o� G��¹��J�t%�i��#xl��+9 B1�-�H!����{zz���G��駟��:�700�1��㡐 X�2�a��E�2d�hE��i&����+-O[���j��2�]=$�z�wG�5��CnZd��pl@�X�L��̷�g!����I��H���ć5
�E+fz��(a��,��Ӑ��_��$9"���^D�kp�
H�,Ƕ�w��[��ַ�ܗM�ĶHy�amۤ�4sݺu�-�Dנ���m^��i�?��>�7�9i,c����d�m�]p��������\����r,n���!
��{?�����Bl��TaIe�P~�KC
����#±����K�+^�sei��qi�~-
�{d�\���8��8v%
�%Kݯbch��3kz[����/�7��0U�2V3\��b��0�@���l��_ha�!���o
���4O�Pk�ѓ�HX�mן�:Z�9_��6[M_Y$|6mnQ��iӦիW����@
��(��d�3����;[-@x����o�?���%�	H��+~%�-1��/V/:d%�XRǈ��6�񬜬|�̏I����L�YDa��Lh��w�3������o�]�j�ZXn�m����۷��o~�w������w��r]�pÐ��r���?��?_�v�=��tb"X��"�H�TX@���UW]Uu�߿��s�9'ό$�`O'����|�/~�+������W��뺏>��+����%qKֶo�喅K����{��?�ν�Y\Xm߲�ܳ�g�E�B��u����:C)�[K;�Uf˯�Z+J�u�2v��%�K�?��Ա�l��&����B7F�<�U�V^y�4δ7�ݾsjjj������I'�m��3�ιs�~�hEɾ����l�޾.������]��ħ1\�x1�m5˗/߿j���#c���e˖�v�i���tڰهG�*+9n���n���,�R�S!�L�B�������O>I3"��������7@(�h���/})� ��Bi9�N5�җ���jrr�$j���w��n��� 1���X�t�O<�u�`tÖ�5�I>2����^���L9XE_��0�$GDV���tř���͛'5�tr�W��%ĳ�H$S�M�޽�ޤ�|f�a��ӳȸ��X��w%(_Mh�.]Jג ���ð�tdZz=�IY��mt2Y����p�_��Y�6�];*_��;��SߥCv�?����G��{������N?e�޽{��x/I���_\[�����>����!������nӥ�#7]���_����r�2F�-�=mHV��#��u�=�Mԡ8��EWX��G���aʅ�:�����l�LUD�}�Rz���5��cͳ����6�Wj�]���d���g�u=������N����rJ+��'�h�˹/(����Z���Hk�7� _:i�r�P�޺�l?+
�%��L�zجm{��/�0n_JI��5�y��������'r%���?}���z��BzQ�������z�����њ�h�| �6����s枇�x��d�49�S�;�Ü��T��E��+9�"# ����y��V-a�'�MG��*�@RF@�+�Lx
���)�jO=��MČt���{���o��t�V�h4&H��m��O�ܶl��M�]7���I}{��$��-D����2о�~�v���уN�?@���h���ꁲj!g�������~�l��!���ȿf�V��<bf}�����՘��`��jR4���x�H���ޡ�u���\����E�9.R���X|-c�
Q�t����x�� �j8�U�i�m[~�Z��B.��w$����-�֥:��0~a4�	G�����	}!�AY�[6	w�ǟ�<�j���,��$�*�.4�	wtKŖI�-ɿ�Pm&&wh�쭚���8�d�֛D%���U�4�}��ʏ�b�z�����Z�(���m�e�n~8��o������G�J�K��$�4R�,�_<���g��U�`ɩ�tH-��F���]���|����첋ixS�[L�#c���W^x��U�6��,gN��M�*:W\&)I,沚���Q�Yu���j�6��zγxC�@qY*}�1B=߹�];�}��������V�G�5��s��tv��>�}�9g�����9=y0O�m������͓NY~�O6�ͫ�&��V�y��9�
�[o�y뾑���� l��;��7�H5.���O}���ڿ���}��e��v��Ԑ3�8h��S�3�:��{��yd�& @\���������o#��y�E�0c��N���A9Z�Ua�ʄ	D0��9;d��"k��`���)˖aJF���;��J�7�����zF����랿p�]q Z�2�j��$�����<��ɧݶk�����~۹!�Wy�J��?�ަ�c'\�&�KӬ��������O�}�vh�����e'� �1W�֭[G&���QQt�?# �L��p��VD��� D%�zz{�bv�s�!�U_&���)�c�*j���F�tC0�e]4o����i�z2��䏷ȼr��%�-K�Hb-G�}$�P�@�N�6 ݢ}Ԋ�J���)�t��t�0��&0�=#E��:9/.�ȳ6� �@ �m�	�a�.Ai��U&�R�Hvm�O#�4F����:��rJ���t۶KB�n�f��I�[fl�`f4	˱t(��e#~��f���f�V�>BLwF6���'
d�CRʍ��ꬤ�ft�L������tw$:aMƺGEe]�gݺu�t��O��7�}g�{�ڦU���ۗ��9���4��������0tP`�&��N���ˡ�+�(��b\��dhQ@�c�FM�uD��#]���f��ȸ�R�]<�Lt�U�(\�r�˒�K��e��z�rM?	#�֕j��U�6`�i�Ь�I�(.�ê�H�@��
�#J���t��d��@��_�_U�vQ^�J,-IY2�g�6`cB�P�{�*ڏ`g�B^o~~��s�<���_o����v����_*�(@x��i3H'� �
8�O�M�'M�h����2�?�֞wx�sZV�sn���|Fr�N�$A�L����S�1q&$��К�8��X)���cV���тy�7��_�j~Ң�M�<gRt3�J:�y�u�	��V+Uc�脦ҫ�b���a�[f�&~�@XBG�m`�y\-FX�'���¯2B@�F�LT_��f&AJQ�2�]�hт3V�>��O8�Dұ�x�q��}��;v옚��BO�*Z)3 ����2Ә"w�� �#�t�Z�q-��x��Pw�%�$�{�1?��q�
i�ZZ����[s��qh�.�V��6��㶖�U+u��*0��oNMn��gzu��z�=EfN�[�Iۑf��ġQ�6H�f������Lŉ����3��\�h�Rf��(����2�x�m,+��aO��J�)M��f����v��
y4��:L��SSf�f#`�dR����D2��ig/9j=SE�QPա�O
�g9HG]ZG-���`
������ҬS�7����\H��a�;p 5V9T�B><�@���8Ad��t�>m��:b�UҐ��D�n��c0��a��	
48M����,VQ!5��ۉ���T)y�gH6�h�`��@Y����u�o����z��z��QN6&�0vm�Np��g#�d�D+�"�v�gI2 �^u�U_��Wo���׿�� 
<�I�����j��\s�z�1�%fY�F)H�2��H���ܗb�u��ע,�l��Gx�JX�#����;�1 c<������U���Iz*jbr��Q�f#P��/��'{(���G��@�J�f��0A�]n����s�U�^c�F�.Do^z�QU��� -��Hu3����W�r`���69ݜWA�%�
�c�n�O���5�yMooOB���Q�cZ��>�￼�;^��7�}����td�K�)���q����y;q_��#ՠD��u��ִҘ����x����ho�`��(!����!� 
���G�hѢz���. u<9����Я�m�F��u�.�����s�o2&�T#�y��.�������g�uV%k֬y��+�:�7@��{��m۶��{��G�w �]�$@���2�nsc��!�]9�_�8U�r���+򛰩�EfQ	�sB��pF����8z'�%lFӒ"�k��0(��	���Whe�Z"�4&�\
�E��*�aW��ڨ@ �wh�Sچ���$M���(:?M������M��m�g���5��8��;�a�Jz�NE���@�T`i "ˑ�?�LG��u��>�b���jҭZV���Qd��3q[&�����Z��#͠�qˮ�7����#�_G'�K�������+���6l r&AYհ����{R�)wB���:Ǐۥm��U�DHZ���:��>5�!���<|;/�A��ul�n�r��m�?pNIԦ�d���S�J�V�xӴ৖l$j�9�)�y����=̒���X��,���%)&�?�V�l%Hk��-e�8�d>��&'�6m�D�{���>��Rp%�{��#H&]3W�3����X/	�_�,��8:�����?pt��CѺgo�hܖ���C�*潏�$��(�A\�^������ =�V���+0Wt}hhH�M��PVTe�ۈ����ݷt�q�K4>�ڈwK���}K0j��J'���w�\Ō˴��.α�ֺj�������_z�	'����A;������h��K�,^t��ƭ[i����B>�e���8F���dS���E/<g�ҥ�G�蜭�	Zz��/[��̋+VL6pϏ?�$�qO�g�ƍ�Kkf�����t�<��C{�֘�5_��~Ԩ�L��ւ��٦U8i䷴yM��)�E�t�Y�-��=�<Èt>X��[n�_���h圩GgD���Fp��܉$gr�\�9Ε�V镥�ƕ��� `��9#�GAlV-���R?f\kW���-�糂\�P��,QW�ݏ�� HK^k�0z=/� /��SVJ&5x��,)MĪϑT,ӼZۙ	!�@g9Z@3�/(H]�Qh��˽I�_l�c���!�r�!Ճ�,�Z+�ٹ�A��䐯	�g)̿!��s��3��2qh�g����=;G���/X��ĕ�����Xu�)w��#]]�F�T��)+OX�d����_��/�b#�c�{��~�ig�uc����5 :<�e�nN�,��O�|�v��6����u��O�Q�2y-��bjhmR?��,8�E8��d�T~�Z*��x��z�/^z�嚹�����Q@]�UIՐ!�X�JGXKϴ,JUD�Ŋ����������W����+*=@����Ps����\�U���Q'�������4̮�e[��;�؏��U+S����my����7:񻯾س��SܦM�q�t�'��sV���k�E!O����<UsB�U{����~� 8��C��x�ܭ�D��Ooظa龉	2�iߝ��zl� ,��0hM(c��6m�D�n٪���`7=��N�#��k����_�Y�k�G�޷�i�	ZU3���m���7m��tʎ�=�v�;�֪}��ç�j�;����kzx#=��CQ	��ltb3�mg��z�l���!ϖ���iҶI�t��e�8\�b�%٨ؖas)��XI��s۴�\1WRQ^ʳTϹ�2�%\��MF������-G~@֨�QF�4t��B�^ࣶ�I̄V�r`����"�2��D�d��L��mB�,����I&&&h5�u��FC�b�a��L���F�0���&3$t)���i ���b����ь]=���D����U���#�d�	ic�)�ò6�n)g�����o����V�#fJ�'�$��j��H\�YL�(H������q������4�I9*[DuX���#����$�;��O�y��̑�0�Xi�0��$���� -��/�nv�٧�ڼ>0�r���H��-��:��u���M��=[FG�m��OӇ�Yςn�_�-�s��;����ha�ۼ�:}�f���"@Y��"���x�vr���f,���b�yF�#�JŠΔ����)s�	94�Efz��9`��#ӓ�I�7��CwۥCf�4P��E���0[i�IĞ�r��M4 �ى����Bw.�d)�t�rt!�@�d�3<G��?p�Gpt��OS�M���,Nh��b$3Ьچk5��`0=>�$���V6=��2[�1aH6 �m�8����6"*d#��Ǿ[������X�ض��q�8������n�[�يv�z�ꡥS%��z�X��&L-�uc���ZBƑǇ+4�B� ��YJ��6L0@T����{��l۲m��6T��������i��ח�;n��Gvl0���;n�E�����7�hڭT,��ؕs,3�ØvP���h�����ϯw�3ͱ���������.ZeA�1�Z!�n�⥈�MM�߿߾�+n��9���}q3�_��睝g�-���>?�Ta�*�Qz�V���)�s�n�E�Qya�s�]������I�ے�cS����� M��j�R@w��r=~��r0�,xk&�,��z^ٯN�AQF��N�\#N��Ĉ��x�F3誴=%i�ΰ�g�-:�K�}Ή]�����s�Q4Yi��\�!�g�t��)놊Gx&�9%D8����l���^��q��p]8WF���m��
f��6��i���2�ɮÞ�Q�Y)�Zjf1S�"9��Hq3t\�P�  �yP�J�/�**W�V`J ���-��ļ��+}E1J�?�]P�U�@��)=�y��ո����G)4Ѥ^�[�����~<CbJs�iӦ�[�nђa�d��}�co~�u?��%�\(��G��o��TX ����AP�P�\G�Ag�u�����Z�yc��H�V�]�*j�b�v!�T�*�py���I3�r�aY��|��>ǒ jP}��|���4^���W���?��?��/D�ꫯ~�;�I�B����G��,���|��*]JY	��Ok���V�KLB۴�8���s�r�a�R��vӝ?��Tb�d��ĝ�>~�������~���몫^���w�k|���o����.:���q���=�#Ǳ3R��I���� �֮���D��Ж����i�\��>69CO�3<���7n�S˖-z�.��������dӁn��jZ�F��K2�K�� ��`��_�2}�r�Jӱ�,YR�y���-���ݻ~�v:w,��:�C��!�?�C���irVy�Dk��344�jժ=�c�=F����ad-�dax~LAɟ.��1���q5��r�xTN��h69��Q�Kg%\)ѯ��;D˺ NrledAE��4�x��b9��8Z�<�Pea, �8�i�	�z��*��$~A��5�nEҶ���g:CH$�$��l0�	�y/!���#9i4&�d��L͛7�������W�DOd �1�I�S�&'�7N�	��,[*�tyjv�Q������5��n��[@���D���4�MdX�Ⱦ�h�9l�F�
y�TϦ��q*��
H4m�L���>��t8�g�^ʕU����˭ܘ����C��f@R꣦�#J@D�0��J� 9��9ɭL�l�\}	L۫���b����h���e5�am8��`�&z��1w�������-+3����B�30�9#��@ �~X�G�(2���T�a	�����:�\X]��4�Ky��}I��`������c�����Cw �Tz>����$U�>���}�	��Pw]�y�4���e/%�3��m�`���"2a��]�~�D��y��nߧǟ����պh6�A�gn��?��;R@�`��m~�[��+=B9N2���~I�1]�n��Ȧ�N�w�y�-�HI�ڶ�������ၡ!R�L<��ӫ�8�fg��������F�Բ�<A�	2�k�3��4Y�7o�.]�TEM�U�3�-[�[�����	 g�:"_�Q"\Ԋg��6/Z��u�{�v�S�D����:����g9��A�3J�P3��|rl�ܶL��Z%t����l����MI�r%��T�!��O�X��F>r��?d���䙐)�+,Bn[L����Ix���[(�u��c4T�7pم�ě�Xv��N��s�ʴ�Ê�
�$�� ��.��:՗�����O��p�J�$k���"ߡ��:�����_;+?��!�� �Ǥ��;�:).A���8ü ��a�~�'�M��<���X���8���������pǕ����|ԓ�~6�R~X*7��n=�k=�a90hk�*H����6Z���u�}�P�`�z街_p������r�?X�g�^��%�������^{>��-��Ʒ��U��{�eVY������z���Z�y�Uu���6�'�N�d��.�<��F��PQ�+=!]�vz��c�2��:?�%��}��n��I��Zd;!BR���-Y��ߴ�0����bA��A*L��d�&�;_�f�}����j&w!X��F��\7D�+:�U��� L2{�'U!���߄ZW�B�)넳Nm�Iw
��n��+�n���?z�կ��?��q:�Kq���R����̪\v��#�ɵ�!�a�i]@A�/�#L�?V�����4
��L�nK��p�]CX�=�S�1�U��"�Dż��jt�ri��:qV4��eVfi�Z~���3af>x��&#���n�[�G�
3�!hy`$+��u�
Y�g��LZa؈�y�q��|�\,���>t�%�,�Z�4N|�2r3Z?V��[qO!���\EV�����]t��c:=;���*�?���G���~�)��R�����8�N�F725��١�I^�2��a�$�탧��)i�-t?�+39	�q�`�e!�.�&}`BCh#���I3d�e�[#_{0��̴ky1Wۛ��c�Ǩ2S�2!�O��b�YG��tC��K�^����J�Y�I�2�[�M�
��6�(HL����:������W�d��+N[C6JD�1���jۦtZ��:�3t?A�|[��3Z�u�/%#�$MH��3�Th�)
�;̘�X?��g��v��k�XƑON��i�m$q���|f&�3�gRZ�YO�ɔ?5�����(O+*��N��My*�P�B��BS�����АG�C��#�R�R�}șr�W��1����˙�F8%��0�f@g�@,���¬��.�з74���3� ^��K��޾�����M�="�6����U��"7�4�э�Sե��h#5+f�;5��(U��F#�l����^��w�,�鸁�,�{y�m�V����#2��ֆ2�9�g2\#0+�LI��I��R����/�v_6w3N�.�Ekٯe��I���VI����V��Ōk��K��&�o��5�*���.]����N�7o^F_����9}�+^�;<H�j���]���m;OZs��~y�� hv�@�/^x�E�,ۣ?�mbd��<���҉�n�J�lo҇���N���cI�I�8 �Z�0�ŝK�2�&IV�L��8BL�|ks�[�꟞?�pw-����U��ܿ���d422J��eӾ���w�'��{��;���Y8ܝFS~cU��"� �>�çe^Y��j�6��w.���G�s����孠��e��q��:��ȼ%'�^��w�M_�W�VU<����||�Po3iѦ�!���h�P�/��L�U�T�]���u�eu_QM��(gk5�I��Ta��m�ke��EF:Kh_��4��E��h�:)73S+���3���8�ͼ��O����4l'PL�æ��*-�F����T!Z�����<DV��>t�]*бE��� N�e�UN�SX�*7��QdP��C�U�sA|�1���=�e2!�+�w�6�Q��a/q��L�2�.��J?� FX@�kn���Y�P*���DV���D.a�6GO [Ƌ��Iu[d7&ʈi�,�r)hV��x�H��L[���\$h�\���ԦA{s�ᤈ���}�|xKN��x��'l��2�J*LH�j�Hh& ���M&�i�&��ķ��,-���>6x3N��.�<�o�Q��_{<�k=�!q ����[�A�v���XN�6_t�.���}�{��9x�C���֬YC^m ����|���]�t�ʕ+;��:}�##�;i�\��#K\��P��U�۲i[��R���Y�z���v�Y�N8��n�駟����aS:v���7��7��Mw֭�p�+^�(���F�Du�M7�@����I��J�p#�i$1���+&�Tt1O7<�Ԗ-[�V�JjO˙q��;�ݎ��?����N¨zh�t]���o|������O�3��f�K'=\����z�J+/}�K���&8�Q��;�yԘzg�I�Q�M�_�Zd�Gb�Z�c���H3�AkK�;b����C/\,����$�, x�y��e�Q�ʈ="ƽ��*e�� �u�P�{zz�_
�F#��R�����ǌ5�,��868�3��`a�C��������y��%�W����A�C�q2��m�8mc��@��J!��'EF���ѧw԰�������M�!���qG C*a�rJ�^�h��u	IЧ4V�:J�$�̴�;3��������L�7%J�IUZ@}�ڔ��}��������@�箻��Ƶd����e4�����RCK@�K:'x����r����v�U2<��s���i��#�	�������Kn1�<���{y���I����@E����eՙ�:l��a�w��gM�'���dp��/�^8ť?����][�bŒ��H�wo�N� ����m�Z�`#[���2�Q�2��Wⶎ�{:ԝUt����2���"/����#�1�s&�����(.��}hm�Y�/��e��?5��ᣵ�	$t��U�3���\z����¡�$�z�/Y�dddd���NWm�޽��?��^�������;s��&�`����Wk��:�Vy���Rm�u��P�P�QG���@ �����������s�}rs^ۏ~^�4����9�?~����9�h��}�i����5k���0g�}�ܣ�X��1���޾M�6��@�I�ֆO����s����a������o��wg��l͘��PBh�9'K�kQ��PDؘ?L�h�ƍ2�m5�Xx#�����2�(9�i����='��;�c�y৿��-ς:{{�C,��
�X=C��؊Է/�4�#���q�l��@�4�G�Z�6cFDx�J�}:V�:�O�p�B
��@#��)��~�A�a!R\�k���CIKL(y$��#T��AO%�x�kz!"Cr8'�|	�'�9�3�̟4*��'���6*3#.-%@��"7Ml��%�je��B���	��
������Ѝ�<&����G�(X���K���DJ�'�+b9M���������%뽇Oru:Kݘ(�:@ް\�+D^|0v(����xG�oa�&�0)j=��j�Qt��EC��N����T�Bât�g����#���,��j�Z���r"3� >.��E	�Ғf�t�i)��T�����MVߗuj�'`HU���l�Bp�زԬ@t�1�+:9�C9^�^� �`�l�]à��K&r�+X�	��85�hLtiQ/���_��g�>��W\��ѧ��0z�g>���$��tE��#-Ź9 F��u@&)r����\%��ぎ�5K����7�MX9C2��"S��������caz_��HRԇ���O^��I,���E~E�	��T@$`;��B	���D��5��_�O0:�H���3��k"X�	��r��.�ჿy�?�Z�d1�mBxw�����"���>9Z�9���1:Xlm�������;��ݷ\}5f#1h��6���0���h&g�sv{��Fvgӊ�Oj�J����2S�P�0V"�R�	�77���7�>�m�m�F��� ���Fq���9�X68����9%�d#����-*V�Q~�hii���\O��TWy33=��F��bZJ�8S>��۠��ULTŤu"a���͞s�K�
	����(T���j�rF*�WK�U�G�qDߚ�1���F�7���j��Q}`�G>��ˢ\FG%&�T�abH/�|.K@�Y�|Aj�Z����2�M&2�D���j����Gn:$������\Βі�x�,�eT�AahFGǹ^����1�֨SM�^���e0G���
Vz[[U��\2�c+Z�i� X{�,�L�D/�0Ű>@߶�Kq��0D�vn�ߟ�?�'ZJ�u[~���>G7�^p�iӦ�Af�K�3�`�����3�u�Q��e���S"A�-'D�u���PN��D�@��ڤ��4�Q�ULp���8��GX��pO<VW��4�S�d$��Q)����ԯ |��͗���;^�P���k��w�ȳ����w����Z:[�f�ѱ�럂IBt�+N;[��bQP�SnJ�7�h�'!�x��<�����TDF�/�i �D�r;|F��@b��<�=U(����w%�GG������^����*Y�2���uV'�z��	�#a�ɣ˼���I��zTTz_�B��r�P�C<<>>cΜs/���͛���u�<�H[���v�S����]�n������^�?�О={����zꩾ~���a������������V�#Ǟ��8w���6/X�hƊ%[�l���x��3��F��ӥ����RM��>�:j��c��aLY��M'�ނ`a$\iR���Ο/Q�P��+���ݵk�����Bqh����V�`�*�����=���g_��W�P��29��|�d��?دڦ��c�1E吴Z��ഌ7BПn�W��+4��[���w_z�B�m�g�� +�W;>>��7�?���S^�x�Qϭ������l~z�8y��>�J�H�a�:V��`���$���.��Z:��)( �T >�-�2J���"�A���q���!�Ja>��f׺�5�r�� >�F1���P'%�����^`��/&�B0�8�u��4̵X`���+-j���
vxz��1�������ɪ'��8/"o��2^��2���ՇȰ��\�}$.cf;���9VŴ�ϟ�d�3��<h�^k_C�]��I�x~��*«`���b�Ë����x���$�nu�X�Ҋ@������-�� #� ���A=4,��f� �t�`�U!�X��
�)�FyuD�q�s*=`qU�c	\5�+�L��� �1�M5
��0���Y��Z/q�i(l9-H����ı�@��Ѹ��oߎ|8������)��R.kw�q�%�\�v��֎$J�%��;����b�#ߺqƳ�-RF�;<�J(sʘf5�o�%ox�{���Ɔ]�T�OĐ�r�_���^{��7�t�M.���K�X�p�t��m���.�:��Ķ�f!�:�q���v4�-8�L�v�f���W_��[���[n9��N>�D��[u� �ǲzv��
�»��nPu�6����G>�����o�Ϋ��ʣ
.pl���L���=>�?������p9�@ғ�1���rmʴ�,��y0v�P��Y�/�6�K:��~����@����y-)H���
t����3�"f$��2��G����e����5�ȍ����k� FFF���e#%�l|k��>'3���`J�LA�p#�c��r�ʓ
�Pw����ߏy<�yE�΍����-Fˎ�tB>V<�I��&�����g�R{N�L/��Cy	����B�P!�vKX��MQv�F���z�k6>���Pb
��(��o.�'�`��i��U2#��[�Q��5�ᤓNϪV������>N��6��b�^x½{�Λ=�R�e�b�4w�\�Xڴi�s�y1�� !21� �b�T�܀���P��'��z��zc�!��=3E7���6�D�RF�|�%!��b)��'�^o����ɃE\�H3�d��kk���\�K"�)���2#Fr5&
2�,
�c]G�Y8���9��d��@$�^A�����&9�=�~2�i�Vfx�9���Y�(@M3��ԥ��K=�Ϛ�?ƽ|��8q�}��^ҹ�4Y�A#B4�)�|���Y�]ϓ�̙�a�z�~����;�lz{��p�Z��j�gφ����!3s�̭�o��,]��442���O��a��~�I����g��G̚��f�`~����޻|�r�h#�qn�u�>sB��l����BM)c�L�c���y����Z[[_x�y�\����HX�O�`�J��&D{{'��$	�6��j���^��1ŗ`���ƅ�>���۱�\v]��36��] �~��{N>���ӧ#e\�>�7���'SMAZ�#f͚��l�2������j^���TSN��)f��9zS�&��x�cO4�����*�)�z_��ڎ�S��m��.��T���=�6�P�=ϰ,�F쥂i�`�5�j�9�K
�m����
�Hו�[u�-�(cӈ�-���,�
�@���a"t���e��	�WR-IȣĖ��oˆ��%�6��fx��g���Y�7�r!�5�Ox�|k�zհ���8���ב���������'��)p=�a���/9B�Y�bPk���Y�Ҕ��Q�6
�����m��,&���`�}�$H_幦�[
'�]"�91x`���a�4$ތ��c�Ⱥ�s����9^�^�LKR�Ví�X�b�̕<��S�ŭ��l���ʕ+�Z�^G�<�#�x�;���ܵ�����>r��s���-�b�5���V ��|��R���P�)��@�u��>UdL�9t�D[�w#=w�psDS����	�� V�
�o���}��S�zϻ���/��c�=&LJ�G���E˗��0U�By?�L)�c�B.y�0lv��6<�1i����E]2ES^RD	6�����w�kN�������~��A��>��/YVK���[;�'%�}��ۿ�_��׿y�Uo��l9(y#�e��D�l|�9Ö,����ڱ�]�Pt��0wZ�F�"����',���1^-H��t�� ykG6�{X`�^R�#�
U����L/�=b�q��ha&�lH�m|/���U�Q��L��t	
��M��M�[e4����C��9s烍���v��9�i��׫�pMP�A�8���.axX��&BQ7�����H_O�2�.L�ze(pU�^u�~�f������sdN�R����'��F(i�[���\�ƽ:�5A�Y\ÓF��LL�ZH�,3#�j��	@��]�Y��TA���$�D�P�`�Q8:�}:�~�M��d�<�d��n����j��\�I��64�:vD���,T��rl��^=���{pp�:�8k����p�M��� �,��|�.�|�+��n7���#�_�riW��_?�n���ј��e>2��uv{��#�;w���X��F]Ռr��~�Vii+#q�����a�ƘYFw�_�����B l8��VD�Ш�mG¸��0��bgH��) ��xT��&����}��L�i4����9a�������;6��a�+NYY"*����ǅW(��BS�k6ج���H�FH�Ԣ������m��:哧��z�,eYA`�R���#�P��'/�).�� �?s�H3�h�K��w����A�	׫٩�=5���>0oJ�p�tx�ꉲ[LkC�#��-��z�S(u͚}�므a߸q��j�c�Y�j���#�-���;���M[Ǝ�j.���ֶR[k���wE!�'������۶m�������=cV�.yU���:��}�%��!�����
7E�!����h���F#�KAa�p�G�� [҆c 𻤏��*:x�%���>5�ju?
�j�,�Ƴ�By u
E��]�hN�2b퉄��`���P�&�d�@�]U��i3jn�u���:"Q�"�?14[W]��텊_)ťP4@� <L�*�K�J�6���u���9����o)Zߋ{��ӹ�Rk�ͨ��T��k{�*����,�����FK����E��a7�8H&S�h(i��8
�?��J��k2j� M�A>^�#z�G$�rШV�����Aa%A�񻲃�(&ƹ�!�-���H�Z��RC���{��&�Z�m�V��{�iu�q��o揕}0�DW�ܔ�r�Z�jD���o!yk쿱��4�KxBi]q��O�U�Ғ�2x62T�c�m�q#v��Y��W��So�����h��=��d�a�iq��^�	��v��QQ�2��ZB�hU*�8B�`<u��G�#�T@\k��	��el�4[�DHL�po��c1>C#��q�*N�E��!�Zb;�2y�a-��������Db�ˌ�'�+���/}�g?���o�f: �A7_{�R������.���~ ^��]/�|��T��P�P�4"� ��@��3'��x��a'ި����p�Ȏ$�˿�$j�T*�by����e�ɯy��~���'�ٰa�H����Jc&*���~�S��9H>��=:�R��tR�S��TP;�|���X�\>���~��y��>�`���n0,�Z����>�	g��㡡[n��u�7��ף]��������^lmm-�G�22��1�p�����&#o�039��gQ�U���u�|I�-�v5&�(�H���wk����
#L�hB��.,!�w��!��i�IFSƈ�ZF��)�8b[���'����a��G�fq��Սz�~�z�.`�Яp��Pel=����C]�9s�ҥK-Z�ïutt��������[�A��+np����V0I+�$IRr]�,����ɍ���Ӓ׃MZ����|B��u���?��S��Y���"�m�j5N2c�H����w��)K�0�Y�lNTr^4ʲ�l���������ޱ����7{�w-^��U'���<�*4od{��|ъ1,f��:;;�-;�'���p]�jU������䔦ŉq�8⽆���b�[��U� �VS&��ɗ��!��������t�д�=Y��ĥ��k�ҿNur���n����V��:^b�	ٿr]{�5��Y�J-��ζvX��>ZrӦMCo�q�$@~<9���ה2D��Or��Д�mj�e�L�ʤ3����ȋ*�SA.�;����.(��)��>G�L�-�%�������ϡz��Q�C��s�=s���)�������q��k׎�����̙��oq���ٳg��,�`���]�v��:o޴�N;m�%�=����lٶm�]�����P�,��CO��MC�	Hk+�$Y*:L��j�T-��R[���y�?�_jQf̘a�1W íyKrS��Rٖܴ䃁u� ��x��+t�\5����>�Q�QX�j�v:���ʞ�;v�5mɒ%U�ںu�8���k�y���n7x`.��3���7���zô��
F~���o]~���F�o����]^��h����^��K/���ZPmIx����\��##Ƥ����(�w���?�%{���X\z�������X%a�8Nu̪�H#�y��⣏��k�L��3K1M֒%K��݋Uú�|�q�<�H��T�H2!��N�B��W�h)T�����\�p���]�W����Yw9)�f�֥�o���3%%�y�E��pI�	I��|�o��}���Б
]���v���6����З���o|燯��u�?�)5U�����ۿ}�O˶�)R�3��>��_�u�/�����w���nx_C5.{����ȋ��'f�i';w�<�5�c�����x��v��!f8�ړ�=�s��_�����c���VMy��k���͖�#�M�=�y��o��Mo���o�@��>��KV}��>$ɮ�����F�ʣ_5��{��:��q�)���Q��-�B&uA!�$>�}Y:s}���?��=�Lȶ��3���؅����~.��$�ưs.x�Z��S�Xd�5О�t��[yv�3'�t2XH!���X}����O|A�p�0(�V#�l�"	5��BE��H�IU��"x��,�q(b�)�#�M�z����c���/��g�>���λ���H��ls����w�)����pG�A�"K�Z
J�@]X�bI5�e\����C=�� t"�K٩*�h�*��4D�(�)'ʪ��'�Z��
n�U,�U�P���v+h{f�Q�0��"U$�i��@u����-�(s�;5���������#���=c�O��Ǵ,Pm���z�� Xg-�ߨ>�뇦w;��z��J�T���֊���.�[��B��p��C|a�z5�n�H,�Pl4#�Ŵ� ���� +�f������SH5u��,S����2nQ�0c�M��o$gN�Bl����[��P�;رm�y����"��@cA�U�C�2����[��yl�l$�؃Y54���]%���m��r��^ކXq��ā%q?75yk��D7\Ŵ��6���7�r��D��fbԠӋ��,���=����s۶l\�r�qǟ���Ϗ�{qwL�@�؎��Jm�G/[:82
ׁ�	�c�2>
ۭ�Jp PQY��(�`�Q���Tj�R��[��x7��d�:K�"Ō$!��L�q��3�`������C��:��Ր{��+J�c���KW��ׇ�R�T�����"G,Z�o���r������KX�)�K"��"�7[���#�?(�z�n�o���i�� �"9�tw�kJU�ϜIφ���Ϳ����٣��>!}hJ2}�����v����3�l`�6ps٪ٿ�w���Ni��彽���������{���կ@���78�ۻ��%�l��Iͭ�9���g��Rp�������۷;����5����������:J�׬\啕o��W�w�*��Y-����=D�t��e���zN�#��u��Y>F��N�:[��c:J�����0�����k�:8HŢ1w�LM�c�z�`��O����?>�Z.8�V�{y�m��e`�>���FÏ������؜s�Κ=�lYdL�ՙ3��7k<���ɐѥ`d�/���,˯V��OfX�pw�����-H����%��iX+�<�Ƥ�R�W��"ǿ��N=�L)�T-�\N�Ԣ��5Wþ���h�T�q��4�)�b�tb��2��e��#~��ǎ;��R*�UU3dEsC� �
�r�׿��ދ{\�ƫ�f ��}��1���ԧ>����QH�1�Ba)�������==}p�'T	�(���G�-[������8b��MOuwt���-?1��
)X��	��Ռ���h�r��Ġ���'GtpU|F�ca�s׀���h�XGTs�,#�'�Ǳ
~���6B���{D15�ֳ�)���<:���E���ju�ҥ>x�'���7_�/���];����M�Qm�#�Ԗ�'7n~vǮկ^Y��"�K;�A���_���K��{��vu��R�h�!E�J����xn�-�nא�DMڈ�������m�C����E��y��k�đ�,�ҋ#-��Kx৴yħ?{�&��Z�t �5/��t�E}񋷮Y���s���0��[�L�5f�3?��d�����z��3�H^N��S\���i��K=+JI�M�)��
�E���91�a|۲�;�807�(2@:J�nQ^+"os��z��W_s����l ����� �DWPh�.�FTRy(�>���~��ρ���qa����M̈́qY�fM=�Ţ��2��[�C���B�|��$k�QKeLAHSa����I�l繄ɮ� �h��і%.Z��j5�Ѕ	��üWb,�k���5���5K��|eH4���۔`71�@%(Ǳh�k�F�B�����_|<���:
�x�}���[ZZf͚����Q���J���g|��(k�cǎ���:vL���\�d�u�eI:�Ǥ�T�/��n�ӧ�=i�9qi"� 5�a�Of,;���3|}F�#�ݐ�(���zR���5+���~_���F������Ƴo�� ��J�|#eAJ�"�!G/�s�9�uWxv�����kWpx�=O?�t}����z�X��&���DH/�Md�6�QKK����ܹs������=�H����vȗ�=�9p�ɍ�|Ф�s3[I�Wx,�I<ʜ�m�����=�����w�2+rX�����?*&�1є���H͓1l�3�0 �J�sw͏~���L�\�x1�60JL9"#�}�CNi��W����yiq�-9�Q�������ىI;x�BL��z����`� +� �8�a<��3s��Y�|�ʕ+᛿�����Z�z��iv�Z::Z�[,�`�E�u�Y�ٸnݺ9�f�}�٭��g�\~|�N@�mM���n��6*��Ղu���
R�߿�p_��Lӕ��ӄ:��rf=J�J��:\�$cM���*�
,�}�l@�nz�9�SHw-�w"�>o���--��<�k�������H�g:�����k��\z��rD�s5���~GGxY��̓�����`�Mq���wK�Uad�!��J��/�}�����Mz�o���G9��S�་���ҥ(�h�	ǯ��9���~�a�A8?�U$��������1��
����x뭷�|��?���y�+��UA�n���_^w=��^z�]?�6vP��?����r�g��V�Xq����p���\�������e�q~I��G����u���؇?��BAo������k׮}�����]�X&���MY��L�D�L��.`��l��k�N���qZ�2��r#���G�q�s��Fq�j�%�\���Դ,�=4x��o���_�aW�󑿻�K_���>��{��дi-w�ul���N4�L�u������k�x�]/���1G/��J�y�6m���?~ڌ�HK�,�-��_���+��=I�*M����a�"��9���ѭ�G`�}��v�rl�-_l���?8X�ȸ�	ô���ߛb�������։�.XU�9���>���_D�`7�*4d�#��g�jV�'5�KY]����fH )���,I=�O���wg��n��8����Ҳ���X�L�
��TFKq�L�J`��Q��.u9����Դ
�d�y��Cr�KZu�}2�S�I��z�K���=]��)&u��C�z ��9���
�;Q��XU8�(LKÓ��\�&%�AT6āT�BB>��d�䫡�W,tQ��h!��	�Ը�wS{9�#Yձ�)%4���j��T�$�g��$�Z���U��h�1��hzZGWW�����\-@�/�ڒ�'c{�,Ő��s�Ah���H!:3���%!���vp�e̍��	��n�Ɍ��Il�F��7����yP��p	!RI�*r�s�ǐt��� "d��d�"�/K$ʝbEP�c���L��,4ΙHR�dP��DW5r�#�&�zJ��$����)�^aÐښ1GD��P½�T�X#GO�Pc?N�O��l�c���S
�@ʅ"r��rq��"ɜb�-2��c��K�Xk�{I~E��̡&LLʀ�}PX�+G��;�j���)f-\P�>44�_G��ys�-%gG�w��[��ku�~���^4�3P��,����b��#���n�F*�N���ZM�L�"���9�Fp�c�"Cr�-�S!�?4׌��'��J�z�o�M��f�6rQ���	4�CЮM~�N���k���c@V��-F!�%��Ġ�kx���`r���Ukԑ�5�<��0I>�|��D[*�B�# ��qi��<��x!$��������,sE�bL�:��DzA�4_�1ɿ��1&�,D����W>�9��U�r[��؄)�f�jR�ڰ)�>{J M�{���FOchv�.d�y�����[ox��Eر��e�&5�vuy�c0#�{{�{��vN�)=�o���p,�:����n���i]��o�e�T����q�cҎP�+
�%�u�]����ӓDB750ruE# �z��I�v�M��S��h$2a"$�Yix�����ٰ�ڜ��7v	m�S$W��#ؓ�?�۫���\*��8�k#�8���j���H�-f{;2��lO�c�u���@��]}�m9��Ah��N&0ldZc
V��qV�.��J"а�΃�����\���3_���\�&�(�5uޜ���W_}�O��3�n<���X�f�Txa0eW��{��>��-�>��_=\�6̶ؠcl&\��J����JM���u'��D�2�`�П��?����>�S����<�@*�7�u����3�ud�O��6Ru�R�6M��۶�\��ď|����*��wn_�p�~�H�"�h=���TI%d)�����AI���r��ʛ-�b�\�N��HRJ�{'�}q�~FR�}we�L^[V�K�"h-"g6$����8�Sa��@a1�$�0����ӻvo{����;��իO���;ç��I۶�2d��o~�?���~���_y^��������/\�t�D����%ҕ�^�������|ӕ2ldyo��yz���#C��O|��_����KiS����?��W���5���~��B���8��@�Y��?`��O�x��z��h�}��t�(2׎�G! �6�,�(5�KY`/+�9+(ߴ|���0/C^�%"1$�dN��8�X͋����|�����A�2/FK��1��cH�ifʤ1~���%B9	��}X�Nx$`m#N�e��!��g#��O}xx�W�8���ٳ�.[D�U�X�0˥r+���G�8v�+�4&�a��3�X,ej������d���� &�-X)p�r�ο���FFF�<�uӦM�b̜9sWw/cb�xf����(�������p��MK���4�P�,bH[~EV� ��;Gs�8`rV7cgAN�P�1��Ȱ�a�8�:Ɔ)Mӥ�BYR1�$�D��C��>��<��%��b���F	e�'��30�]��>��Fف��������q
��#'�x�㽨��|I��:��4e��G��3�l۶���{�*��ٱ��U+W�����Ҳ|��R����|�u�|���]	�������;>2�W޵k��3f� _cd|�3rv�R�8G'0o�غJ�ݒou�ߚ���vM�M���/�Ҝ˼��>�t��B��+|8l̞<{��	�RV#CkbQh��j<�G�dpa�af{&=v��������j��7uF�p�J.o�,9��เ���>k�8�������8��X���mw�y'�VXޖa�=��S[?�I�|������Q�i�w�x���z=Q����v��kkh`�<��7��Ѡg�O����G�5�]FO<�}M	j��0����i�-�Q�*:��Hd�����wɅ�Z���X ]wnߍ�s�GLY�g�qꚓ-Z�1��_�v�֭[S�Z������������gpp^��Nx�;�	r`���Y�a4J���c��=�a��]{z�9Y�T�F8�a��O|뺌����VC�y�|�bw��Qz�U$H����?ܱc�'n��5�\#E=o ��1-�����v��X�BQ\)�EȢ�V�,,ۮ�1||-��rpW�`'���m����ԧ>��W�Jj5���z������������'?��8Bp�/|������m>���>��M���\�b2QJ�X��R��տx`s�Z��*����z�w�	���������ɍ��0��L�a�$`tM�tQ�Κ5Kd)��K��ף�>����v:���w߲e�@��Y�f��툹](I�߻w������_�*� %%0N;����w#��Z�(*��?��
��3τI� �d�&k	A/��-o9��^t�ՠ���U��xi8P֦|!���?O�_�9&�Ac�E<��a'>��-2��`�V�����8�B�PZV�"���Y�m�8p��!�x�_�Z:K|�u�� ,HLN�.�i�}(2��3NG����Z:*�})C�{�
1*0��2�y��s�1��F�)�8�d�XB�;#a�)�g�	gCC6C̹��C�M0�j:�\aO��/�L�s�ϊ�B��U2�WlL���%��+r�!�kz$ɮ$M�\������7,���ݑ#$��J"��H�C���+��2BN�]�C��##C��0A2�5���b��hs�6C�|#��<\=T�nv���w���sgM���^�:�m8IHN�&!ؤ��0�Le�{)�f{t?��$Tp,�1����5�h*y�e[�jaÌ�1k�5���M����
+F\����;!J�q9�gV��Of�RI��
�%	o �
Zפn"�OŒ��<Z�ӭS͘/B��6X�=3E��-A��P3��GE`���az��E��*��6�	c��3�3x́�!��B��8��I,M�a�� ݧiӦ�f7�PT�0���5w�\i�W���T[d��j�f�B�� ���pM�M�����w��9�fk����2���d��°��Q.뉒l��L�=�.���-��ģ�H�}(�K"��BR�B6��1�T3��Ԟ���Ll�� �(�$�U��#L%��΂[���"XҰlt�T0㪛�}=���.^;�|����$H�)�v�lj��-&g䄘�:�s�3MWRf�%9��T�ȡ�k�.����R��M�K☯P)����R\��彠�K���SR:�\J��q�M������j�I�G1)m�F,�(����Uj����:U��q���_���uE��-b^]��hwo�Z-UC�"N�Y��F~u"=H�C�~H�M����|%�R��i�F�,� ���b�|����N,��p���^��˖/:�5k�\��Y���{o��p�A�;,���e�ܠ`b/��������[0μy̏�
2F�裺^u�ʥ��Θ�'�ф��p��a�*c0�,���G��l��%Sg$��8K��슦E01�S�����'�)���偧ju(.���K1����_?�3���@�k�`K�rRZ�l�M����1�р���c�ןް���ώ�j��(�b9 ��0U��իM]ߴi3��A�%w�}/���I��X�S�vS��r)IBC��<�6���m��E I#������f�#O6澮t�M'˙����JJ�/ExQ�F�b�/S�	�[�qO��F�|L�/��/��{��5���{g��~�����t�|���������UǯJ"�]_��Ӧ�4l%���A,�K�^x������~}��^g�؅����޳�?���3LӮ�p��W������{{_��O~�� �Q���C�����/�d��8^�^����$i�*�Y͉
�����w�+��
��`���N/y�WXCp���9�܍
:��Q5����&!r�)���x�I��,m�o<Ip���\�sn��|&���`M5E	�V�\l��32�"�z9/�:::|j$�!a�LBhK��,]�t�.���;w���IHh�h0>>ڪ\.S�h84�����f¤���J��N,�b�6���˖-S��m�@����"�h�1g�w/\�REF2�)����ݽ���{�Jm\��� �֨�)WfHX"� ?����x���1�n���!��&�f�W=�%d�t�dlt�����*��`i�����yl0��a͏��z|���288��ъM��C�_�<�z�I-�۔	ˡ"��kD�Y���+���3�)�S�C��\T�'y54�3�f2��A���C&�a������u.��^+Sl������/\s�[W�XqªU�j�֭[�y�񑑑�v	!zq/����>�聾Aƶ2�Y��,^��w�ĭ{hc��M��b,������������t$�#�N2��D8��P���L��y�DNc��a��B��?�����y��TW����N崡{#���;]Bm�ZL!�P]��עڡ�~��ҥ� ��k��)5G�'�I�+���˓�c<_k�#��<sul�;��Vp�W�-b� �9�����|��9��
�=��
nÎ�6�:e�� ����(�Z�[$����a6�|!id�\	wZR̕]0�v� KN������̀p���)��s�^�η��ڱcHo!E��::[�̙����u�����ƍ��Xż:G��"��h5�سgϯ~��U'�x�W:�U���
f꺦�#)��m|������k׎�������,�T�5�����Z�[����DѲr�w��X�`�#���C
aw��|��k؅"�a�,��Nl\V���۵k�����Ó�H��+_m����/vQ�R�9i
1!�:P/��B�8Z�ca�^�+�%�"jIJ���]o�U�v"	�ww���{���_��jJI��#M�o�G�Ⱜ��:҂���(pDp��Q�Z��g��>p�=�\q�`�Hr +�SO=�;V����G!Q_\�g?��1�cZ�������.��B����#"�y�Wlo��;.��B�*�=�g���7_��3��L��j�$/�����������,�>"a�F�n���\���������W�Z$��BN
(G��b��Oa>��!_2~KP�7���I�R�=A����r�����p��Eդ8�ADz4��"j�����/��tG�9��nI\�Ο�O���K8��vn$i���KS�J���C�:��Ɇ��I-��TӒ��a�N��2fT
e'��B�I��~�b�l�P>j!��X7���$`�z~=�U]S|o`R{��!��g11�x
��-݁���fZ�[CfՖP��_^_�(�N�1����5���q�Ģe�hr�K�M��F8G�m٭�TrME�]_�E�n��|T6^wt �&,"!�sl�r�����	�1E]MS�$&�z�E��A��T]I`&X�.�<��	S�&����|31�����=*{�V���Q���ZT���x��lF�U�ԙ���D����������Tؚ*��*���uag��೩R�K7D~����/<"�����E~�����!B̬�|��Z��:�,�U;���X��:�wT��b �	>G� <pB,�I���%���ah��6��e*�e4j���q�0�|���z�޳iK���s�t�f��-۷����{�tׇW�E�疢���#�k�?���C�^�lgq6ott�"��Z��v5�pC[
k�#	 E�̥+5���]�sY�p���R�q(=���\���~�ON׿���y�}?�b�x(S��N15��^�����1�0GA�K���fR�r	gT�75�p�SU��lMRH� C�p1Ǹ�m��U2�L^S} ��y����:��*��8�Y��S(nb�YW@�[��F0.����X)�eX	��h"�4-H�8c�Kܭ�	��c5u<Vk5��T���b]K$Z��
�?"�{��b&{J��a�ȇDN�	 e�q�\SJ��$�rD���R�@ǒB����´-P�C��ma׌3�b����6m����k�{�@Z>��V�ME�ji��'<>t1V����0�8N!��������O?}��GKq���IŊ%����ܻ�o``ԭ���g&�^m�:F�����<�b-:�h��"��M8%�ECx*��?�F����@Ռ���M�6�\��)� �"rJLE��7o{����X�ѷп����ѝ���	�ߛ���q�ڸ�MW�0��c�P(h�F���h�3R;�O>�h�"Ԟ�d�(� ˅��恋�?�~�_^�w�E�τ�4+:&�М���T5S�����4�n�͏>��_^��O����_���$'X�U"X(��/���������_y������
� ��d�`�\����"D)c���-�P(���++!���S֜����F�>�@{{몿8G�9'���V��互*��B�Ȣ�KZ;Jq2�3j�y�A�v��G}�QC�k��ݻ�����:���@T�_�qT?�ۏ~rɲ�^tIc߻�8��>�o&�G�&�g(gQ���J�?��_�0�4+��"�/}i�Z����r�a<IE\Dȉ7��g��-R�_F-�aN�]I�5E�/�������N?	���S$٭�9:������iy��a�xIH��ǹp�S(`�/\�p������_$[�l���;��̖�͛7���/�c���GIkk�B+��m%l|RcyÆ�Q�4j5�:؋��� Ί��b�3}�������дi��:^��hZ����n)�৹cc�```�u�>:Z�|d~�4΀��9sfͭ�d��e˖���]���>�����bxL���J�����CC���/^�ګ.�����p_/O?���]�sul�w��]��x��^p��g�	 |��;�\�~=��g�}68	���U����O/u�炥�6�;v�����'�ϬY�f���`�����?�!������8FCM��a����*޺u�F*��Ŗ ƌ��t�j�F`2)�_��)>/8x���d8J�]�!��81�	��"���f^-B�(��?Sf�B̉�q����]]]�.L�v�]w!�d��4����vX��s����vɁ��9����]{�/<���7��%�A����?�h��)T���=k֬��:jdddמamp��4�a[�o���k�<:�d�'������P�&�g�7��I''<5Z�L�AL�����-7e�4���Ȭ�0ZdAx	S�7N��/��4�4J�/�҄�|~�Ҳ�<���\Wšq�C�M��*A�%�i2����J�bc���
RbŊ��Ӑ�JQz�!n�`�/��3��́[S�K�r^���2�ԙ�^Eat����q�5�����`�;���p�g�}d�����<<���"�k_7��ݥ2� 1(9ń0r�!��F��nA����#d �M��ߑ����̞u��G�md�s�mI�L偣��(�������T�6��`���૷��� ���;N:餟��� ^@bk)/D
ƫ#�j���	�װup*�z� Xn��+�,o�hY�
L����TS6��s�1�#��뺁c&e�4��Ib��s�0�0�0~ ���%��az�68�$�����8��;��^����o�Ýױ4�B�?a<�,T��u�^�5���s�=�?�d2�|�4�c�=V*XaO���ꫯ���`Q{�1O<���ٳ1�*���k����
�ndh���~V$�
�5ػ`���/����;w�\�j��X�ڵkY�o�֓�Dz�������{��XorK-wwk�%����TïH4��?y��k��ф��OQ
�j3|�c�ϐo��h��9fW%hp�DM[��`H�r:K4�d�_����������Y�Elhh�a�*�I��Z�c	��[䘑��[�Z�][������g�־s��D�٬S�OE�%�0��q߉<���.�Ff�T�o�m�^�>OS�PM�^zp"�E[^Ew�K�X��/�8H�֮�rg��Z��wð满Ĥ3}挽=݅�2�t�E�n+�u�,c�Q� +#�J�:2�`8��� B��p+q����1��m�}΂�y�ʝQ�*:����Ì��j�|/B9	p:�׃�����$��̂��H=��0gUl}C�W��qI}��U-�G��2�c��<����.����Zl�FW�>�ôu��T�;�';zj�P
%����SHl�s�����?t����oWJe��#��̑9���7^v͙5�����π�^��h��e,SɊf�'av��R�!��`�~��ЛB����fd-��'��-�y�"�`�S� �5F��
�d�3��3ڈ��g��y� �>IDA�`��Ķ�R͌$��sk-����dŇoZ�T�%�=.�$ʱ�8q����������%B0ө�'2��TPѰ�1��He���w��K`p0��ͤ`k^�`���o�he����#��HD�L�m�Ň��$��:ȝ��4��v���zt����D�z� K�2ڋX�a�{v�c~�P1�8�c�`�*0�hL(�~��	�b���n;���@ﴯ�������TrR��\�@�Q��Z��C9�T	E+c�kŤ�\�GA�N2�0p-S�J�;������Q`�rl���K-�z;`�JJ��`�*ըXw\Y���ƭ���!��E�6,5J�����۰*jV�!~�vuiŌ�a��ql��J2�tl�I���H�~��H� �Vu�'IO�PkkkË���!���h?�Zac.�*��tu��& ��n�'CU�0�t� �%�:r=U�F4>>Vsk~��6xY�C�F�"/���Ux���,/�tJ��5`у�V�T��� g\I�NU�]���T�jkبΙ�D��=����&�z�Uo�[ހ)'I���5���\Dk��K/��w�x��Ws��b-�n��(�|�9G�s�i�)��~��'�?�̖g�<�d?j�WS��������'�X�1�er�^��nq�Kr�I0���e$�"�M�m����w��c���~R��,���1�J%�����?�c�K&HY��]CS�j��o��/��` 5Uj	ډ^8��=HL�ϛ��m�_li����>�8��A�&��/Yd$b��g��e��#�/��T�X�J,c�?̔.���0�{��h��Wm|~���?~�Ձb�v۰�Wdo��o��������S�=]�!xV�	
KLKs}��5���� ��?��_�eJZ͒��L�y�30���5��P9䖃���" eHb�h�����P�`w*y���Y��~돲/�h-���c�d��y�	������kB���X�)@Y��o��<(>gΜr��Z�#�<2R�H���*�`�Θ1c۶m	����,(��2������רx���*^S�D�x#rm�P O��*R����-��|EN����hi)R?�����7>�FdPk�W�$I`�Ç�L�Jj2~;�(�u(L�u.h���E	Uˠb?߅'?�-Z�Kr���4�S��Y.ϝ;�1
��`��::;�O`!���x��e˖�����׼�5��{�vð��J�#�nXg�����G��'"  ��IDAT	6��r��k�%dqI	�p(��4SlT��(��L�FN<�ƒ��>ƃ#���`�h!H�督t<D���>x�R�R:8���.�:lp���#��/�:����q�\� �bz�w�_��`�f͚�h��p|Q���v��744��5�626��/�����֬9��R`��,p���rdw�����~d�h
�C�.G�Y��r��T�w�p�?8��=o0>`���\�|9�DX�02��C��u�)�j�#�w������p|�'��Ĝ��6��ݡf17��������q��u�:7[²�Vȭ:�f�S�~�u�,u��]�<�;v��:,lU$9�$�T��Dq�4|w���ȁ�I8��V�z`���"Ѹ�L��%�ikG�I�F��w�?W����5�:���Hd�"�,r&����)p.(�9��5@���`^�����񨣣�QnEyC^�����ZB��12d&$�1m&��sR\C��#Sah��1���~���7-�6'�Re�r�����8\)�����&Q3~/ݐ�1�؏yv8U�q��;�{�{��_}��)�?d�����ǀA���084������P�xdl��,3�Q(e-���z�X��?�O�t���w��p��`�;��T.�Ĉ��H������_�W�N�w1�il.����㘠�El��ՠ��y�nq<묳~�!E�'�#�裏n�}��)����q2�J��RRWW|���{�_��u�{��%�Yo�����|��O�()�i����b������wm{~��Y����բp���V����V-AG�&��F�9M	1��LF�!�B{aP���`����_��Or	}�W�bdT�"�Ґ"!����c�B6�P���B�k��C�>��=�,�����m�<7�%JF~ʿJ��ʿ�%,Gr�K'�&����[���lI�1U�<�*zF������D�� ג܊�W�U�	)"���Bū�ȪVmp�!������)4D�8 �B!����/�7�|aUuy�|5V�BtәHP$&�I�Q	�[�����qD��R#�Ó86�W��Q�a:.U��#2&�R��o��]�-��Mb5m��)��<��H()3�"zUX:��IH%��I�#<�=FM���Y��U�=5:�38����8�xǽ��F�~�ig���|�_�����Va&�p��rP�E;�*L�f�Qs��=�i�I��hb��hmo�EA�0	I �@1��ŶgO��fDI�-�u�(¢�RË=/�T�H���"�^i�ꉁ��66����h� @2aDX�#Puk�r�����W��3���/��`�=��6�N�]9��Ӌ�q�}��j����Rۖ=����zp�#K�.߽{���P��G�:nC�����хu�OȽ����ƿ�^|��#�̮�����K_lԆ������W���X��]+��)Z�W5T+]S�͙}��.�O<�D,�ή�˦u���c��x� ��uBi[�0��mm)w��"8�ڵ�[1����I1sϜ9�}-�8��J5�n`�m��D�`�Lk������ą3��0������&�{���L����*ҷ�4��a���i�e��T<���䚋ɫ�O���3gY��܋/���hokk�֖,Yb��܏����jܳc�PO�̹����Ã�q�XЁ�m$��FĦv��g�;�~-=u��(I���v%%f�)�#e�����:���(j���.풟��<["Q�W�*��y�T,��A-�u�Vy�S�lٲ5�NX�nY�����,]��~��� �D�]�3킀���-fޡ̫��{�B65`QD���q}��=�4�O]a��/S���b��B�Ϡ�-$��P@�~����	Pݤ�I�9=`�K��LV�@ݽx*��KH,4�_�j�Iap� �
 ;;�#3�],��@����n��$��������1M �w�W�I��89)�����)�&\]������@�χ4AM�f���>^���`m��4t�zEAT�mw�B���k�(Q�������~�V���|�R�����0��H�FL�S�8�JW�*�(���t������� Uf�[,�pddd`�
glYG<R���
e��+�
N<F��z@�?!��b\C]N��EcY�@(����� l��`�R���4�d�����x���x�?�V/_u�e�b�;�p*a@%�H4�rX[>U���&�����\)P�Gn졄��q%�3�i\��7}��o��-g�}�)k�~���A�-��������������N�����4�0��:>.N��Q��D%%��#��n�����e���=L��'��a��袂�<�=��zؖ-Þ�S�jd�r��~dw.��db��)�Z���l���ĪJu��h^�>a#�@���G���D�'G�?QX��*�R� �cC��`�h����Z��mUZ��{����^��}���ަ7��E@AE�F��,�h"`���ƛ�(�Fc�ϒ{-(�� �bC��00�І�3o�������*{����1�����?��������Z�d�����a_V�\U20y#����Q��G��F��3�w��Ā�<��]��'�����?�g����}�����������xn]U@'�L���pU��-��E�Gy��tU�����"�'���J->^�X����[hy5�*�vI��n��y�@5ܨT)�if��Sʙ�瘝4x��?[J��sЛR��Ov;7T�`@W���x��v�eJٿ��5�o��0�'�|�F�RR8������.ۨRZM����EZdѢ�D˃h�4yU�~`T����P���$�H���)��#���PR,Km��H��]M�8e���cz!��4&S
�a��eY������#�6B�%a�"#IW���뉔9�[ p f���ϩLL$�h�>���g_v'�dj��8u���<���h}��׾fs�P�>|@;.^���3�����q���;Ӫ0��Ƹ�$ G_B�"a��E&� �Kɚ��Kp@�jo���?a��D?�F�:p0�3AmiiA?(�)D�K�݊�;gT��iN0���ڊ�ރ�?~���4�,��f�ҭT*CCCX�F�p �|>����۽{7@/�fɒ%���{��;�(͟?��o�7n���:8�U��8�m�������V��iӦ�z088臈$��\�bJ�deV���b?�|K8T�A&�y��+ΘlS�VV���0l��և��k��y�jތB	f��c�e�F��5��� q����լ�l���Z9�/u��[���mȤ8##8�W���MOO3!$Φ� �Z[a��}�޺T@��`!L4,�-�c�933��ۘ��Q���\�r$�/�?z�4픣����
G�']�)�»,��3�{qA�¬$� g��-b�g
.N���?^��d�\*�תP(C/�����R9��/��@rн~[����Q��M�1�I|�3�U�wzV���`��ƻ��<u��gSb�7y��vt�Iy��j,am�BA�GDg��>�l!4=�Y*mb�A�	�S}��/J6A�.�M�?4�
& �G�9ڃeZԢ-"sƘ���4:G*��eMO���b Y@)�%���3���c�����6����`��&&&0]c�8��[Տ)�+�F`巷�[��ubM<�i�y6;�o��{�#�¡�o}�ozǥ�^z҆���w_�����j�c/?a���(����r�@��_�N�!x�u�T	Jq��"qq;�IP�0����_�ڳ^��ןw�y�����- �x�u��W����7���с��<Y�(_��Z\�SZ�M��Ɨ����o��.8�˺L����1��8��.ۄ�F~�1R��RW"QB{���~L}߼�h�43��R6�Y���*�j���a�n��M:$n�#fa�O>z?��	)�=��֎䵗�*ۀR�h����_ i�ƍH*�V��y+�׷l�r���??����_�PwE��z=H;2�*9�s`f?���2;���yݲ�AŕW^���_	�C��o���~��߾�]t��ص�����ZA��T9��F�Hݖbf5�� lĜ��Ⱦ��o|ĕ���t(�@+$hԊ�C\�i�s��Q2P#P�*\GS��tļ�4�P^/J���l����JAx_���ɾV�Z"(z�w�*�艥$z�`�0鴘���)S��m�Ų�&����G��@��~��%Y�)��NP*9�ƶ")�OHD���b��,��BJ:We_/ ވ�����O8A��"����*�p����"x��,f�A��/{aP7�H	a��\� � �/�B+��n�t�2�yA��j�
� �)"A�H>��� ��d=DϷ&�H���_��o:���|�h(Dد	�+�P"#u`�bѢ=���S;���� q����mw��%��[�|���s��]�l����ɡ�C��S�r=�Q{��Y�v��Q ٭�Z[K��b5���j��]��oI�J�pʏ�]���S�C�7l}CqP� "j�J�p��"�|K�����Dɜ���Z���$��&����V��3�?�-����-]���K/���/����t������G���7:�b՚H��?��=�]JE�Xİ��OO���byK_�BM=��a�<��� �k��+z�:8p���g�u���zpaL<˶�T�@��`D{�4�{RP�l�J����2>#G�h8�C�Vr�4pgYy�9���x@P<&w8�.	6�j{�S5�e��E�MRtl"'�����AƦ!|м�=6�Z4,�l�iئ�o^���SO����`��sd����%��ų�on\����a�AG:3���4iث�1YN���zww���k�b��������V�\�hɢ���رcbb������G���Z�z���0�\�5����L��`�R$��m��ԦL�c릒�S�y��p<��_�"���� ��fFa)w����K.���!I�f���.5��I ���������3c0|L?�.Y'� *��k@��aĕ�GC4� ��d,n$'�ޣ�SY:��#jg���;�"&.E)yX�M�̢��p�~���Ћg���!>�c�]�IJ�~�`a���Jj(kQ�a���s��QW]�hX�*��
DN���-拋J������sr,L/�O��!)���-mh4��ѡ�J2W�*��P`!�����1��U��N䣔�H5s+v)ԏ� o�Ǯ��4�f��Ue�V��)O�^+[���9�kN.ʺVԘ�=\��%��Y��Wߩ���:R��Q	`�YЩ�7�]P�SM5UDik^ �#�^��<33�N�^��ut�����##����ؿ+-#l;�HM*���e� ��z�y��{���g�~���ϙ�]�9`�T���a��ٿ���t{(�F(01s�f�ܒDbqB�:v\V|-�5��n�����3~����,0��b���uç���CߵLC��E>����yP�\���s���z��c�K�B6]4�$+����~ha��SȎ����Ӓ{?!{Ю G6�v��DF�C� ��|%9
c�^L�w`=d��Ĕ&�2�A��=EU0�/�lE��$��Ҳy���G� z�k1	Ұ�	��ѻ�O@e�����W`���������O_���ky��g�~d��H�kNt3�"�=�g�y�=�ܳb���+W���	��z���$�����tZ�,M��`�
�C�^V�}
�����ZH0�E�<�a9��f��A0L�z5;0$Ͷ��d\sf�9,�<����D!��{� d5�]Ӂ�$��F��+:6.3���YI�)�%kM ��/��2�h�q�Fe�=�-~6�]Y "#_JJA҈o~A�Gꙣ�r�`�>nf��@��I,ak(408(�|�����UW}�`b[$0��}�w\|�E�x���[��ޫ@�c�����7�.���s�=��>_K�k���5�:::x�q�2b�bw�*��\��o~�O�;@���η����հ��H�r��%ߢZ�7l�ph�.�p��O:i�O~�P�=3R�׀=}�߿��H���qæ�~� �#E"�A���pl��ьZ�Q.|)��h�	�-�ˌf�E`�w��}�g(����rfdd�sp>� �	���������,�I1E�@��F����F�K �A�\��+�p�/R��◰ x1�x,�Tm����ڡP��)*R�L8�x�d���o���3���8T�ɂ��w`��ٳgxxxռ�s����ٓS�>�����7a�W�M����.5o�<^�pA�|��/900�R(RhN���K�^���؂������)O<;��#��j��T)
]���P�#ʼ�ny�ժAÜ=�� 8Yӵ�M�k�,�-�	�f���-�䡔���,�cci
��[Ht��!�(°��cLJ���������"/)w��Ʌ��[������ �r�p��a��4�8|�
1�u����W��`������ka��	Ʉ4J��,�f���8X����K���8�%�(���,zF�Q�u��,݂���@tӦM��i8mbxf�����(�T��dk��e�'%iOj%_9��ė��RVy��^�J�RO��u"�u�r��'�V�RK@��{Am��}'I���T��"��boll�}p��U0�����'ۡ��:��`>�該�VR
�Y��`#��c�|AA�F �8���qu%/'�+�X��b�FͳBIe�)�����T��-��Ik,�1l� �b�&SMLjQ-_`MW%�8��	�>W!����3��A��	�l��/��Z]�$�N9����c`j� �]WA��]�����gDxؘ1�N\Ò�H�gwn�;�ct	h	g���ׯ9w�5�|��_i�ݛ������Ҁ�����`JC�ɺ����k׮}�[[��i�4L����PH����<���:�c� =$���=���WjV��ʬ�8%��*D��|���ˬ�#�(���P_j�"��B6;���bg-/	���sA�r�P�(Nlr$X��alP'vJ��@�^x��ߎ�*����̙��j:�|�'��#l��M3�j@��t	g^x�w�}�e�]��@^D08�rKyȚ���̔�JK�1&�!~{���Yǫk�haǆ_�aM;��i��{뭷~�C�%��߯�S�������+$��^���g����~��o����n������J<п��g�4������n����(��`m!UQ�x�y7�t��,'�$;�g)�$�6g�����F)�S��v+�ypW�, ݼ������%�Pn�-�-�$��.��5��d�a�^�
p��A��Q��m{��׽��Icd�.GT�e�K���O?Rڵ��Wj���Śq#�l	Y���dm^׼�{~ݺU�Wg99WP�dH�pUЊi�o�����?��_��I�����z�c������>6dt,���'���#'HQ�v�?g�޽{{����X����_����/\��SO=��ݵ���.\HP	IS�F�����cPt�?�]���ƃ�E��!��JEI���O�x���Ύ���"_W�o�^�|�hY_����[5'h��]c誁B�,]<��f�'s�2��[�\��HϩrA�_4�ъ�k)�����q��h)��o�M����r�<93�/ī7���VN������6�b�F�Jx$6�y��;{�W,;����P�$�T�`55�&�t-
�F�)
�A�G�b�������;q�����O�=7c���N���/.O��_��X]��ޅ}s;��,[n���'�v�s;������׼���������ゕ[�|������膵'�[�v���F����^�|�k?
V��C S`nx`ң����cӊ�kq�9���X�]�J���ݔ�����#����5Q+Wr����k�� M�^�~q�,�x����a�y�H=�%�	���E���^�(S�R���z꧿���6��~�a���í�!�R�i�F-���s6#ٔTބEْ"���`7Y6s�y<�W����a�0ۺ;�?11�:6� �C��ۋl��
�<؁ "���4j�,�t�ɃCC3SӲ�Q���U��]��q*�8[ONآf��_���xڳ;EI�#�(�����<{�)����D�$90�S=3g����9IZ��fA�ϔ��b~���1�/`�S�1�ԋ�F�o�H�AB��&�EI���j<�
�&��5s96G��w1�x�_%�	�wV)d��>_m`~G�V�0�'���PəH:�?�LNJ���CP��q��"[o��FP aEs���AX�ld���CIT�U��5��C)�s��i;�/_����Ԕ���rؑϮWQ3���,1
|#�MWd�Vb0^ 5�Q2���������C�a�@�S@�%��03B�����`������B3Q;�����l���c�C D;;q�i�������v�A�ML���[�bDPl�#D�L�X
H^�Y��wZ0y3�����k��_����眮U�~�T���f`חrj�uMlυ�#֐J{��O�H�n����������[9c�	*%�e.:<X��а8<��i�)�� ;&���I�È�I��`��\z��0(c���͛k�a'����O�cG]bnHۭ�� ����_�җ�� ����8Ru��::��Mn��Eܵ[.����������ɛ��wl�0�pǳ�4*�h����Ss�j��?x������q(K�z�g9Ddʪ��R��9�E\(�
)�R��a���f� Y�w]�E��S�kȮ�Q�Q�8>���+?�`</��AE�RmL&�r�#8�؊�{!\ɗ1�z����3��P�3�]����ŗ\���\%E���4K�����+�>�����Fqx�<�\@SVCe+�\�B��+���+.��Έ\�5�L�����{���Ɇ�k��F��{h�C����1NL�Un�������n���VN�\uj����}�֭O�v�P	�퉲�W�oe���I>�F���w�~��w���#O�[��?��
ږ\�Qy�Hݷ���<[���?4�(�������,�d������, V�jhU���'���T�>%������j�o������~�������~�gc]ٽw�)ϪLO�{�>� �I�������e�]�+�&i�` _��k��|��喛 ��i�A�;T���֭W_��ȝs�9���ML�"�������?��o�q����oy��82��O�^�}����aы�]|�����'���;��Ua�?����������.0��]��r�}�}�{߻����yu�[#ñ�����9N�2�W+��U*������'���kc�}�&�.�N�_Tƚ6o�<���Ͻ�i�/c/v�*(�t�ҥKל��khh|�Ν`^d�1�|���#�_݀��1R�	�j�O�Z$�m'�,	.VxWWX�z23� �����d���l:��*,m���;�Βy�i<�,<Xի��ܘ��L��� �utt�a���<c;�/��C#�[�{�/�c�ep����[�޽`Ü9�CCC�v�[��co��cF�^+"
���4F�L�s��y�V����f҃�Ǒ1�Pw�,���9Uj������&:J���ɧ�"�B|V�)��ZhGg*ň8�)Gԣhj�M����Q,�q��.^�O|�"�7乐�{��СC02𜀠�_��"�z��������I:X����"���ث���X�!���kIYZӚ��x��?��R�G֍���9��)#���"�vK�0!���R̤�$f�Ά)��1�N�ȨYj�ʜ�<�1������,S��-�-'���`u��`� �P�j�E�y���E�z�S�_<N_�Q���I��U�2��i#;Ts:�s`�F��R�sA&0��-d�3,ڬ6T� �xxR���rf�ʶ]����h��!ϡL�,�z'��x��T��Q� M�aH٥�1��W�F.�ش����mp����6�\�fbb���v__<9G@����=��]���ɰ[ס�L4�cw0=&�ԛl���h�U��ԮcїL2����\�l<վ��@mvF fU1݊�6)����)�6��ę��4�d]$�(�%'d�_ �eہ�$��.��J�8#	^�T�,�yO���Uaj�H:7`[.�"��
�	݅:@!̒�5��%B���X8��������lHW�Ꭾ㘈�"d�-���8D�{�x9+�&_��NU�Yzp�\J�e�A=�C��2Y65;Ͳ��T&��胮�m ^�g����~Y����|��[���b_��)���7E70�d��< �)f���6��xIK� .��B$�d0�N�yO�d1�U0E��ü�Z>��`�<l���DU����ͬ\B}2aZR��^I�G�:��]���
��>��7�U��\p��o��(���9�,�r���7����~��ؔ�w���+_�ڦM_��~�Pp����B���g�%����7�����/�D��G�]��������u� �U�]J�O3�D�}���T�RxEZ��ۉ70�$���>����w`慍RbCVBI���B�a�f`��PQD��(���[�&�w]$d��t�^Tu�VSGfŰ�`ng�r�����}�=�{����F��W��.Pz��°`�vu�oo��������{�+~_��<ʊ֏+4C�\���.Q,����b�@\S�
B\������߻��3?���N=sߜ�N��<�s��%��#�B<�����9��{~<]�/~�(��͛�HU���W���^������>r���*�x9z�� 9�Q�1�c[�=.#L2B�5�kɘ�-�T��%:>z��~��(RǑt55gW+A���L�i�B�+$%�j~8oAߪ˗Ο�`�ܝ����Ž�av�v���;���.ZB�w/šșy�K���C�(1-ۮW���J�b�˺�מ�||b�fOU6�������:[ZZ.=�X{GO�^9p��駟�*����Y�c"F�K>c5�f�+�vq�]�ѰA�S����s�^�ءmO��0WqD�k�*�L  ('�޽o������~f׎��-�|�+��������16� ��MN9�?rx��䜹۶m���x6K�ʫ�+X��O9�t��A�-(�V��sXjyS��X7d�L� ,��$h�L;�PLO઀a��-=윅5�}�,S��E0�w� 1�9Wx� ��?mW��
�P�-��3�E?�xP}�Y`]xAѴ�o&�8�p�3.$�]`�G��UC�B.UE��t���& ��Bbdt�{��"�044�`������j=�Kߝ�s���ކm�=�R��~S�tQ_zk��Td�->�|�c�r��������|�\�'s%�Q��5�i3���F�(Ӑ9ORM�Y]�Ô�2�h�%��"��Z�� �&VI
�\�}ǁ�*@3t�/�"N|���u��P�D�P��t�*>Nt�������Hv���9���E���!������kZ��y.3�m�e=P;Ql�4��_qIǬ��(_�=W���I!���L��*&5�o����i��aAWK����y�P0�b���%�h�f�-�mӕ2(y�LF�=��L70@�}�U�� G����ߊ%t��B9$� ��H��Q#(�Ý*3�	Zq��<@������Av��[��	�çv�E��Y�Tѻ������#��\#��a������hX�n�UsV�MZ0�C��K�[9���S��c[:u��J�U�"�F`���~xߩIL)�:��sx�^�
��i mV�Q�qda�#�U�����EaG-�$��KQ,�b���c�:t��s�_�M~�{�F�&�J0�"s��!���7����)��HEKi\+Fv+\2��4X!X�����Dä6��i�i�ٰ�� ��@Bi�@�Ő�(�X!
V;Y���u{��[y3�8%�U]q�|"��>��x�u�ͣ���P˱M%Rge�&�E�T&9���$v�1�����GFl�]*C�l.recH���[vE؅[����������;��@�Mó�&l��7l��R@ݪ*!��a���@�������׀��ࢪa�.�w4w5�V�H����x���Ϻ�~���ێ�nUtx���	���M̊�W���Zf`��C�!����^|�Ł`���,[��R�\�K����{�n<�d�/�d7l�p��w?��G�xډ��Z&�T���8�&,3�?��.  ��~�;��=w��g?��]���Hҩ�;J�df��MLI�
e6�rx��3�Ɖ�Y~`�.��,N93���،������`&����C���A�b����o�����'�����uZ l�L(8����k.Y���˫ժ�%Qr@���;�2VO��ҥKs��2;�ߑ\}�2o�����O}�S ����JԂy�sO,\���n�Ї>��o~���?Q��w<��Z��e�<�p�N:�'?�	��<��ox���ڂP���c�W�8yd����e-��8�,>2���ڥ�#�[D|V���X0�HV`��ڰ��L�J2��U:����V��ᗭXq�)���L���?�̋(ө���������۷o{쩱�1�j!���i�u�$�%
�
0�Ν;E����O��+W���>|�p������m��hǎ��'*�J'�~�:)�l��:Z-%Ӝ����-������Ȩ�����?�8�c���w�}2ev����;[�n}��U}��MOO���Dx߮����>x0\ Pa����
8���g����xBVFFF��^s Q8Ĩ.QX�^C���н����D}B�� B`=�ve
�&)�Y����+�B������$EF8�-lq.�h�.=�Ò��pu��@2�5g�=á�߱%�^��uR�1���d.	�|ʈ#F,)�=��aW����0��ߩ*�^����&������˗���<1ܛ�3<<��]V16^o������u�J�NM���: �]s�j�.�B[�D���y~�r�f�9Q@�fL�\f�E_Ԕ̃뤫�y�)7&Y&JN0l%����=L`��|^&.���v�w90::�˫�m�X$Y���7"�B
3�mF�lMcv��X>����S�+����!��Ժ��_�C6#j�X��4Y"��s�����:eU0�bc�.x�(�A崎��r�F�����7�)g�KF}�$NM��P�H,�����|�A��z��a�����NŒmo{��g�u� 0-�`v@����?�kP�s�.ķn� �k8�u<��>�v������[�:a٦M���{֬YS-W@��ڵˮ;� ݝ�p�g�}��y�0&oy�[@_�;nٲe�%�5�GG@'�ٴ�d6�R�T�l��ߎ�?��ł ���y�CU:��R� �A�86�n`wM 'S�9-�|HML���`��l:�[C��0@S���<����fa�	�])`B�`ʨ�Ml�MAz!�Y���-S.�R���%#���⺤_��<9eu�%�1R"j*̖:�O�w��dN���ɪ��'qZ��WR��,ޘ��ɔ����	qaE���&r2'�.(S�V���&jD���ic�dr#��3L�=]��з�R����?����Qk�7�����i1�h����3$�����+��00>*3�u�x�:���]�Yf�����Ĕ�W7�Ö�/
�Xu��(Ч">~�'���V�]�T<���yP��^��~�_�ş}��Q�4�+<CQC7���d�l!��DF$��?�Ã�|ꎛ���-�s�P�Ql���L���ƴ��e�{)ۜ͌4���.�I�"5��'�<�!�֩�}���/�G5����"`�x�����|�E>֪ �;�vVT3�4�PD�;㵿��^3�`�?�&�����Ü���e 6����u�/*�4�b�Z'�ұKV�w���CX�+	=�U���R-Y/Æ=��S���G��Y�J\pJ�,��`O^]3m��ԶG.�����8PuµN�sh�S8~H��U'o��/~��Zs�!�W"Y�(RJ�E^�(��c�弬��8N͵X���� �����F-�|.�����	��4j0�(�rx`�^-t�]��V_oG��Ů�p���!����!P��Fw�986Q"E1��a�KtJ�+́8������<�L���zE���^��v��©�:f��?0xxlddtU�(a@��X�Up�OˆHT�.`� ����)Н�:�9T)�cN��qa��Dc�OW`�J�zpA:3e�2 �r��)��3����D�����Q�[�a�T߬W�jyQ;��Ax��y%�2�Q�j]�;�PN���-{��|���ƾa�����0WEQ�|�*�tW�=�С�JȱiG�5o��2��^���]�&&cP�2
��.�,�4�|]��s�R059�z)/a�n�;rJp���~�ԂqDcY�xRD='C�
�I���P�^��L�J*7@� LR ����ڒ/ �"�=�:U.�^�`AgW�aj`J�J����ð;��F�V�hC�NL�0BbAD+'J8N3����h��{lL��&6�t�fb��W�O�4;?�R��)8n�&u�O.ḷ�G�)�5#�@\JljΔ�x��v͆u`LN�W�@9����撹�I���X|�S!L�<7IjB����V������_q��:^��#Ug�֙�/�r��)K�RQPo@���V�1��`���\l梴�o�d�8���KEĳ�O��L!( c�TP�Zjՙ�ʴ,+�R1���
�q�s�ci~K�b�|��E�z]������	��԰F�m(�"("!���l�
�Bm[�)�jzF���-ct�)F?0�BT����2MO��4t\�E�
�*��4�0���������Մ?3=�bi��������������w���1g��U��U�����5K�C�����:��ϫ&:�"��bS)D1uF~әg�}����,����{`-�t{�O�;��P?��� 
�z;���������[��[�l邓N���V� �op���}d%�utA`�rI2���OX1d
4$���&'F-�Ę7d�9ln�0�G5m�7-�Hԡ�)�jE�.��(�&Nc5B�H/]'�|�ʒ��2�H�N\���"�amvy�@�� �*dH����.Mj(��<v�C�'��L�;Uӱ�-�⥘�Bdu����3e I	�k��pHPb��vN��qu��6�ɒ�2x#�OYa�����&�f�K	U�2�d�l<�"��t?�����<�O��v�1�I�P.se�
�g# Tl�b	�<����T̝fՆa$��$�g����(	�S�ԫFҲ�Q�:�>�I�bf�&��8j��������e9�����ai�y��J�A�p��tE߼y�#�<b����kp�,Y�/|�}�{ߝw�y�e�newBb57:�Rv\��KL�׾�����\����K�gWS����?٣���]��HZ]�v������9�e�M�;0Aa`	��ku�I�CEG�[Y����Ҹ����e�#;6�����g~��{��Ţ�8m5FN<;w�C,B
:��R��/%�h�3�@[����r��M�&�^Rgtt���{�g�dgQQ�0x���͛��4�,���f���/^��$�Of.��x#/��w\h6y��b�������d��׽�u�}�b���	/���σE����<x�x��_�2]����~�E���7�=���d�[�h1,���N�7�=�U�����'��ǟ~���������y�9Pظ�$��\%���۫8�Ç����f�u��Ird��H��E'�li՘V�!��F�X,�ԗ	/�����c�^�^�d*~�8]ńX������ո49"�ۈ���X̵����M��J{{����"3e�Hd��+0>9bj�X�a`���Z��F|D���|�=�M-.i��..P�&�eEh��۔gd�1I����ʣ��-9� �Sa`���"���j�<Cyf
��ֆݙ�nd�˖-�Uf������}�V�^��p�j��[�D�cM����R�=L�f��?y��[�IO�,�Rf+�ҝ�@�,��K;�~�nY
�O=���F��,�TR��S��Xp�m�r�)�CXp��v��x��T*\�R0v�dY7\�­�8�q]U���f��eQ���g����=Sk�N�RU���1UC:�z�_0%h��Y�R-�˱�JJ?���4)9������^գ�e�쿘�B�S���]p�m]�?�я&*�A��� �plb
��]wܾw��מvʹ瞫H�:Ѩ��瞉�h궮nP�ȇ��_��,<��e�ҥ��ǧ&�OU֭[�pN��~�Z���IELU�åStW%�逈QbȐ(&�{X�yugѢEp&��~�#��_\��W��wϞ=���,M�U���][�n��p	l���;o׮]��� �$I^Ôr��7��Q�����'��i�fx!��k�tC���ʆV�X����[�����uwvv:�}6������:���sυg��M��ԝI̮���ά��V�pH�{U5_J�r�Px�3;����["@R�
LIN�������{UQ9\&I	�����gXQ鷔�+�.��\c��8�3��q�ę���$8�͛"K$�5D�͐]�qkm�:�2��6�j�F�����!��8�I!�q����G� 7� ��&"��|D�`E�
�eڸ�6a�D��@P2�>�8�TҏX�n��N�3�b˱~����Z�'+�������l�zX�F�d���ӓ�h!�.L�V}Z8���K��X���w�\����ly�fY2��Ɯ��k���F{UF7XHN�"�k�7cY�⥵�D@�x)9	���j2��}��)>2����&]�2��B%퓘���� �A,��'Y��;
l�>��_/Y�2�b�R �~!���7�q��?bN�@�5�sι����qjL�W��+�'����u� e���'?�I�5%��I��ZL�oC癧���=����,�������J����Ҷ����l�?6Yk��wZ�Jl�ȝ��#�]�|��>w�;�S��Ǌ�?��ɕ�l��/9�D:���~�����;n��c��4hY����3��tEQy�H�K�Ē��M��ž� �C,#�\�����b�u<�j>坢A�E�Q���mO<�c��}�ËV��?~��:55u��oL�w�>$�u [Ʀ������"yR!��8Ƃ#v]�LMپ�(o��̋ ^�-===��;�'''��?����X�^�l�1w��	zu��5D/��N9�^��D�`�L��U�L*${e�y��C�QȞOnS�;�b͐�F5]�Q�R1�5���vhW��J�\��S ��0��HG���BƐO�D��E���]��_���G���\�g�6��R>_���b!�l���h�i)|�� Б���"�K��Я΄5�P���]E��*tK5�h��%��|�l��� r�V�j�WkC�[�)�*��j���}m%SU0���-�\�p����AK�xp�,Y�j1!��p�6�L�E�I�lN8�f}����b[�8��S3|-�`��Ԭ"p=K7��Y.��0�>b�]]]`�rN#v�� �2��[�P��u��ىZՇP��k�˅7CS����j>R�Һ6�q�"��&B2H��ɸ!2����n-!Bn5����\	G,;���#�hy-b���~�h�
K�=��c`���d�a��������io�B����R���%b(���`��h��\�0�*�sQjYy�i��s���ɖ�s/��943��$F�R�
 h�H{LG�ammV��*i����Ft���x nQ���!�5�dYl�Z���t�g��k�.Z��}�	�a�{�w���w.]~����c����d��Z��w���a�-����+��}�%d��իW�*��V�����zu�̘3�]q��%CCC#Cc��a9H�$����i�h���[(�8�HC%S�DG�%$)c�i-�`�����͛��xr���sz��j���W��������7��������՜���u��V�rla�tИ�n��W.Y�YjΪ�'���~��EU���m�<X��ŏ�/Z�r݆��x�:3U��H���|�Y co{�;7n�Xw�gw��2&Le��s����.NR��H=��dw��r�I�"/*�d�R�~m^0^bJ���4!���D,��]��b]4�D�G��a��F))�Z
�*%�R#9?ґ�Т0Pe9AZ��PS�TR%ބ��T����YJ�(J�D��'��&�.�~�)���(�W���s�|4e	�r_�lh_��� ��tR�2��(>)��YI���ޚ�d����3m��
��&�a�R|_�V�z4T2R�c�c p�T>��}0W@�.�vbTj2�� ��ym̮��IRsTz������3��㏯:q2��~>���1Ӱn��w>�я�e�*b�rS���7�u�]����0���o|���_���>q=�J�UM�g_¿�Pk¦�i"m�r���za�?5	��5�%�T��s9�T��Zނ��4�$>^���
���Ь!���Ͼ��{��(���g��8�F#�qp��M#a��}��*�b]� �,�O=�W���d��0����xZе�&�Cf��Q,�kb�-6�D��C�-Y�����3��dy�-�|�O?��]����T���r5��\Nv��=�y��>����ll����q��82Hut�R��p�ĩ��*!�չ,���3!RR��X��c�*gEc�000�`߾}N|��a�Zs|"�0��[���]�p��.(棑��Ƥ����� ����߿ .ʽ�5�R�#̺)����)�����R)�N�Tq�j�[?S��[Ш`�,�ct��T�G#�,�X�Ps��
{ԩ�]�
����`����/���
+W�����`}%���R Ѝ�2x�
��c+{����u����09�P0L�cWW{���4ق1T
8���l,�Yq�܉&z�s�z��ᜑ�Aօ��"ycKKkk�lhx}�;35���jhKi�4R.���ݚ�o
��K�_�F�[$�x�[QJ��ar|gJ�!���d��h8�֜��:��{{�`x�1��-�C��,/]�t����t���R�488���M�b���K���`��Tﲭ�vy�7��x�+��gC� R�}�o���qښFP�f��c�^D��^�.O�Y<Ji���n�!Q�!���͛Ѳ���j�(�%GTBY�qQ,��20F/��=�4�fS�8�H7쀃u���sٲe��S���w���`��I�P�I'�~��D��C�J�(u�R���!�W���G��MR:�J"�qQA�vƱ�R΁1?�S�-_��/}鉧w�z�r۠�	���w���ԅ^x�g<��c�<���u���՞yb;L܅��1���[�r�\:@��X�pa�s`��:�-2K�6t������5�TX�v�e��On�yA݊|�S�!�r���u��;:�8W�с`T'F���j9hmO^��7�����'x����իW�޽ۥ�����,�S��LiӦM�T=�����tLemi1���	'����ɉ �F�U�g��1�����͙3g�`( h�d4Կ8x(�9�/"]:�q���R���D��7��ȳ�+��k>Ǝ�8�rM�Ih�����2djr'�J��% Z�O�\^��R�3�p'b%E�DJV�Ͼ34GI1^�����h�hK��,�4S�f��Z,]R�F�T��j�Ri~Y.��%��]�}��[/9���W'�[��m���UF2RS��y?5��K���
������Se�
v��&'�bx)�m�'����sE�+0E�7�:�凪�h�^��������ط� �[4��P3����9Ҿ^`��O�"ō(�Y��n�j=.������/��WW�CEU�{r(���հ�­���9D�yϮ����ƙ��ԏ֢w���, ���q�]8�Oǻou�\�6�˶�Ђ����K��N֑䛬�tM�z�'�ȁ=}me=v�\�=W�����_P�cddd��\7�q�j��3ė��׶l�R$߳��3�A���� t�W%�<�p�nI�������]�O^��Ӻ.0�"�XR�n��{d��p|�3�x ����o�|��^}�go���ke;{�(o��i����8��{c�F��x˗��x �P�x�Gy��4K�f�/�O����	PP���<,SP�z/���&ư�t�9��"����8.��{0��'����R�����&�F*����f�*���BYu1QG���$�N�[���p��n�����dɰr��c
<��� ��/�bTA���I��/<�~���j֙�R��$����\�������I9��� r&+SH.N)�>:rу�{��]/�{���0G�g[���^�X���+�; y�5ಞ��끭c�6�:M���X�f�~�m$H*È+�TZ��J�ӞZ�W�|-�,��8�����(��c��#FV��j�:g���o�b�m���S�̌�8E�����A��j�jCv#����W�'�5�^S�q�Rƽ���\�/��lf}"�))4Kj~����%����%o\��C��W�Z�0�������������˖�0���;����>�u͉'���mx`d"�t���6U���4ǲ��:&���\�r�sN)��h����t"GV��s�B�a�����D�\��ٻ�!�=�L�W�o;E+K�T5)Ā�]���Wh˷��'�\#��ݱ�Xyz�T��x1� �Շu�(�C4D��5M$>�Q�Dq2���?G�����C˔��Q�8�Q!���(�bi���YvUY��:���w�}hxx�G?�X���Ut��z��v�xW��1T��-Q'(�ڝ�I���L��v���!0fqׇ(F�Ӄ�Jη(+T\k{[��_}҉�"��?�(��~m�Ӈ��}�w¢y�=�T�(+A8V�ۊ�gdt��U�z�g���6mm�w�|���m�v��%�^�]o��}-�Z>oZr�u�O�������j.�g7,���jQ��&ּA����iur�WHyh�����|�(�aQx�j>��WX���ð�I�u�Ӆ��=�é�6��q�{�3@�=s���d���܉���f���Z�--����716>00`h�&L0�����(�N;��aT[Z����?8��nd��H�W�w��v@w���\ ��o��%��sQ�٩�4���8���z�]Ͳ�"d,�E/^��v�À�U8Ś�G�����E3m2�,��N�EA�QЍ�ScuP������0t�'�V���4�:(�?�|64����FKc-�wB�PEe��ܘ��&@���-(���^<Ndw���GVetEi�g����sR}��^�Y��"
FT��#��\㒜� -άbwM �(�G���Y�V&s-VD��u�5+�Q�xSW���͉a���7UShPJ�e�3����s��F,�I@)��鉔&\��U��W��T�S{�������S7��=OM/�䒋/��S�cj���ƍ� �����k���g?��_��_���
������u_,�0�;v��C-��ݰ�\�x�I.ېA�Z.�	�V�a��0�S|����4�L�y�����^�R�{]꧴iӦo}��?�0��$�JH��E���yv��	�b`W��,�XlHX)�P��A���8�������?���֞�l��H�U4�$Iυ����5p����;��f��]�ů���~���0uU�������߈G��� v��ɖ,�(�c�x�y�����4�Ph\b9���~p�"y�+O�z�	��}�_]�&��9�D�2�Z��ޑ�K�9�#�n�(� �10&V�YWqa�P�:g¨�b�ƾ:^r(�YE��OK<AQ�פP��lE���z�,��V��%e3xw�q�H�^��E��MlX�!}_�^��8d��J�E&�b�1!��ײ��#R�.M���.��@�@S�+S��3�ʡ@P&�ٗ��֢�\�j�3֒B/6��b�����!M�����t��P�8::�1ܨ�v�.n�)6Ǣ�{�ȟqe��&�V���$����|���wg]�� /|�M#`$INLL���	X�T�P�BH�"{����G)�|ɝ�,�4�O�)���#+5�؃�S�d��@��j �����͓� �L^�,�4*g�P�X���
��&RS*&5ՠ�L]R8N��l8�.���8�����s� `K³��dz��z���۲��5k��j� ��p��ϻt�C�
[�p���	�7��E3j�M��č�U�yy'rRM�Ӯ�)O�aM�-\*v�p�UWWWm&�F��
��(0���::�K��ߑ�| l��B�M�q��o�A$�����h��e��ДE�oDϥ<9!���Tf�^p@A�Z��L�~*�7�5<*������X�8��8`�J�6�(�9�+��4��dk�������c��	����3˽Y:�Ǆ�������M��u��M�I?7���s��1�;P�%�r���2��z<�v���Y���%�!q�	�|"'���$�^��h�xq�T�:g����U�L�Mg�&�7�&���T^�M������>KM$̼zYq)�����kf��kI�`�籼�NsE6�|gT�tk��$ϓ䛐��ds������
I��R�.y*tR�qN�Ӹ��5�Sͯ3�ٻ�W���ZN��S�=}ӿ|�{���OYC����rˀ����	Ɣ�����:ZZ�H�$ˎ��g����go���?�bѼP���R53ډ0)`�1JЊ�}��}����k���#��2�*��O�M����#��b���²�%�
����od�IX���$ҳ���-��>���X2�g˻/���N.
��ȂS����K'�G��,�b$]�=R�J�a��ZU�ہ��>[W�\4Vk��+��������������o:e�� ��O� �I��S���ʑu�G���a�������_��7�s�e|I$����!��֞������s;۰a�pT��s�̛7���E7$�Q%Q���eJ��Yp'������ ١q�9gkc�z�,�Kh�3�4���xdkD�VE�k����G�^:�/�&h	�S��l�����a�Ce��X~�P�)��˔[t�*�GX}�ࡻ���_� �5�e��1au��|@/�b�P��zA��@����ZZ����e��"��z�
F).-�l�>�0��ꅁ��A�(/��^����|��4��cOG7,��P�!��^@h�T�F�U1�`�f�h||� f搐�>>�¡a�6����6j����h�*l�V@�
X<>�jfx��`��802��=݈e@q!j��2P@P�B�
��qu��
�OES�^��?d ���Zerzr�n8�{Vi(&b�&s��yJ�P9��)�&���fRX�}���3���D;��c�ʕ�۶/Y�������FH���t���ڵkW�\��/�� ��~��[ZZ6l8�vp�0?g�#� ����4k����k�g��d�6�8��(�<f�x"����WƔ� Pe���3�j�L�9=݀�*�����U��5�|K�IN���V���Z�c�BX���`B���vn�B�j:ah:"����e�`L0q�zg�m�ܘi3�8������(�B@�:,�0V�|Q1,߮���(���`Y������Ka4��b��;2��_�ڮz�a��&�0n)������PKI� cIJ�|҃|C����8�3].�R,085ݷl���Ʀg8�v���x(ɧ�v���l:��g�q��e�\�ztH���NL�5��\���ghr0J��Ŷ���h��ζ΃�����v�w��|E�Ptf0���_�z-\gb��͓�TX*�k�]�*ث-Γ�T�,3���d�Y�z0�C�鹰�-�l-��05��#ãccc���:X�W(�$�س{pfz��SO]�l9 �	�q]��Ol�H�PQ%�LjkVcP������C��~CV�(�G�f�B��;
�4�~�<�`��~�X2@��n��]����\����_xf�,f���I<���~����|)1�<4�E�`�*�Yh��dRQ�-X�!����lI64��Qk
`%�%f��db|���`,�� �ĭ!�u����A�j2�a6�C��PRh�(!��a &r2b�C_�"T�Lb����\�6��Dp5�c�������D�	j�����e�/v}2l�e��5���:���g쀅�1B�?��M���		�=Z ����P�9����F$�,���.A���p
F�"�ڼ�#�X�5�t+��)1�j=(�)S*X�S!��?�E�^��ꥎW֢�5.�-[�,�����o�f��.��BrcaRoL�8q��)����4t��r�U��n��Ɵo~����ߧ���Y`��������+`-��R�U����g���Qy������2���y�a�_�"�mN~�l3�Ǒ��om_�0 ��o>���^~��n��#�<b0�s�;��vMLT���cA���}�IK�b>oc3_j��(M��H�Vj3���m�ݶ���g�u�[����v���P�7�p���%Vo�����6jr�t�M�����]w���w�cS�B���j�u�����_��WEkZ��������K�䍯	�o������[�PK���&��D�/I	��L�0B)CWRU,�A
.9�~�0�{�RwQ�o����V����-b�s�źhr�5�R����1�:z�%ZQ� 
�[��G��Ęi�/෸VǠ�.����f\��a��=�y�8 ���0Y����Sv&� m�g�x������)�E�cP�^Da%�Sq�2��pę/��G��ꓽ�pe��'j��q�$&��sq�>����2�l[e�N�;�>7��#��_��̲�L�W;U��U����	�mA���2" 0t����{媓���0���3cQGAAQ8Jhr@��C媽w�+�u�������=��^�z���]���k�������f%�B�M��K��K���Nc���T�$�K�w9��	Z�2�SJ�6f1%o���p�D�<I�9b������{��Yr��*�!~�e��W�Y��82H�Е6#gBe7�f����czz��-�/_��:�j���[�!n����㚝 XXt/��C�7rZ�����G��f�8�7��#R����_���?�L�r������ؘ6�8p�֨ac�H1 x磹��Mڕ�͇�%���ɖW�b�Dt���JͰ�N,Y�D�a>�&_9k��-[���GFF�{��bB�	j����ÓD���_��1��<�-�(�M�����yc�V}eI�X4e���XM���s�*��M��M�?�>�a�C�p]��G�)��lzp%k�b����X������;p���xx� ���\��]̯�T�!�
�~�����5	����p���W�g���)�3U�j;$16ƑQA�j��闹�Y��t����N����;	��7"i��V
"�Ge��H����ީ�o���ɯP��D�.��È��!�j�P�i�r�,KDܞ-�$=A?���)a�z��@�������w���YЕ-ig��+��<��񝊗��G�^G������ۄ�9Z�d��2���=����_���8�������d��D�0��L9L5��r��O{BN�KTU�>�>dtu�}3IKf)Ǵ���=�'��g�,<^s�� ��=��|�_����.��ګ��˧?��#��"�s��֬9x`^�[3�.�V�T���&���Y�W���~�+��+�٥lj�0�D"յP43��}�����O�9�s!�1"a۰�����ZM�+}����&��v
䫱�*�ORg��ɜZq:(�(˭[��y`Æs�l._2a0���#Ө�?��O}����v�40x�4/9�Saǆ������lp���b�����i��i��(�kN9��'�|�ξ��w2U�	I��f}������W�͡������p�oy�;	g9T�4�BCh�qp�X�a\�{W���~x�O��1�Ţ;����#*�:�}�4�d�F� �6I"��̬�LP>Α��W��D���Х	-&f$)��B��L�Z>q��@J�;yD�����Dz�T�I��iJr�n���
{(|�7�RcnV'������1��S^��Ѹyn̢��蝴Z�m��(��LO�{��%�|�ei���6Zuߋ�94Z�yj�=eд�&	p+s�}�lߵ�+L�*��Z�xI^� ��w
'��X,��,9�
q�z4�E�En��S���]�!�?OԄ
�&��{��a02]�X�qn't�4-��;k�p��8��{t�X�~���^�1���3��۴�����\�G�$=�à��9�Z���X�W��B��V+���/!
(U���&9�P��wO9~3�uj���h�TVH�I����g[����d�4��5��JԘGH	$�Em���wG��e�H�2Utݠ��i"M��+�/���16~hd���e�-^�prRsl��U�����m]]�3�<s���ɞ|�IxRK-���s�l�]�h�q�����*kq*�_�%:�XpVbf�xB��a��e�@&@����k���h��#�j��kw�KH�L݃��2��\�b{n;E��S$�T��7�uf��4F������aW�4Cܮ9�N ��S�����ynvHw�}�fbI��ȅ-���`TC��U�|vk`���p���ph�3�i�gʓZ�L����α�ы���������l����R&b|":��d*��;qb��?S�@nfD�{h�t|j���X/��|�n�UDn8<��O�xq���"��l�{'�$����&����Z����R��2�4덖S��MӖ�vZ�� ����I��{T�6�_��6,9m������	x�\���!�����|睰ߎ[z\ˏ�8<s�I�QC��>㮻�w����z�)��?m��>$C�������_�淬]�vbt���ըl��`�IkN<~�%�]}Ã0n=U�K���%���r���4x�'�;E�~%�+�����V���L��b��j���Z�͜��b1j�j�%�[w[�����t���Y���c�F䉂m�6����B�����Ű��*
OB!㔁�԰ry�������|��牢Ÿ#�&:��_ٱc�T_|���977������:�=�L	l�!�Q�G����b��tL4�.��)��	��
���������AI�zrD�~��_��+B<
SP*�{w|��>�-�e�4Sb1Ӎ��eT��Tj���ן���z�Y۶Ԥ�����8rUż�ʫ��v��X.y�[������>O�<3q>ĺ��hC��-����+���y����L3�<�f/��_|��~�w�0���*:��I|�F���^�؎R8�ø�r��3��>mAL*��ߠ���9x�<E�i�Ė�����,� !��|�`��J��Ų��I���!�+&o���t7Vt�Q}�	bZ�2v[�@�)��HE(#��p�i5�P-��45�����^v� �6�b�J�b?m��Q�0�CC�y!'D;tDJ'�<�qH=�^~��Hq�~��F�{�W��O<^s��]dQy�y�m�x�9�^��/� c��FY�6l���ɟ|�sB�
U���:�� \n�ᆯ}�k�H�$���=�y���^�e� �hh�D��y��w�7�a�
h��w����9�Va�bncQ�U��/�@�6�L�9G����<�>#�Qn���>����B������O��on"};DCzH�`gHˈ�y�vr(�I����w���x��֭����>�G_���QzE�r�����{��w_���Զm��NJ��uƖ��f��������k����ȹ������z��-������Y��_����i���R@N�;�&ykm@X~��Щ,��@�0I2��ll,��������n
<]�Z;I@�c���:�*�^�C�i�OK�q9��/��RCV�F�*`�T恮�A��Q�Y�*<����C'r'�i�ZX9)�:�ꗠ�Z�Ȕ����z�	�:*J4��i��*�OLS`���`�k�N1F__���p5��9��,_�|Q� VϢ�18v�j�O���������?��Y��'hۼ(��̦��E�MJV��<���F�xE3,�D<^�͞��))������8��wGoƈ�U)�+���4;��J�.��6�t�M����:���;��������\.��:N����H��g�y�!k�;Jj8wP=S%�7���ڠ�>/@2�:f���I�.�x�\m�&YI	]�l���<<q�s�9�dp��Tn��T�G��p�JI)>%� �!��V�cyv�b�n4Z&�t���֎H���x�Y�L��0ã�5�p_�=�	����Bm����|��,^�XΕa1����D�*#� N]�1���Fw8���*+���D�(�X���pZ�u�KROO���z{����Tv���4h�M�p�T�����{����m333�q�x�4��D��Ç1�NT]��V~�����2b*��~��j��\m�:���m���񌞗J:G_m��+��dSP-;���7}��~D|��JB�[XCcf*rT<?�Æ��.n'֟ ��jՏb����_ ��������L�\x�b�y䤜i�'8�:w�Q����+� ]R�Ox��g7l8�X4���P�)���NO��#����h^�����D�	�P���ҥKx���N:�T%nN�E��0m���7���߿��tv��k�'��>�G�'x��Y*,K���. ���Ֆ��Y9�+��mX�0`i�����E�+���J��*�eϬS)��8�A|i<� ��w�M�k�͔���c^RL����}��� ����FDpF#a�l޾���[R�O}�_����z�^���\��m�`>����_��U+��6X��K�)�o�x��\q饗�y�_���}��7�~�[.���ۓY��cV�t�*GF�G7]	>�'����7��$&��+��	��7��=�5c�"TBXx%*�ߊ�5ka|\�4i�y�Y�S7n�x�E�.��W���'>��[+/qL� ���j�9^S��S�`�.[}җ��+���MI�5�B$B�V�u\\g?r��S7����Ϛ1�LAЎ#�B���Y�;"ڣ�|
0sb8"j{)�E�qԛ_��cpgWgQ���T���I,D�	Fg��z�|BM��,vI�y�[�u'y���}�ê�3P�I1�`����d����صkI:�H2bqbCt}�_��/}���-�9CLo{r���B1YY��d'v��ؠ/���!\(%���������<����
��%
�E��65�K$��8��ʒLMn�G�I]���
5y��Ct�
TU�F��]�pS��$Y�Y���h8N�gPD|�X�Q����9��۶�b�!�����:,�����&ID�b&ے%��m�����UtGd<�f���ŰH ����E�&� �'.�!�y#�[<� �ꑑ�m[��9�9x�	�ly+0���-G���9�f�A�I�Ē�~�-� =
y�zHB�&�m�&�$�#@v�[c���&��H��o���2�b?�8�E��m��	�������p菍�4��?Z�h9�WPi����]�|-/�\/r<�,�[��l�����'׽:��P��bQ���M[����)-���cY��+ǌ���Q���~��� ��a99�+c���G�a}'��ɤ����t��8�g����{� �6����۷o?q���bi�b}t���|.��g�}|oS�:�,��m�WK^\���Ua����mۚ��u�/L� Xâ
�Z&pKR�^	�˄�z$*�1�����Ll_M '�Vql}W<Yv�Y�F����u]"Dx����P�E�T�,�^I����&`�����b�3�Lu9���A�@%d���P��^e&�h�:��r���oDX�رc�2E�fE:2�J�eī=:_����ZV|ԯ���QR�l� CN"�V�m ��خ��ryx�RX�C�Q��kM���HƠ�@�6�4�}��+��)W�����	R��y�}��2��AdШ�󪁍s
&e걯��ʱ�q�� �h���#�_,� zw�ju�٬�j�N��gW�X;��[_|�I��-�w��dc暥�a�UF��Әi���>Y��Եl(l6g&f���R,v�Sn�"HƲEK����w�5��R�m�hN��տ�����韚��M2��v7$L9��O���vy�!�w"���T���(Ě�/V�^i�_<��Uwf�\�P*h�Y�d�nd#�6�)��\�Ɔi˖A}��(���)Zпm˦�K��"��W���k��_�UB��L����r�-	ox1bA=������tIz��h�hCME�KŢ,� rJ"�"�]�Ƞ�m�eME��~���/���o��{�m?�uM߷�ڵkၞ�~ݖ-[	,B+1J���n����-�K��,����_����������v�t#���Eq>QB'x���?�N$킋����ߊ�V����~�[����?a��k�y)����ai�[D�~���y(Qm���*��a��q�(D�������+
C�E���u��1�8#��Rn"m;��p�<��K03Xf�H��:X7f�/�1��n��L���r��aF�⨩�D�e��+�9-?���?�t��;��S�q�u_��?��~��+e��oɝw�ޒ��xq��'��e�sVLٻwTH������q�߽�G'�R������m]�/��/�MRk�f4h#�,�����L��y�k��������Q�'ݤ��8&��o�񚋵���^+���X��Rox��o!A�r���ߔ�6���L��������w��`�7\0�|��׾���������}/�	%,��!Ϭ�r�j4p.����2��@��>�HI��rڔ>�f�Y��S��F
1�2^*g@9��-����ꌢ./�
���n��h��^ ��V���^��nUj�f75�"0]��i�ʂ
F�4��cH�gh
xɶ�c��K2wK�a��F���s����:yZ2X�G�u�h�i%%���W��T�������	Q��u%,�4�,#q�P/bz��>-C�a�JW.\�-Ux0�ur��m�,GQ�Y��F(�
�]Q!��4"7K7��1tXcSCִ�6��ZxOˍ�^�C�z�N��7�&�4�:����*x�𥙁I��$p&ʦ^�@�l����
9�S�l'0��;L��X�T��>
?bߋ�.T������q&�'�ڊ���ɂ���R������0�H�������.�?44ĥ?n������5pz��F�EWUiS�0�1�XpJ�B>B����"I�f�ĝq�x���$+�q�I���vE�� �\҄-Q,�C�_����Q4K����4����j�-��B�WF���������Q��9)�Hg�r���fuN�$-4*�р���'�ߥ��W�Z�P������a�{�c;��Ll�.ʻ7OP.1�s��g�\�ɳ=�e���DvT�t�PN@�����2��{�o���х1��s�=��*B�W�I:D���������f�T�/�9�����U�8�8ה�-��Ǫk�;*��K�u\��jp�����Q�F�qX�0J�0�6��V��!�#����,�����H��T�{�.���������9a�R�j!�_�"O2qE������
�G*O1�/��yq	aURRg:�� �I 
*��������T�u*�Zp���sZ����$�E��B��T��SO^k�1X�-�҄�����x"�\��c�l��h���Y
ίrËO��24� Օ�vKZ�{�6������� �W���k�����X�-Z��x��>��O�sΩ!��YZ&�I��W�3�ټy���[���J�s�J�������~�Ѓm�pf�:�������~����uo�馛.��Y�=�$��y��ߜ�g�����T=�f�i֮]�6�}&����q�FZ�_���g�����,V\�d{�}�nVM͔jVem�\}m�4Z~�	3M������e�~���z�������_��_���= ������C�����6mڿ�C��?��?�߿���������^��0�˩��z�<��C���K��
���>�iCB�M��B�������W\q�m�ő�cǎ�/������/|�ŧ�vr�Y��[}��b-�2)+��7�{�ΑG��U�Y60���Ȉ�H+�(׊m���>�O4�`+<ǍC��%S��{5��� �����8B�#���}S�)��z�+D�jr�ī��w2�x3���^���%�x/�R@���\��s�:� ����A�C?����0Êm`�4�l%��)4Z�P,S���F�Fd]2�<�]k1P���D%�1!���! 0L-����1�,If$��i$��9�"�P��^�K�[�(�X%Cѐ�A�Z����rI�z�	 �|�c,n�Y���+Җ����q�1dC��F0&�/,�����\k��lJ� .u]�Uԉ4!Jc�P_�٧�Z�h�^oւ�����݇�����X�MU
cYj9	
1A���ASB�]�&�����I'7Џ�7����#�ھ#�U���6�|d�P�1��Y��1���[�L6�Xac ���� �d�l��3�J�z R֣�=UCD7m��#' &د�.���A0ᗫ��b$Ř&�5�Q�q�Nc�fĲ�A�ԴBHf�J��y�� �Z�ڮ��$90>��d�:*h�z��V�`W���9�ʉ+��iI�A�}�}�:fX�z�I#� �ԉ8+��2���a*���~�iZA���e=�U-��n��b^!HgW25OR�����r
v��T"�ÔNm���↔�)sIJ�x���ͪ��4��N �{�b�#��`&�ۛ���\�������#Xy˦��J�FW�BO�^�C��ҏr�$�)�X�G�bOEI�U|;N�ԟ�c骢)1�`�%�t���&��Ģ�R���b�=��Ȗ	Nl?�T�y��f�R\_K�.���c��Q��H++����Q�P��&�8���D�ø�8Ͱ�q $`O������z�V���)�6�$GLY1 }皼�C!m���9?��˚��'L�S�TIw��`}l���*M�ۻ��1)���ʕ+֞�?%#J�G@�Y� 8QГ�����(�	��(��dx�k��W�>�i�ԩ�M����6v��-"�8�!��F�{і��,L]��Rci|t�9;ϥ+�$(�iadD�'3�F�{�ӂ�9P��r`/���Eɍ�¾�T�ǌ���',Y�������� `�l�K�
�o���%�1ڱ������CYA��X�a�M�4x�!\I��G^�؏ԋ��EY����30xIH��0�o]=?���8n]V�� �GJG��Q,7%���*v.B��L���-O5�3��xI�2-�������Jy��+�)� �������u�؅�&�pץ�0f�<��0pp�X�tC�]�5�V2o�g�as�,t�S
v� ����g��X��W7t�_����{�����k������0��hRW��O��ǧ*S'���|	U��2��YT�Qb�iJjn��?�X�$�pP�+aK��Mx�w����?���Xwƙ�T9�h@�d�����l�¿���`�ۄhy���o��&�7N��7}LNh,�0	tX˛o�t�`�ٳ�[߹�'�H� �BQ3�J5�ܤ�P�Md�(N'Im���=�J{�F�����5ާ��Ǹ,x�*��0��s���P�T���|�K�k��{�gl�:0��u�;����s�ŜI_�o{q3�|�U�����w����}��"j	�L����w�z�z�#Ŏ?;���]�q�����m���H,M3a�bˋ;��?�7|�o}���b��n��ǚ�����J��իW}����~q�i'|v�~Yzu�o�񚋵�dò��91�&��&@�lѰ���8a7��	H)�|�I�eY7���Gl�@ө�NQ�\N�VƐQ���a}��(o��{�'�i���� � ��M��]I�jM1Z�&e��/=�uf�$4*���Y�R�\�'fޘ ��2��x��p�DP�\V��~��\dL!�%���	y��Ԫ ���Ѱ�KP��8p[��EB�\x3��ܸ�8�qGt~XI���n�}�ؖ��B�cNh�&"�Q�ɩЕ��TFh�}Vc|��n��/�t�2k����b��l"��B@g.�B�J���
�mD-ݶK��%K����aU�{�9�.�Lõ,������F'���72:A/ܫ���U����s��Im�+V�(䊫V���OOO�߷��X�]x�����w?��A��0�1��Bd6˂׍:��批\w�!����$1�Ō5NT�16=���&��SVg�yV2�Ϻ-Z1��@�����ϙ-,M��Mq�Z�=�8f��l�6�\��'{��wc�Y��?,�Xg�<\y���lUoNMM)]yJ��FDyw���q�Dg��AʊZx��A�\�Bq�Հ�B|�V�T���.��#?ƈ	�Q��,N��p%�;��h��1j�lG��}��Q�6 )�)b�N �2�fgg�lٲ`���?~nn����l;w�k^�z5<ǭ�^�(m	�Q�s��w�ʕ�z���0��qI�����x	�{��e�T�F6	�\�W� ʘ&Y�(���N�%��jZ*�ѩ�E�-X�c5D�Ԃp�޽
���񘩚<֒��q^	O�q~]���7�t0[Q�Ng���\�Oge�ƫ��P���~��N �9W,efk�4%�@N{zzT욋{챇z(��k��w]������������2!|ºUs����/�\��]�v�S�7n81�b��dZ���|�k؈X(,^0��թi,�����Y�f5\8�p�:u�x��p���`z5^��3�Eԓ� �������J
�j�F�-^�?>>��4�H��Fb������5U��8�od�ۄ������P��=�0��2W�h{�"%Kxn۶m���W_��s�=���;�d�q��Z-x�����S�.Z�p���?���a����� IG��H"�s�֭�\r�%� +���u/�Gh� ׬�@םy�fWO����M���0�Ǔi�)#���X��}���>�������1����۷�r�;��A��?�=��4P��|��ߝ��^T��T�xZ��tc�nL>��%M�4�~r�EԄ�^��9n�2-n|ذa��'�|�����ӟb�;)Hml^d�>�q�w�ҔQI���_�Ȧ@�����Y��g�_!N��@�ɑ���ʼԆ4l��X��c���ˤ{u��+e5H�� ��656�#�<266Fm����|��k׮]�t�;�k2�����}�X�E�U}�����׽�u�����)����X�u���o����0�2�� �]��\��G,��BS�q̲{���qt��o�񚋵��b���۲-;I�7�M��2���P-X��*�D��(�\a�.v�Z��@d�j�� Q��l?"+�{4VNU�aOd*2|�� $[����-:Z�ґ"ɶ�<��R&�:P�/�����Fx�o@�E�[Uu��xrU�!L��(q�PM�r�A��f�2q�LB$,=���?au�fC�����SΪi�zD��]���Y1d)R��9b}#n��`�iw!�-���|1�g���Q5z��a�c�"�|R�2����x�DD�Ms�R�����j[&
�d�&B�B�kz.�a-�33�"�ђ%���X�Y��N�"���л�Z��=�!����J#����3�ї6�&W-_���r����%���+�8�]a(	"�Y�ҡ���rc�pe}ǜ��>�3�h��ME���f��eK��>�e�>$Ѧt>�$r��K���(]��sQ�\�ak�]rn�u�=�sf�OU�Hcâ&k�Z-�&��b���00͂�g&�x{6vm9N������sBs�Z�]�22d[�Lb�-O�C/��O�
�^�C[R�8�>O�C��G�/(�;إ`�P�����zT7�Ro.n
CR0 AT�&�Yl4���7
��r��]� �B��jz��R�.��\���E9�@����=-�����!�%��K����r	��w��t2��� 3�j�-M��T���mW�x��F��6!=E1���l���	6:�^�u��,�?95�~7�k�R���Y�����m�t�M�ؽ*Lˌ���Vܟ���rQ���
TY� _�b�>����b�� q5�Lr��Dhh�+s���
� ��blt��Q�m[,)�h@�24�!��ݛHq���r�.�\
�E�,����f'��$tU�殒W�	��δm���IX���e[�	��1 �x��S�#��R�1�0L��ڛ���Ȫ^�s��I�5�����,�!\���%�����Cc�N��V��^δ�f���#;ȪKz����D�kU��4d�<a�k���zc������h��Q��r�m�-�f}����m>|�63#P.q��B�[�Ltr[:9���>�:M�U��tU��N����*\��8p@K$����*c�ǔEk�:;�h�y]��\>%�*D8�W��6�`���8����� ކ��qI�%�� &�&bŀ@��Ac�6� �3cOAƞ,D�Z\�j��+�a�O������{K��;nŪ�7��F���S��J�E��jy�.��s`�5ʹ�2�qD�g����u����9����2u1E�V�X�|�JD�),�����ػw:r�AzxQ�pcdx�J��H�`� W�vH��L)V�G�0ϯı�$T���-[��}*�hlA]&p��!�WB?;/�4�0&~��r ��|��wǞ��?���o���W\Q(�B	E₂���0-4����͊�.^bڈ���[�i��б��/XХ(~c�q[MEk*b�Q��
��R	L�@]+���r�~�w��R��t$��Ȟd-.g�4��5ǹ��1�� _�<r��/� ��
bIBCN�:0KSՁ� �v� �8M�h�N������ǘ<p���ſ�/��-w�q����sjf�駟������5�\�|��۷�_�2�g�{�Vo�N�ժ*"��]}�c?���{����� ~����O~z�[/��{��ۊ%]��Hj5\���?E~��g>���>餫���0Z���N:*����ߚ�5k�A]��*���&��R*�QcT��AԀsiYN���u�@�b�C<w(��V�"KQ��q&Aq�h#�[��a[þ���=�x���'~�->�6�1�Pv�_ueP;�
72VXB�T��s��)��_���|@�r��D.�;E,�6�L�PF��BQ/ʴ1s"��5�-<J�W���g�>4�*a�����&'�����m�����l5�ecw��s�Tg�׫Y��T�|�E�A�����a�ҥ˖-�^�|yb��v��}��ڵk���SO=u�#������!�}�"���A(�}�T��H����z��4���Z��, ? �����{��"'"j�r����鎍�!DU(��8-�뜫�0>1��q��̞3�<Ӳz�o���ka������I 9ƴ��.�-gzz�oIp�7��ꡡ��+W�&|q����	���]��FG�����:P�V����[�n]�s���w�n���<���?�|�Fp�o����~�b��~���.O��;7n�X,/:�U�V�5mǎ۞}��g��7�a�Q�:�#M�_X������h�4��إ`�Z���ޑ�����M�6)tN�q�K3�tnn����waJ��%����E��!�8��'i�~�����y��(�1W���W)�/ݟ����Z &�%�F�!-*W³����遅�ծT*��sϞ=��k֬����LC}���^{u��"N����H}���ԙ�Bw�O��&F\�:��`��+"���U&U�B?�M��ͯ�L�(z���Ck�Z�\��Gϲt��"��R�2��F�W���*W{�$,o�3��W䉍'�u09E}v˪E���0�����ٳ,3P��V�I�KT�iO����g@R@�y��N��p� �Rʕ���I.�-�P
�Ia��gnr��g�߹ufff�SO`�Q�B0�.Ĉ?n�P&[�l]a+�wZ������H�Ҩ��PM��<"GV	�
8[�)�����
{/Tq�:�K�p%�����"��
(%̪�t%�{����M���W�3j�>\�lӁ5�S1$ ����R(�0����˪�Ih�·pcYH�,83�J���[K�%�?��ԟ�seF>��n��?��70�61�*�̒1r�SR©O����bP�K�,��ہ�7�̪�t<��Ӡ'��}==p_�F��g�g
|�R������"�8�/��r�Ǟ@�T'�ˋn�.4���z����"����e�]v�w��葆!_���~���D`h���ْ>���b�Qk�#
� �pp��ȩ�;���ʳa4ǫ"����_�~�?�5\0<� ���YB���:P3@{S`�*˰�f}v=�p�cY)>�r昊�8����$��84b��W�7�hCi�����6��܉C(u�h0ܝݷ�����+��g>s��w_r�%��8����σ�GRS@�W*�O<��ŋs�k��'�"�م}u饗�3�{<�
F�,��|_s�UM��=������W[���EQc���7E���?����M�䧝~:�E-̀�R���x��Zl;��I�>%z[�Z��h9"�;H���FI��H��y�5&���WAL�H�	�Lb>�tOQ_un��،ӥ	�+H�6LoP6�,���JG�q'�ɗ:��I�:Z�������H6�/�����K�����b	�!���/���z#vO�f��ӎ�I�;��]��i[ż�PDΊq��Gd�ɓ5	���1��f%1jF�4e)�j�nД)<>�XM8C!���-C��H�H� :RA!���n����@��2Nv ]�&��3����P*�|:6=c���w� �����.�g��>F��V,[�|��e�����g]�H]�\Y���n�TF�����hV�r�����������)��1=U39�<W�ƌa4J��hUfG�������[hF��vT��M6��YX�09��{����S�����W��$v�bo�w#�{!2�ڴ��	�7v�$�Q��R����a=MJ̦��Hw�|�ZйӉgˊ�_����Y9n�j~�ۦUX0P��'G��YTo���AԊ�ˎ?~��?S���ѿd�I�φGqWnp�/�ܻ���n㬕�c�>49�rf���h�VR!ǞLY�B�A�e��h
��:�﨡�N���li�\��u�LZ�a����0.�l#���X��m����o5c�aK��'[��/v�ˎ��Re�����oȦ�˛~�g�E(��N=q�܈I|RT�RR�L�c���y���_f��v=)���:��a���d��	��}`\{�z.v�>MB���ϛ�wx��4�.f���y��E��&jT\���x	�!i���B_�2!���$ERf�M��Ʋ�lej��ݍu�6�3++��Bc��ʅ$^B�FV�ڜbZ��c䆻z�[#��(a$�O�$��[�3硸bF������8���/����E�V[�d��o�����El�l��f��-�2�D�@��^�@9�Փ�R�E9�`�My�R���ވ8ńc/8O*���~̵w�t*�&�g!�Gwpbf
�`!lfǩW+�`���J\�5�{>��&�����ꚤxu�B ���;^5&#[��j���.C�K߱cǡ�U�$J^G�Ҟ�����άj����f3)Z89�S��x||���ߛs�.-�_�u[n���ME�-�l���}�(�]��o�VN�=$��K�BwW��8	=ܯ�B�8�BJ��E�`h�h� ��L�FTȭ�j���-/k�h49�G���,�=��2��;���K�\����'���L<��}�q�-_r��`��W��ڽ{�/6� �ut�����J�X�DM<Ⴟy���\1W��ߺ~��x���3so<���+W:3�Z�RR6=9��s;����i(^wA	������{
�(R� r��V�9+�6���u4�uv��p\m��8I쇦i�]�����\.A��<곥n�B��=�B�*Z��a��`.�������x��Mc5'�(��V����:kl
� "nD�X�!�S|���aK���5��sE�.�;���^S��d�"H���^�(1t�)"����f3�:��$��f�N�p��hנ8�#�=�ΓHGN�e>;xY�avB�Pi�i�ǏT�h���|��w_�j��7� �ݪ�~��τ�w�dQ�y瞹c���\�(����,�t����伳֗��۶�UlIݵ���K�e�0���x��(�`!w�Yg<���٩�� ���~��|��׿�<x#��"�Z�ঀ���^8���{�0�t�G����v_:g�:����m���X+��8�Q ���<��`��*֢��,R��1����ĉgA;�y0�7LW�**X�O"� g����tp�w<�2���ב�6�R�&bⰐ�%��m�-���x�߯�1�9��Nx�g�̒%p��g��s���#Ӻ, ���.�b!�A�t0l9ufRp�ǡ�CVШee6D�&\�Y���=��!h~XJ� ٙ�B&ؠJ��>�fHV��~ �Nn��4��� (0R���O'S�;Sm��7�)���i5C�@}��^�θ���gG��~�j�6D�W���ٻw�wܑ+���X�%�X���.�Twq�޿hѢ�ޮ����@/�g|dl��=8���
������#gH�X�|������n]���u
|�J�r�|��.�659	�o�`e��p6�B�&6oޓ��KOX�Z!��0+������ ��gDI�6�H[h���L������'w���uw#^VO�f���O?����EÇ9x���А�{�3�<�~���O>��;�ܼu��7�w�i�m~�M�6=�ē����Ƭ�0磣��vǜt���y�Z�g��?u�`Q� �"j�����T8�.̟��%�@�T.#��X�+�a$�$'O���l���{4rƁd�2�(�;w��Mn�J큫̈R�/m#��6��>R�ů;~�KCt�f�1::�l!~<d�9����7�ps#J�H:�~5ۘO�x�D��T0�q�j��]�rJZ(�R�R̀��23Ğ�����s��Xw}��1��h��ĝ2(aJHD)LNj��ҥKל�
5��"��$M�����N��?gۏ��ώ;�$3)�לg�l�v��Ԥ���p�0����� �9����k�*�3�Y��^�pj���R�� ��=��*�n�AC���Sia������pS�xX�*�{�<�"�A���� )~����*8�.$��9��.������ݵ~��O���q(M�J�sxgP��M�.,+W2A����Pƃ&�I�����<������k�Q�F�Չ܃����+Q	�-Dc�-  C���@�����\s|���\�D���#��<b����Iٷ8�
@{?�u@]_���-c��߾�k�+[.s�.���F8�L]��Lm�*�$�:���g�����/�	x���:g�pNC�w��!���m;x(�����|`i�q�L-��/K�7�(y�Ap�	'<��C���U�hz ԰`���_w��z��c����e63���[��ֻ����Cg����R�3©� O4��01�D�	�'!r`"��
'|`z��d�'�X2��k)AۆZ�7M�%^3�0ҕ��W�[�@�Hm�ͤ=8:��G
)���'r�?Y8a6�>��&�3hӗ4��i9�bHyMD{�_��F'ʚ�p�,#]N'!3#M�<�p�[�!<�����]F/.�+���~�&���B/(p3�.��������Y:x��?��?�R-����L��6/�����}����w��w��]pup|3��`�#�UC�������]�]?���r�7^w�u?��mؖ���Z���`.δ�_3RT������""�,N��� 3�"	���`�"5����;8��G� ���^(�DD���0HBl%�S;�o�y�F�'QpU�v���Ԃ��ڥa����L/e-��]bfNhd��cF�﬒�6C���Րy��<����0f#�"N��n�?���h�blX�["��ݳ�<De��#��"��4Ҝ�ZQU|��F�0��*�\�J#(��4c�s���SBXi	b_ð|Eњ����^[��W�����9�_)��P)�}`�S`��a�Cb�F��@ӱ��c�#&��K��}a֥H����0�ȇ���	DEV.��׋�GQp�I�N>}��Z�S�hT�[�tynkV��@�1�`X�x��'�f"��G�&G�G�}a�q,3�y�Y��� n��c�6SӋ��i�Tܹ}d��-�|��
9�T�5V�����~��%!/h.,���L�{�z�p����)*�"#���Uco_e���ﴳ�^P.#�r,��'��C�|i�R9\���/��y����).�t�����9r���vt�Blڻ"�U�V�-�_q�����\m��jw�]*Kʲ��ʹRe���:�Y�m��F�`w��D�L����^lJ؏�b�M�1����bۮÇa�C�#	��� �45p}G`��I8�Yz��hw������݄~^RT�{����z���A�&�b��.<$�㵽�汖^��Iq�:L��q�^�J&Ņ^pmn��Rw���={�_��ѹj��գ٬U�B��ʕ+m��v(��[.OMMM���?���hXD���(կ�Z�y��XU�@nB0�B�8�O�թɃS3��A:z
�%��1��l��@�D������l4�6#͍�M8{U�w�Cwxx�P5W�Uʈ����\��\r���A��I���Be/���1e1G�|��A�7�s�I�����;���T����G��~E����I��dH��yI���H�q���-Pk� Qh��>��#^��"�	��+����ل;Ѓխ�s�/���5�p��"�R�`*VP$�X���^����\}�iʺ�������g.մ;�����Qm��`b��&^"Z�SO=E7r��V��\�ʁ����dwuu��v�Z�mD>��(����!DD�TGFF���l���|��556� ��kX�����;�Þ�f�-�J�b�f������B���X f^�LM��f���l!��آI
+���Mx!��(\� �r��{w���{�l�.�T���tf_o��v��	�j�b]��2�G.���!�i����r� ��H��j�ޟ�v�~ӫ�ٲK��$��1K3UY]�G�nT+��-�c�39k�� �%�X��P�`e+�*�D%��kws��I�W����Gw�?um>g��յC�(�F���y�Bi��RS��HF����!��8������\��Y�S�8��~���s�Ɵ�}�	��N�H����a$4=���y�V���^�
XQ��E�'¨�p$�C�X�HBC����f)o�������#c�4���1�����=��U�D���e�Iq�0K���>՘���Q��3���x8!�@n�baǇ
��׿���^�^P$6�U�W�cʈ��b�G�d-^�ri�z����=��'��㲑3�k���'�
�h����w�����C��A��@R}�Z�/z��jQ��?9a�I�xqku���7���<��hQz٪	7�^�A����w��������,#�l����Ʌ����\��a8ߎ���D�>���C&t��#���� ��B���$"l:͢e���bq�P�A�=6�H
䣯����L�(�鴴L��k͜SD�e�(�pp�����":jӇgխ���)v>-�7���g� �AT$��~�A���W��$�|���lb.9�x���5�/��B��H�
�<t����P��b�F*	{{"]':b�"*!!K4c�w�]�!em1�,��!���]Z�D�d*�����mj�,)��L��T��9���P�y��	���K��#����D{�D�6��/ā�L8x8ƀ��ҥK'�֥!
9�",^r�Yg�q�p<<�O���u��Y�Y��98X@9B�V|���å�F4X��O|]a3�,R�&-Y������HH�d� s��V#�b�v���H 	be���T�Y���Bt$�,�Zԛ�d�!�,^�)���x��=��1;�NA����l�u�]��-Ɩ��fa5r��2۰A¹�$�����p�y���mٲe����f��z�)l���s�=w`` V����A7ba���$)Z.f�	ӿ�ݽlٲ�x�\~kl�^� gsy�3�j.��m��n�"�x��ѩ�U�{Q�m۶�zf�g��'X�J���9�ǈ$;C�n�6����H��%8%f�M�R!��7<�;�n�w&?�%�G�6⺽����������8�`�E��y�`�i��Z��x��͛rnr�Og||<n�o��b>g��lL�f��t�8���B5��Ŧ�5j?pm�{eu�<���y��,�Ҿ�L����		��w��E�����%��ב�*@�%CDa�d3l�W8�<s(���#��8��N![�x�`͑�FM��dK�t�~�`x{ͫe.�F�qY���s�M��8P���3�<s��2���Jj�8d*�M�a�X� #m�dÆ�z|�M�6�zn������>^s8g��-���R	J6�{��S��
�RhN��T� �L}V�������c�'����)�1T,u���%����Jp���1��詧q�5�ಛ���{>��~H��W5�8RKjB�t%���M�ʱ_���6��=��jM����;-�]��O,a�T�p�`�7����@���V�\y�0>K���q��%h?dx�������mv���N{�����&�����6-o�믿����-��r�'^{�2:Q����C��� �=�$^DؐD,I��D%,B�|YŢ37ǌ�xa@��S���?��/��w^��75�방^7�I��|�c������l�6;�W*���#[$�Hk;�^HܜJ���z�H�T����2�ǔ��ZV�z=�i0K6��:i~�brh�#�\��<7V���^�e��)2�x���1,��K� {�����o�Dׅ]M�u֭[7<�������o�袋�gC��2ͻ�{zz���7���X����"A�}��`�?t�Go���5k�\q��Mt;i���:��'l<�T�b�ڵ�>�����zL���V�7�x��Z"N�l:&�Qw�M��0��To�m�T����60U�lz>�+7��@��g�Z�5
yÉM�TC��!- 5'�y,I��Qs�5D��D�־��`)�]u�����\�*��&1<
2��m���q�[�,����n��(H�Q��d7w�6���R���KH��|=�;\�I��2����4���<��P�*A�=����Ғ�4�8��eSp2g� ����V!K! ��J��T�M����@��M��d��_�r� �B5Mj@dc���1�I�e���7�^�蚎�ښ1�.H�*)�NM�2�O$Q� o�N��� �D])'/w�)�5;�!�Q����X��v���}ܟ{�Y0EK�2��k=����5��|��6=�7U���{ǋ��욜<1B�ƒ��'�X���YZ�ZȇFGz����]����B�U���&)��nh���`Ez���﹧^�b!D��<(KU��@,������N��SO��h�0�M"z�i�	�PA���rU��	�LAb�Q�����n_���./F��B�2�w<���{��?��$��O~�Q͗�n�V��O��/,��W�Ǘ{{$E�7��}�I+!J��-���f׬^�����7n��k�g�ux�����t=�l+�2a�98f�Ȗn&�9٨Oy᳛7/<�x�FmMq�H#��|�K�Y9�=�ƪ��Ѣ�m�P'��
f�se�<宆������SV����E�������8������9��612��(`L1n��\�u��ԩ:�벁�쯎�����:�S��<34��XP��(x*��~j�ܽ�/�w�*�+s�:���(z��g�����J��Փ+��޾C�:H�@?)J����9�Wi�N[�S��v���T8th���C�	�|FT	��Pݏ�[�����BKMR�N=@���3'ˁ�p� խ�{�3�h�	j�鉔d�LLv��ʐ{��]J+Y
� �&�|
�{�u�3�UCY�"޼m�֭��P�x₅����`~�e��J�-PE;&�܈X�N�kH�pyC��d�;�S�f��T�i���Q.�uhd̏"7	!cb뎰�aŚ�}}}+%dv��;3$|��Z���==����Ï<��3�{��/|�������ѣH��ĭbL%���*��W��}�fm�yٰW�;��gU.ۺu����>���6��ւb	�ҙ�$/^�ⴱFu�91�mYn��?4l��T||��e��'�&Fg{�r
\�Ν;+Hs��L�c[�����Ԫ�g�y&DP�3�e��f3q]����������vH�V�	, �q⇈����3��ۚh�	^�]�\'�t��R�:�"I8[�2��\ Y%<��qdW�W�m���<�c���@_AǨ�k�ҥ ���u�:9���/Ƀ]��ISR"_�	4/��x^�z�V�ƚA}� �*���=�q:#��~� (K�J*Gtj��������,����˭�˖���v�E4��F@�T#hbI�Ĩ���D��D���iPP净��*u�vYvg���;s����<�{�ٻ�0M��3w�=�}��y���ꀅ�cʗ}���t����C�}�o���O�&�T�\�j,X� �\߅A��p�j&p@$Y@�+rq3e����_��P�9r|xR��m+�r�]��t��Ǭ[{ƙg����k�x_��/�+_#��?�aoo��c�P.g��˛Q�o�T�LWy��(�s������4,
�˼�[�v ��R�D$���;7���,3�������&?��sW��	�BA�Ҵ&�iNb�F#$&
!Q-iI�[y䰛�Q5�L����'PKǑf n#���!�N��f��=ۦ����9sD���9�����3O=w<�gvw�#3%iX#He-`���;��~���<��ޟ����љ�º�8�fLQq<�`�9s~����>b��$�}�]?fI��P�]�[u��|-GtGX�`��T�F�\�,��\6Rw�1D1��FgY>��-�"��XG�R�/��)��ywLK���5��87�*"�����h��o,ዊ�R�KJ8=���0ݒ�_���
q�D��7�R��͗4�}���a��a}/H�7�4b�E'gV�G�[t�W\�� V$���w�����AB� _�響}啟�2���Q��˴6m�d��*��!}�aG|��� ����3���.x���Py {י��瞺��{ɂ��W뵥K��&�`I����z�vbd���!���~��?����ԁ���w��݋/��Q�d qt�2	������,�%��6Y��y�	��`��w��w�y�&s��$#�ܹs��_�[��k�\.�ߏ�n���l'�8�=�zd!�,��S];EsӒ�ԝ扈8h�5��;w��F�tU W\Et���M�(D�xظ���BD�X6����UDp
I,��,�j<��!hlŚ���S��7�:�&�55TA���B�������C�,��EѲe���S�?���֟�~���;w�8tvv�W���[,�����������?�ѹhѢ���j�*{�W�������vb���6�������<�F���pǼ��"�k1�ʫ'�xb�ۈ��C$fWZOKW��Km~e��ի���V�\հ�+.����F�l��j�)�$�aZ��Uf�^��5�8�{��S�l=����Cy�	��7�aɒ%���0\�W�^t��#������������=����s2�<j0�������%.����<::
_	A���D�0/`Ws_�>�g%���rR���BjDDO�ʉG|ea��K��>���p	���][qR6,���1��Ar�"!�D9�OE�	;�(�,73	�4	�5�B�$���5��*FtۆgG�U��K$�	
='� ��Q~�+
��ѱq�ut!�Du�
�m۶r�z�QG�t�رc����x�]FE�X�Z<��#l����c���_�z���?�s�,�w�^=P��� h?�;e��#��
�^�Y����jp�fX�A��@w7/���ZQ�V�5FG��b��4A2a`cJVQ c��h�0Ë�J�%˗�(�	pet]2�ҶpP��{��_���R)�����+�%	^+r#������x�">}T�:T��e�qЊ �!��� �$X�_p<*�ATdG���o���M�]�N�`�R�$�ܧ>["�$�!E��;i�}�D��3�F|��@1���� �(�V<���'��V�`��IM�	�Ϳ�����g���c��V-E�	�!�edw��y��l����rȐd{Qnp�ڵk�����~6o7�I@jđV5횫�=�3�'Mu��W�ȵ��/��(���ry1��y-m�˳�:�ӸI7�-��	˞�)�f�!ZͶ�4y��qMl����-�i���G�y�@ʻ�@>S����+$�
U%\�#<R$�؂���2����瓟�d����w��t[��K����mp�K/�#J	�-�kl���3��4���<��Yg��������5z���k_�����_�l�Ҽ����z�9��u/e^cC�-Oj�7��E%d*��J�s�r�-���b1a�ƈ������֟3=Y-���Dǽ��?�����κ��;�&h��r�:48�����	x�-��s�������c;<»(�쀎`g�?㎻�ٲ�i��L��a��5�RS��2��p���+��Xs��+�Ӽ��W搽n��R9�r�Y/tA�f�eqd��'�fXu���^�n�����N:�T��	��c�Xu�%�~�O?�ܶ����3Q��D1@;	�E3� g����J+�/��/~~�1Ǩ��Z��0��M$+9M��?~�+����3��@�����璪|暯\s�'�A]~��7{�Yh%����g���|ppP`���,6��L�o����+
�
�r�cb�X,���o�4U����2"<����rqt_1M�v���={v��s��e��ڵk�2'������þ����ء�x=���ad�&����'�0E�O���{P�m�yx��
���F��;�Ʈ"��3;JF��&K�v��S{�V�a9����`6�+2��ۼ�U�����a�R$S�?�0�C����Q�0@�h�R4K��x��?�p��S�6�����(���R\O-��jk�eVo��Y�f��]QFw��ݻ��gAA�>�(���]��B7#������o;$���<�}p���5kd?�{�խ^�W���LB�7LWF�iJ1�d&=6��-kv��9�-o+��Nc䍱��/6\$C�E�9�tV�@u(#�R��U���a�FtٱJvc��X�)+�͍;W,\�ܖ-s��V�u]79��1g�<����?r)�	��Qb�wm�W���@La���EK�i08ۖ`5ѝ�d�e�L�\Fȓ����@�l߾��٘B/������Ƒk�2]�bMU��ti��d�<S�
�r[.�����B��i��,���G�cyS`��"�
�is07N�$��;�-q�(&�� �DX
Q�'���`�M
��P��F����#�s;�� 9zjD�(e�k�Z4����	a�LU���'������j�F&Ɗ�D��t5�t�Ri�lSM���;>B&��M ��n.b��j*��:���=CSp�%�
s3Ͽ�U2�E�-9f-���7n/��RCQػ/B����S��2e�eI��#S|��o]�b����_���]������yO9��O?�Z�N��j	������.'����	X����]F�G
�B��{ݒEkO=��_��-��&&+ ,;&��.W���e�V�����ŵ�����
r�p���]���w��yKΊ��݋���@GKc0�szgê�cނ�p���m�1~$��v<f�-�YĮN۲�Ce!��cX/MKXI��P2��R"|\I䆫��|��T˰F|U�nb"�>7���2+��'��"����`�~^<��u[R�4'Vh��s���m���alY���3m��V2lP{�_C�����W1J�J!e�)K,4�`�S���dD�7��m�}��{m�FN�<�-N8f���{�o}[�_��\w�_~�3�ᠨ�\$vpwܒ*c���PA�� YC�DO�30ͪ�2�A�0�a`o}�)�c�ٟ�ٿ~���pb���g���{�a>w*ȱ��1��ʊ��
X���4�&1!#YR)�1��U�K`i�&2�k�j�s�M4����m�ݖ�	xX�5-�4����KM
c0ix�"�Ӹ~H� ��3�	�LY�I&�:P>��e��R����(Ln�`D
&�V�64Q�3K����Kϼk��aL5ֆ�ǡg�����������^���yO�&i�c�rx��\�N��᧗�X1��U�(��_\x-�Ș�nB��O��n������_�fPݸ��^���7����n'?��{Y�x��ZjjF@:~���N_OqD�r��L��������۶n���]�BOtR}�C=�a�棎Z�!2�z%w����9��;Z��*����w�&k?y���?�q(��U��D�@�P|���\
��M��Iؕ��C%����Ɠ�<Wf!7�Xμ���7�k4�E��*b�t�Y5NB+�����'�<��S�MO;���|w�56Bl���ݻb�	�Z��|�C=k!6xߛo���s�ㆎ"+���p�g>��o���|�;�w��ʄ�-�+����>��O|�a �s�9w�~;�o�z�?��������r����?M�d�����J�\s�_|���c��~�=w����/�������U7Bĝ[�f��~��bgt833z�|�rtC=��m���?p�����X&��&U������ɝ;wzDXTr-pծ���Ɏ���;�#=w�\)���%�W��u���#8kZcc��X�M$S�E.M��������N���痧��I��E�x�:�˾�.���LĈ��W*��!p�\�H���P�D�ԪV����?��O���:�m۶�~akww{�Čh�V��Dh,Eɪ��}��W�K�S�9��TX�`~�%E����j�@�XC,���z
�ӓ�;�ƍ���Pl �#��k٩�"�n�vi��ou��P.O���s�/� ��H�%SG�pM�C�k�
<`<�N�biٲeB�
�mCCCm~�q������Y���䆚��H�K�'��H�8x�	K#��J�FR(Z�6663���#���8d)^�����e�[`�W���@l#��c���(�i��`J�z#y�M.�<$V"�iy��EpgMs�sE�I���O>u`�(酠,B�f�aޱ�� J�?�e�A����Q����W��yw�ULc�\s�(�j��w����-j�T��ױ�Rj~�uZ�תMSp�|�2�U���@��0��[;Hy.�_"��ް�7#۞?���/]���X	�y��6j��-�QWR��xV+�� Eq�G�r* ������x���[7��.Z�x�ڵc�c���/_��##��6X�����(��򦉋�pD�������G���wx�8[�%�
;����BOO���8�<�_�64\lcL�*I�� �8�*�"h�R�<{v8Q��:-��'Į?�����~��b���E���ݛ��BM��(J����D�\���<Y�.s~�Aip�T��D��^��
��M�|u�[`wB���^��vx�(�1�q[���>.4�X@���"w�`�3af"k&�f|��8��u��|�9@�޺u���s�g�x��s_�ɓ�0��|��\v�e�eGR�:���M<�
a'"^�,?���ib�$6i��MѴ�}�k��w�P������`F����S���L]�~p�E]����1�2B�e�Q��zk?H���f���<��t�ҴU���l�`d��O��4��ɇM�-�td���"g����&��"-�Z�#,
�.�4������,� ��{J��Ї}�q�?kVf���~�z�+AU ���bk.o��D �r3?�	��� ou�x����>[��^(�8C�-���+�\p�%��{������;��o�D2��p���w��boB_+�CuB�z����:�Bl�u�Yw���vv^�2���O,���wƻ�n�2�MΓ���}��[���"t��顢�"	��%G%������?��s��N��~����?�ĕ�o1G<3���n���f5׾����Z��[K
Y�x�_!�k6R7��I�k.�����E�Y���#1P�H� �{�Y����]~���o>����(� �Ԑ����Ã�����s�6o�Y� Q�BAY�-����˒'�UE���>?�m��w>��_�ڜ����vQ�Ì,f=<��?�Ǡ#~�د���%�:��O������?�G'�=�C��㥜"���_^s��r����\���]��̇�nt����ɦw���9'�Cn�)+�hf���)+fC���V�!���	�,qՇ�,4U'|aX��n� cD
��Z�j#�d�2	�J'�k��#誐W	�T�v;G��)�3bfH	j`��&GǺr���.��������ҋ�[����H���*�g̃�m���lV�]�ި �3��~�)$�x�S�=mRA^�`v�73�nkl���m�,
�w���z�y�$��p|�)�#�PxD��@ܹ����FU�@F�<5mUk�,N�(E�橩���TSw����'4��SӲpQE�<�<R�ٝ{�z��ݍ�q8t���������|~룏P���<��*�{�>��^0�m\قa��=[fh}����2A��x���;7
��&���5T�?p�����u�mȽ�n�>C�kjvi���"��%#�&"F�sh�+u3[��a�Q)��|r�VAF�΢(���v�/�FJ!ӮD�S�w)�x���J~��w6�uY53��y�aM�!��dwF�w
cCe�#�r���^8��W;
X�m+r/_���������/4�"0L�&�����<���`%[�Fh���<"[���TTl�Q�!�h��M�yLΙ2X��""���Q4CIƎJ�
0�fL���Q��7�U0�	�����Xш7gAT�+Ӂ�P J&$i庾��sM��,�r��AF�S���]AY$�Yq�� !�|�Lj&9�՘ncZA�ٵ񡝛#�eb�ݘGBM���;�T��r�fB:�6,��RCX�!�&O������Ji4,g���X4����ʆ`�I91���JB�}��	z>��h�ϝ��Ý##��?��,9r5Ĳ������eoy�0�i�ds�#2�
1fKt7���cA��S�*�%s>u�g����}��7�|��Bq���^��O_\���.�H�c���[lF'F�U��mXW�?�����t��e�����}]��_�G��;��J���F'ػ�962R��)5s��:Fvr��Aq��p��Ș�*��ٖmf�F�F�y�A�k��+(r_�Q�쁁��n����,��a,��3H�t#냈
R�t�����dp�@~�1�Ɗ��C��f B�!D��iĪ-Z�H���eI���.����_�mG�b'�a�d1 �:'� �B�Ÿ9�"5A�a�<Y,�;
s�8�]�����X���	��,"��Yk�d��e���#�An6�q�BTZa/!�?{�+@��!�y��3�FY"���]AJ)�xWs������n�2n��*�u�g�
ud|���4Ԉ
BJ��gI��KDO���0�R�H�y���X�RF,����v�$`)��)�K}/��8��&D"J��	L�$a� iŸ�JA��=�ɢ�%�@�q,60!���:��ʕ6���0T��6#w(����t.! Q�LI��vR�^|ه/��?旊|���A!'^�n{�-�����V�m�gQ�y�������s/�a�9WߥW�ɥW|��#����̙�@���h���aډ'�޴����D��꒦�y�#ઠ�lc,�TZ3n���1K�fˮ���[能�|-�suU`s��?��?�%��n7�$	�>���ر��s�����۲e��G�#R��,[�졇z��eǶ���Q2i^�g��]�[�{�w^|����u�<���F��k�5_�K��V���ȵ"�~N�w����Ɨ����nϳ�Lv	��2��ԧ^�v�ҥhFJ�G�ˢp #�q��O�K�,a�m�Q=^BɕW`��~;l$�^{��ի1�!�d���r���믿�#��7��ͫ��d�Pز}{(��֎㊪�q��N����O��Ы�a�=mٲ��|R����K�D뢠���f?���!�vԂAģ�z.{�@�ĩj�K���Ta��Ĭ����Y,��@Ψ�c�{��-�-�еl!��-[����=g�p�=�إ�c��ӣL�7�u�5��p;3.�c��&���m�b�6%�����Y�Q�ݭ[�����e%�$�C���^��y΂�b�3��&���������e�����ؑ˧h���2�]8�5�����ix�B;b6Z�ǂ)_��@>{+p�&$�nFV�����h9\�$cg0È)O�� ���cUa޲��䊶�l��U8�*�e�a�yI�F��4��dJ��s/n�60Ʊz`<����s��eQU��r��R=0r(Ik?��H��$�λְ�����-�f�sn	�����,j2d^�̯�A�p��vwuu����>��ώ�P� p��^8$����!/������*qW\���B�'pR�U.`�����:���ݱ�A����$�,���8h����FI��SdWޤ��rJ
O��I	2'�NT��N�"�x��*!���ͥ��d�f{F��EE:��1�S�����v>p�:!�3�Q�������	h��p�-\&���D�c[H��^gh�.þE�;�ޅ|I���$�<��B�̣&1D��:��xs�T8���_���}``�+�.�B{^|	���&''Gǧ^~��=���ŋV���>pՀZ��tt)k ~l�
��DzU�­�9�Ї�ScO=�T0<�}�vɪwvvFB�j4�lV�={6����(,g�I$��`f8m1�0������5,xA��ֆ$]px�	KZ�H�๮� U�_w�C4|}a���%bLj ��;��L9O�IN�l�U�痈4xm-�vw�a������S��(H�d��'�0!Qxa�\~�'�n������x3R�%������݉���}�d�''�,�4%�rB:�lF�c���#j��T���I��7���f5�&�s�"f����@e�jEԴ8����v���*r�������Ō�]"��2I�+�n�gz2k��Q)��'��ͭ���;�t�VV���	b�{7�`��}�ן{�����;���+�IeU��y��Ю�G�2QrUS��$�O?���~�+.�����/X�`yJ�H!����@�9������C�E���/��3�=u�w������xoL�^�&�Oci�k bX�O,a�MV7o3Dvԉ�y�)Zz,�dEEU���O>񔧟|��޴n;���Y3�"� ��A��3"���6_İS��)6l���<'�e��ZUL�PcCC�o_ۑ�7��bG�Iq,�4U!6�04��M/o|��wvt�����歞͎Zs��e+K�w��9բ_��^�
f`Y��KP��U���h1$�%�����*�$��qbWI�iYDx{�%<.Ք��4B�T�j����#z����^����/v�-�{��<ugX�VF'�P�u�4����nê(���r�n��*��<eL�*�\��jvhy�T͕��iD�¤��-��=5%�!���s�ݹb��hn����옞�4�=�&�"k�)�YN�G8�+��E�������r�R���,�?BȊ,!��C�5�$�3��֭|CI���:�H����%i���%��@� �UmM5?"7?
BŪ#���*5�c�1�HD�l�Ps�a��i`d`YJ���A��JQT�emwh�*6���$�R��+H�"��%�EW%Eu�T��a�Ǯ]��_�%����-%�Mv,�����f=�Aۊ�7P׈�wc�}!�U�*H�����2Y��źA=����H!�ަ���e1�V@��zC%)_�ł5�p<(���<="�V�>"���+��!a3���2�Я,bUO���Qdn�dR�TT2�pYb�a�$�v�j���
�#�Z$��v,ɦ
;�e	~L��N�'v��,ŭ;}�$�	<x�π@W����h&�G�N�ao��X�b�':c��*Q\�T�+�`(Ö����J'B&���Y�b�a#�"�����>A�6VDHL|,̦Q)��
F$����@�i�8n�a!����>8ީ"K�\�^�3�7��x9+'a�Styll1�e!��5�-+��.�TB��b{.[Gg�A�x�8�8F�^0�����Eh�P���u2�(�d�/tъ���5�6+�L�Ĕ0��6^�bIfXu�ݏ���x��f�Q�h�:���Dq,��;Ŭ�3;3ktl���OLM�1����moÈU>�'�^��@2��\��Z��4*��fs�����!	�#�UX���-B����,#���5U3Q���q}�H�hQEĩ�j�����.)�GE\`�,�y�'�&N����Q��a����
�wuM�:)�_�&�i�)��	$х�B怞Ĭ��$��� Na�w<_v�\`���Q�"�P%QFY��A�D���w��41�G,�}�n�%�����9��%�[��ɡ��~��+�����>J���[���Ay���/�\���}S��S��~�1=-�&Z?O��_�Ef|�����\���<l�ޱuT[�VW0d!j����4����$�E:������>?��qb��Y���M��ߡ�M�k�E�rܶm�p�gLW�l��t��,��1��-_���矎)AA Q<�.]�����K.�����;�<^��A`$��Jo��H{*��ٳg{�>����dOWwò9B��9f,��1�+��xE�O�_|�h�"$ImA8S�`?)hL�#��+���I��X�qƁ�gW]y��w�y���99�q��5.����A�dΜ9�I��A}N�Q�����N�n����v�o6�;�B{���x����]w� l�޽^�.��"xZ]�m�~a����y�;�l��ו�	������	�A�9����!RUmq�^�LSGN�ݻw?��c��8�l[_��1T�{d�W�H�9Q���޽���K/����EF�J&�,ҵ)��n��6�q�����W�ήͯ]��2]%ڕ)���J�ҳ�>����͛c����$���0T�HƔ7@� ��w�.wvv�|�	������|�����H��/Q���	uJW)��٘ɬ�j`����F0N�f͂Q����M��RD8�x���7\ǂw��VSC{b�:jx�7%(`|����X,��n?V�f)T�wMI�1��q��I�B/��z��G�@_;yJ�"�}n��N�w�ÿ��������[$Q��l�*0�"�������ps f�.�Y����(FXwp��8�p���o�������;>>ɳR𳗘;1O���`"����s1��sh>1DSF��)��yx�j�b�M`,LĄ���(��>U��N��������t�[Wq�V��4t*�K-��د6Y1��$��6L�����F�H�R��]�JB����1+r6i_��l�D}����˲e��C�v�T��UŘK#�O��S7���{ّo;	�m�b�1U����]�ɰ�ȵ1�GT75\S�8����H9�2�1v�e����߲eKi�6�`ilݺ��_��A��;�_x���q-��;|>�p��� ��5�#;�bL�5*��������F_����x�2������o��s�Y��j0�v��Z�1˪�J�<,I�L�J�l��?Utstt\$�(�;|�� 	+�F�x.h�:�:C%�;������B��
\��-(z�����B�
(L��Q�pye$�TgM�L#O[�2PӰ�0�0!{�쁩9��`w ���4�Ð����n|�P��%�K/{����[���9-fw��Bߐ/aa�Q��M��?�[,�����x�äz���}�46�����ь��o|̸N�Z�
�?$W�3ƪ�yf\-u�fl@�k%-�o����z�x��:3/�?k�'�7���u�`[x���;"-_�0�Ø�B� Ǫ_�+���j��Ej�%*���`�K���Z�����߸�g��,|���	�C!���(�'P��K���68*9��<p34�t�`���H!����&A�$ϏX�"��d��%��<�P�l��}�;��c1�G�J��O|����0���+.��d�b�<�T���˩�!"_147��u���+���6̞�Lʹ�-��J���ߙ"V��"�ظ�����F	
�ׂ�a���C�٧?􉫮����^�^�˩��G�K��>{�?/��<���N=�W|�?���c	�	��Ĉ��(�Q���F���']�X,sE$$�QD�Ghx�H��m,p����v�9C�Z��H��ZT��������p�L��aw-X���D*��.�|���ic/��;�{�66U�#��� |E��s`yį��
�2�c��,�k����2e�9��h���2:6�m���P=��$�C]3�+�Z��+ _[���r]�ԥ�l6?00�<m0��j��:r�x���1�`�IDL�}�
�L���u�� ���]WS��u�X3�@�#Q!��M�6�P�P�F��o*	�颡��]¤�֟#ȯ�U�8��+Mm7LH�2�\������肬���2V0�Ɓ����n�h���,ɪ��Y&(���?��<���nE�����Y6��8�l	���M&�Dl�f�=�u�Ok�����$���Z&�5�J�;5Xh�n	�TD��o�Q��A~A>c�`��"x�熮s�?�R�f3�/��GT�U]Ɛa�=���B,i�v����!���t���?��,U�p�XVs�-��ՠ����C�wA�D$����V�"��}�.hw���]�dEbd�c�Ɖ�@�1j�Q�[|�b��Y��@��$�5l��ӄp���24�E4�c�P^P�Y���TC+�	e�L�r�`"���,�:����N��bσ�"ɂ�N�HI-��s�A���q���9��䌦R{SEIW������&��s|T�CuXS����$k2u0�9������ζ�^��}�~0�ݬ�L����P�t2?�Ր���8�����s��1���/
���]��STmN��cC��L�jqV"�{a�����Bg�+�ڐU<i�$�Z]b���
@P3ȅT�S9���bA�h�1̷@�\߃��+�
���� ��Tؤ$��J�vHy�ᜂ�"e�mpF�r(Z�*�t�D�CF��T�<U)���Xc(��D���8����PT��$�*�I6�kPƾ̉���-�?f1��FҕI������3����1�;���C�w�W�ӛ6�X<@�т�gT����rWo��ࠦco��0  !��z-����j�k�h��s�k��09Ո�LH�㫃?����I�|������MO)�I�_� �Ul��0��m�c�����-��f�%�p��~7zM���ْڗ��x}8֐7i~x�m��[_�0w"/Ki:�����.�<^�j-,X���&	-���\�sF�.!��~���n��|-�,�ݰa�G�+
N���PA������Ue�
�=����o��V~j¯g�������������]���q2+�#����H�V��`��!&��M��T1��b)#{�1�B<��P��
o��n,e��ښY�'�#mM�i�#֬z�'DaF�~盜A��GF}��/Oq;��"��~���؆����V�\��$�U)iW m���t�>�~�;�����9�p�=X�ftz>�G�2֮]{�������ήm�L6<LQ{���$>��:�q�����(;P�.�o_��\�q !��]��{�-;�`��͞=�P,0�����˕Je��.��0�`dr�j"S�v4�ES�8����9������p���#�8"�E�prl����}���3:�=91+Rp߅'=BS�-d����u���Ve���	�Ɖ��r@`"�}�(�B�d%�i'	<��f���:�0T�s�B$3��������0vH�r�W8MV1��s�z�DN�:��,H�n�S�\�NLL������eLDg�d�8\'�~��l!F�
E+y^(����WU�2�'%�[���b�|�&C'�[����C����ä?-fQ�/j��D� �C&�ىÄ4��w������ �#Lv{{���;88X��*OOwuu*2���2��"�.�A�g�X������냙��;��f�}�?��i�gͅ��!f�$�w�LiTd���]]]S�[^��xhc9����a�������ྯ����t�
�e���'�|��=ۇ�����ϋ�2u1�h茛l<)���>���"7�r>�\�8�;���f��+�{6�Ɂ?ɑ<�Z�LV\�+-� �4��'؞�����}lZ��H�,Jjjrcצ�]x�UQ:k�*��ܿj�B����L����y��׭[�p�8�4�9m%��$�1�����;�{;�k�a m,r�^F�s�L,k��w�׮]�c#��A�{��U�Vmްfg��!�K>�Q���XOOO�^�}�
�)L���#�P�*�.?��ӵ=#p=�Aq�����E[�
A$V�
�z8�W[����3�3��h��köv��MEf>����Y�ŋc���0|n=��D�.j�	�by����j��l��C툲�R��ЂWI�'Y��"ѫ�'�!@��V�AaQ}M���ep_Q;�H�ӆ��!3�(���n��������r��"�)C����7��m*���z�h{��^w��A�����\a���q��g��w�$���+���]I�Z��4�k�[{=?hg�{�:�)��}��i!�M~=~]������<U˯�[�xL����y�kzǒ��oF_˱mMfG��������,1�mr�n���7�Ĩ#v�HRB�K/��������|�}�U29'bvc!Q�롨7�IN!x�'������W�Y�8��?^SF����؏`D���/\r����ކ���Gznx�%�\���V��rCC#k�9���$YV|��v�M߹�}�.��S&	L�C�.��$z�:l>��2�j��ԣ{��\��s�\�MJ`<��+/����is�ɚNy�X%f�[n����?v�������P�%?�m��E�Ų�����!�
Ѫe���b&�DO��b>�m�!��d2��gO4�>��ǖ�[pE�p�J����l!�^`Ŝ:��h�`>�ERY� �NP���V"Mu��� ��( d�Ю�V��zSy]э0l'4M�[~X%��l����cKu_�◶��OW��T��ftxv��f���,�e�l� �af�PF�*�(�1|p9�����E�/+�`�`�O���)(�Vr""gT%7
)����]Eq�R��*��<�v
|E�;4�o�ߨl7�J�O��Aj�)���C5�P�*y�n6�)� ��(�OP�`.����e���ed%o}]��1��B\Y_�س�%̑��( �p�hƒ�<�EL!� I�/���D�m�`Vd�R�,�dQ�bS�C�2�F�A��U(q���Z�}��¾-N���E�(�EIN/�]PJ�Z�=3�Ba�b�t_�s�G�2��+VFY��|0ysV}"��,L��H�%Yڱj�@�V��n �<"̛( �U�a2H�E�8g�,�L��U�@�GULpƐr���b��.L���A�Kv@Y���NS���˛�TݹE�]g�Få��e.�Q ݋�~T�"��"�qDQ��aa^�r�	!2W����È�B� ��$!��M�ḥJ_&�w,�zH��l�P��v�p$zt�|�y��,%��F��Ƞt7%��� cz1$�r|H�.��צ+���6'��%��R�*�d�iL��͒`t)�axe�ڨ/�}dϒ�u�'�J�f�h�39=#d�F�
a��n�;��!r)*���UC�4���]���l�1^�՝����4J�!���nU�c��^�[�0�s�*f�,��:V�V���\&?�|��S���428p����q�r�֭����o�(�2f5�&�#���^�.2FX�tMS������ T0ܞ��-K�ih�*ǡ����A��Ƃ��`�y�넞��=���5BD�i@
(B�PV�T����	so�
L9f��Zy����	-��I�!$3�}��ϖ�X�XS�Э�!C0��0�E�#`���l_u�q Y�7����ʠ����$6:1��{�6W2�˂[3-�3���LHx$y����nF�H�������a�s����׭w�rӯ��`Igl�5���ؔ	g�����e���u(�@�&���۵���st��������>�52B��*0��:�Z��3��h�d>ј3qf������a_v�w��boB_�W�0|��`���۸�{eجg}���w����qpp�ڵkA�0
Z$QJ�~���}�����o}��Dh2�5�f��br�}���.��3Ϭ\��Xs�y���@�����H�dB�Z�l<�O��#�<2��9��d��/W��B�o+(��#�h�|�H��=�]_��� ��K�EJRh�,���{�=q�]w�]�LB��n��3$�2��7��Y�����D��_�җ����[n���.��AZ]�%�13�B��^w�w<ڇ�۲eo��hfV}�qؐ[LJ���M�Ώ!(If����*��)�\D����b]Cz.�p`�G�n*Y�:�ꂃ
x�.���Q#��f�<*�@���̤��A�j��կ�h��	�z��.N�^���A���<��`  ��IDATv�9�J��^a�\.'~�ہ0�f�DJҒ-��1��sCP��b�K�
~6�,O#�[�J��5Sg��=��9I��݆UÀ��ٰL&���,��W_��0�1�MO���>3��p����� �B�p��'_t�h�؍����\�.��)��D>�m<<K�Ab�>�SN:�$���o��a��41��ϗ(�Q����4;�i0�ߤ���Q���	���6��ay%���h��E*`ڂ�[� g-Č_���SO������e�������Um�;�jšv|"�0�����Hi4^�b��� ���ha�ا[/����'�L�ŌD{� s1]���0�i���4�Wb��Q��}f��c����[������a"2�"2�G�i)����m�Pc�ECɨ�C594(_V��=``%�رc�x��m��͛�!<&�!޿W�u?N�Pp!�`�Ot�I�><���A����Q��d2�>�d��J��_檒Ã�������=@3��������ɫ�<�y�����F���fU�m���/_�·I���ݕ5�����Jx)������̦Mp��b��sX�p��ŋ��2�o~�K�,���%��T뵹s�v�w�J%-D?!hأ�����g�p����F%��5)�S�VFF�JX�U$Ds�f���X(�9�0A�I�OFG�z��e�0;v�󧧬��BOO����:](a�nݺuz��"�F�_*	c�ש���G��f��҆W�ec"a����ү%�:K��H��ߤ�,"۬է9)|���X�! 2mVE
�8B�oz�=���al�������M7�T*O�Z�jnL��-/���Ț���~L��L����z~�K�M�����Q'x�M�����3�F<;��t�њ����d��r�L�!��O�[��ݔ�+Nh��k	IPo�I#P9cf��,�H����z<��v��|-_T\?ʈκ#�(��#����5_B�{P#ѓ$�J�v<����c��	���L.Z�Ǯ[yک�~�+��|�*Ɇ��%!�bkO`y/�{,����!LdKG��wZ�+W[0�c��Fxiܼ�I�=5kB��)�����6�S�D9K�be���r��=֔o~M��zf$P�4��cu���^�G��\t�����o��u�.[��=���#�+�A���'P߷�x5�z.l*p]CS|4;�P�5I0�g/v��R��lP�}^t�uu�u�;���׬Y#�eȐd��ܫ�?z��B�CW|T�5-�4Ч?��o�۷��C؊�8�9l؞j�!�V㈅+:;;|r�!"t`�yӦM���}��k���>}�9� vV���͔��ppU�D��+j�ϣ�Cw��ł�O=y�;[�j�vkYT���XV5�#|=��S%�,tbD�&z�Qˢ�<�C��<��\C���&ǒ/i��9!�1�O����~"L�B�r�K��!��}�J�A	4B� ���+J煘��C����K�"�Jڒ�u��d��
�O{�I��G�\����-&��$,���R�1U�9^`�.҈խr94Bf(Qu���:��9XBI�l�Tld=���*SSh�)���+���ɺ����5��2�l�����Ƈ'^o��d�����y�fq�D�EX�]��L@V݈w�����4�@ௐB3����dR�Y+��_aؑ��,�-��S%Q�]I�v�	���
�����Tww��c�j���dY55��ՊS�	�igU�?�4J��	���� ���5��}�G�@7!o�( �`c�/>=&����c��ĭ�=�?g	�_	}Sdu�S���V�8�Z������W\<�b�C�;'��b"xEƈJU �Ey�<�Hn"�'U�d��,YHCA9j�z���" �+�?H8�*����A�r�b�ٷmX*��n���`=-��G��*X=+�L%P�_,��3u��!�Nl'�=�PTI�������WH�Őx��db
3Lt$�Tz��ո���A�81`�]Js�!�rOG��(��J���li�T��hxbx۫��4e����P��	�P5����c�����C��w("r���/s���%�?�b*{j���3,��X
��}f��]�C�f�j��a��^���%�mp[��FG�����6�U�PA��c��y�� �k5��
>˚ ����S#�w�8�(���c;�Sk�*GP�:�e$�f]�q,�4P>՚�M�z�؎�\0�~�Ǭ���F!���+�{9ݰ$�
m��S�c��	F�,�:J/������x[Imd�F��g��hr*��P�H-ݚ,�0�f3����d]5_Gi9���NW���[w�v`O�jv;��e��ᅗ�l�h�uvwM��ʵ�@հb�� 2�Y
�U��QʛQ�*��dI$�M\����I��C��Q�y�_�5���Dc3�!�b�;'���^xF�Ih�n��<��hӘ�Вs��u)��r�.��=#��z&����~�A��@����$�x_��o�>�����9�t�����\p����׾��=o�����A��4LhL�*��Q�����������r���^{-��:���3ѽ�;�wÌ��㪫��z��g'Xj2��,Ys�3^���NM���KńT��s��&�%�+W:Q����]�w���)�����N��ƇTM�4>��[֝t��_<�������`Y��fՑ�����1�AÇ�����C ���OHb\A�уG���N9�c�9���~�-�~����g���s���7�}�;�ik������}�����-7���������b�����K/��n������s�Y���߹s�3~�iʂ*��&u��,���:֪��=��p�� S	5�]��^Dy�O�8��;�yF��kP��o$*ȯŨ}�$�3�i
!���0���ePc+�
2V�a�A��y�Z��X�������x.r(��mP�ϖHM�w�$�?�5�1�s,b�4�A0�����>'�uq��$.H�"�X�E�a|r
��#�1Ry�䌸ef�����X��-qʐF�`�hx�VH6��<�L�*�޽��;費���/�<~������l)�$��r�'0��V��,� #>��]C���[_���51��W��8z��&��?��n@v���1Y�X3i���$�&�¡Da9���֭[�/�����4������Y�?���Z�ׄ���C1����}�!����PN����4�===0���|�/�PѯQ� pP�4��C�gKsti�C6���n�s���ر�g�Y�z�q�楗^*�Jy;��ܹs���P�=	 h�T�"���ܡ�DvSc+n�[��?�\U+I��\.7K��,P[�R����)��}%���8E,{Bh@gգ��j���e�q�w/ʪ(����v���%WeS�Iy���##+TK,$��ͨW�q���ĄD�7�8����Qx�|�76�m۶'�%�08��w�a�aO�n^WW3�ۇDqӦM�,���fϞm���	4ȃ���jx�?�����Ν;9�0x\y��:;;����CCC/=�������0h�yݽ��1.@���yࣚr���<�pbYL���@����"A�Z������;L
jH�l�st���]]�QG���a�'Q��B�/���}j�>8886Q�E�$Ć�Q��FXdʭ�V91Q�M��)*G� 1���̵:��r�J	R������l�Z/��65��c�U�斧'�Awq|HX�N>��O~i�G}v�9k֬y�)U4��_E�)�R��$v7<~��7v�!���3�A���P&rE�
�[�~���Z�\��>�o�x�_�w_h��7��0���.��?<����Х�|�oox��_���$�V���Nk
��F]�U��3g��dL�՞�9�?����	ݩN)�^��l��lv��@����>h��^t�����q��b7�3n�qe�1�� Q���g��/Ěk>1()��U��cxR���� G �k�&S�%9�(CB�UdBF�������0�G�S�e�����9��_?��	'� �s���f�TҊ������5�\V	gsXO�ڦ�q�iNW�����9~=�[�%��uG������㌳~|�]��U�h�OML`�8?��k/��j�l�e���_��l����/����uMw"�b�D`��:2;�E�]���������$�e��Ûy��?��GT	�6��|I���$S�x�=k��
͞����A���qn���j򎬘�"���(�J����P��F/�}+�b� c�Z(2�jx�M��)���92R���.���.�kb���$.3�JT�,���P"��=lT��bGJ�9X(0�^���h�n�>���&M�y4��e�;XZ�L�����	0�}ѧZ\*��"Ɖw�x���z�Zg���Ԍ��j�nXל�&��xr�E��7F�����޺M�KZ�k����>4y}�}�?˱:�{�B��1��q�Fmv/�z��4<F�!��F��B.��h���C̵T]�(]�e�Ij��íVm�Ȯ]�f͙���񎁁9]0b��Ex��q���8��>��H=�޳�tq�KS��U4iYKR�x����?;�۽P ;]���d龻��Ϟx�����64��<3�t������={L�UJ���xY����xe�R�blLb0g��4��kV������3֏��6?2 �"�2���"8.�9�lN�B�AavD2�#LV�>p��9��S��?��Ԭ_��Ffm?'�b5i]S¿��iX8{��	K��W�j���t�*(:�5��Ԗ��y�j��<����(�,�����1.`[u����3A��n6�A{��N�ӄoU]kj|bʱ�����/Rw�&�vE��]�:Ѥ�P"�����-/�P�	�Gf�IC��K�3���V�;�13Ө!��$�UK޵n�t����)�_,���+�>�⣏=���LP�{L�Ү�^L���E��u������p�Q��m��s����X�v�ik׮�j��B��W^��Dެ���#���Z�����/e�#��)�xǻ�]� G���~��������L��{ug?��/�n�ޜ9s2�<���*��d3�e�FN��_vGW'H�G��	�"/�ᖰM��3wkp�.�N��9[����`��Z9�ǧ&�$PAz>5�5��[��������iwL��4t�bNdP�:�[�"�-%i�4nd����k�1��]��%'Z���!�q�oZ�2�����i��ǺPQ�s�|&�Q�m����Us��@nh�7U�]wW.\��;7o������_����g�fs/n�619U�*�F��;������{QJ�0� fӂ�O��7��F���z;�Z�����a��_��p����1,���A��:��8�m:��I�݌J�^���{��1��<��;%>a3}���ϣ>��<�t�V���u�,Y���?���{p���<�_��zz�9gz�f�%$!
	0�"�fn���M��ט�v�8����c�q����`z�MHB��v�̜���u���߿��ь$$�,�����Z�����W�����;�s��z�ɳnGo������q�S(ڄZ��?�=�o}��>�1�qiOj�|�#����׼
�Ū�q�)]WIE��3��L1�o��
�b���Υ_"�n���r��J�]d%Xwi�f ��d����p��ap1��ݸm�,�!(D�,K>��)kq��*('S��X����ϓ���W1��7�%���9|�m�H+0m#�CZ|o{��~�?�'�:�d�k�}hנ0�f��T�>��Bc�]��C�?�������gBГ����?��C�����^JĚ����/|urr1P�a��-�yBE��n8ҕ�
u˖-�++�}�>��OТo�ݿ���}�;j���P�-��R�00U�۶.G��f�K�Y]����6L0��t�Ɨ��*��C�H"��ÕmA�$� ��X�(%�#.f���R�.��e�������ɵ�lns,g2C2U&��no+v �m��]�Δ�@2
ߍ�ujU�2i��p�m��Bj5�II���\n<uu��Dn���P�4��h��C�B.���n��0s�96�@�l�aNy�R�i����Ɇ�������tQ�9r���J\�P�
2w�	Vs��$&3ځ%B75��w�]���z8�/(�)Q�Ϟ={aj�&��B�/R��<}�`�jI��a������q��~l�
��B�42�Qĩ� Ҷ�T+744	D����e�h�("�z{{����,q���u=T6��H�fY.�1}D�lQ8$V&,�V	9�]�)քL ��d�yy �l%p��j�X�3�pV�>)�$Se���RZf��������>��֫���Tw�scp�ҖӾ��'�(ȥG?G����T�']�kA@m���cǎm���p���D�4g�ע�X�"urƒ٬�R�*�Fd`�B&	j���lLBt��:����٢k��FigiO ���S\E��@n.t�=�����;[Yu�zh�X$�=u��׿�u�Z��U��:�&H��W��.GO�FGG]ۢ�EM�kh:�S.\���Z�a��ڲc�����X}h���(�~;x� =����Ǐ_s��t����������O��nF�(ԩk�d�v�V��2!�d��p��LE��l����K��Ũ�G[^^��˓~+�$L�����2�3��Ş[�R|�;��D�va	�A+����ga�`�ҿM�V� :����ȼ�t��D/@��=�ImX�1[�۽��Z���!N{m�E*q�ߔ���5�{�:r�,��$͸4�_⃤�<p��}w�}wsq�[���|e���5Ф���H�ޭ�M��f�&�殑dtOG����s|��Z��%)M�Re�q;�|����#����`���c��w���Z�N�/"�E�9��[^��5I6���ip�DC�&/���������K�=B��4��8��H���8&$�#]~Ӗ���ۿ�o~��~5G۪
Viځ�Y:\%��H(��o������$�;�B�i�U��K�FB&ٷ�oրI��@Z#C;� B�3��T�D�����L�D���JoHQ+խ.�ckɟ����4aL�'U�0���.����/D&WF��7H��w�Ma��Xc�,�$f�V�X� ��2�;������o�9�4��c:S�Ic��ˬ<�o��B(bIV���l+�����w���=��CL���p�D
�*q�w4b/��M��9\h)�!�"p5��]���Ї?��p�|w+Jb��Q�dQ܇��4
��@z��x�f�G���ɂ<)��BR�J4����.�p���c2-��s9��I�d�R�)�<5qr���[6��]ǐ��4�r���l�D�*�)ƈ�F���Z3A�F�6�f�i%a��05�5|;���y�'�Ch��ud.�����Z���/	]��xU�?�ւ��-1��)p�6��{G�iU��qE�Ƀ�@gN� 9~Ԏ�Rؖ�q��fZJ����L�������EO����[�u�a�&�4g�o��K0@h�?Vp�u����4e�PC%�=�#g'�Mp�;��k������-�����W"m��PQR[^���S*(ȴ`�~0Sg�m��q|R�K���f�����^���ך���_ ���W.//ӈ!��)n�lp�Jp�v���Sy���m�Q��Gē4�5]�s.�������ԩSMf�W�����9�0M}���|tqq�_��篾����?������5���J��a;�n:�K�e����e�ʂ&��P��G@W'_����vi�D��9߮-�<��Q7��k5RB��]X���-��5�Lپc�k~��h�fΜ�&ap�����'�=y����µ��w��h\[^E�[W�͚����m�p� i�f��|zR��"�nʸ\S�	�UP�kj� sT	�~�� s��i|�k5[��~f��M�{���S0����\��D+3s9M�y�m����o�D+k��$��z*�Q���A�>T�9�Zi���[$m��;9�1[4����U
إ�;'�R;��<W���ذg�1k�7��CC�Z��>r��z������l2{h�7���n��
�Y�F�Z�Ai�o���/v�ۯ8H�u����Çx�;��N���9�4���۷o�ص`�S�l��v1׳}˶��Ϟ=���g���?ϣ
���7�H� ������=LgJ/�k�n�yhfgg�5�NŞ2	���ǡ���֭��,]ZZ��-pb�e�f��ܖ���YZY����Ȳ�V��4�+���g�1�BO2���u���쩉��z#��@,B 9���kߏ�o*A,W�������P��)b��"�C9�ŕ�tzߜ�Q�\X�q-���~DP�zi~f�nN(���J#O2A��=5�XM��s˅��N1�i��GO7��2>Fk�6�3S3;Q��[YYsK�v�W��٨dҋ���gP�E�Ў�dL�$�͉�ə�������P��K�	��n�˓��l����_<���u�P ����-��ѕiB�Fv3�~�Ƴ�\��?b_���֢=L'1�.T1���-<�r`�e �[�6Q˶lR}�����?z�ד$�rn.��7��/��[~�@�D1�7��Mo|��̢�0Q�l��j.�D��u22�� �ʢR2��~��tx/D'(HZ)�wB�/2t���E���&
�"��ǞD"��9�Q.H��|��$����߄e���f�
H"��a�t���,e�3���x�W*�_Ŝב��R�b5
�(B<��(�F|��$�±j�d~#�#�K֊�)a�n��h����D���i��m�.=3�@�Hkܰ�,V�6uR��]�0��Z�5�����<��uȴ��'�@��9�/.M�8�)`��rB�oQ.qim�-��%>27"ܤBhE��G��u��E>iH���SC�̠.� !su���g�v��t\���`D7J��>h������m�F߮,�����y���N�O3���>��� �q[7��e�ժ���:G��쵄W�$a.�o:K�v6�����w�ju��{�=8gL7�t̢J2�:Eh2���
X�R���� �8,���e�zH�O(�UD@H��K���w^��*�$��:`O��8{��u�\S�ٹsg�C�X��Hx���\d�d��Gza�H�4[�YXe�/�}��;tݥ-�5�z�v�-����ڲe˂�RLǑr-�8�](�p�tMɫ�+_�uD�E�`9�I������C�����rGm�V�t8W�$�&	HWV{�l�N�&��Z�.�=�4�i|VW��J=�1o۹s�a\�}'��^�V�a��z����/=z�hY[�n-�mC07 
��?����뿒�/�*]i	Rv&K}r-�
9�9j��X2�)Hkw;g��؈E[W9)Q �c#��w�}�Wҭu|��=��c2J<�!6�G,h\t eF�vF�d��:Z��M���֝-j�Ė4��rZ��},Ӓ��?�����	Ѳ�U|��ǁ=���^Pĉ�--����Qo`�>�<}�>��[w����.-����л��ٳ'T@)�2t�K�����^{-���/~�=x@�2�$����@�=Z�rk��c��:�6[���^ΐ K��=���l)�}�f:�� AAt���UH���ju���*-R�3��ݍ��q"ҝK���aЬ�[��Ξ�3��\#�zF����"IzJ�!i�\�-l�f�W� ��bo�e3����IoIG'��###�i�JZ�2�󦧧� ��������MLL���]q��g'���%�e=�|��@�o��c���u-}I$����=����=��q?2�F�=ݳ%ha��%7_IA��?^*��V �,�d��������Ǐ�D��8RF�c� `RveG4�D�Zj��K�!��-R�f��n���*�D���^��m&�?5UEڰA��Eq�(M��*&h�R'�k���P��,��5X�m���%X=B!B�	��RK�R7�K�����J��S.�]��_�X�z���i��Q�g���g���!��o�y����$H�BS���/R#J$����c״	0]AN�k9���,�<��s�0gw)�g�~ nQ�&g��"
R�|�1�W�hI+f�hi:ҙ4T��)䕸�)��;��c�SlX� 7:]C]��lM�Zy#̈́��F_'�W��Y�����V�gźt�1������Al^��h�:��]���1]���aa�q1��w�$]�"�߶���ِ9�S�"5�нo��3@	Q'_6�r4�y�X��[E=���E�zk�ze5�V�,�H���6�	���#�W��d�����LG;�
��4���U]_Z�,N�;Gw+���I���X]YB�N��FȜsTN@�5T��_[�o�2��ܓ�V�����n�5p���٘����ceky��8j�*Ć��^h�q��Ba���u�@�"K�E�m�Ih��+E5C��0�H�Ԥ��UfP����lxեŷ��߉r=��8R������P����:KJ��j��2U����F��T�h�������ZyQ��~�~���b�pUT��т�����ۨ�VW�	��q���ۡ���)O�5�R�$O�\-*S6(:��CUt�w5$L���j��4������ssK�c��k�ą>I}5��}���^��������!��������]�!���y��	�1b�Ν>y��J%[���.s-���i���6�LM�]):D�m�P�~-�Rﳩo#�5ܮ�jD	�x�9����פ��L YY[]�;uꔒ������Y�<�ؓ/N���eV8�3@ �%��*�jH��@z�)MZ
�,Jo��G,��k;���]b\��^�-��������s�&A��_.��Ґ5��`��b]R�U(�#{Q���`�M�>��E �������@����{����!^�E"�i-j��r R�$YBC	֙<us�w����}Y޲DU��JRj�c=y�/�F�ݼg��I�����s�~���=N��;?u�VzEA@���GhE_a�`��T-�b��R�>�[��Y#=�3��?;�c�_���и����>�{DZ{��Y��0�-���ޑ��q����}�]��0ے+�h�-�'��}*�X�mT�睪�J����JD#W�H38�M-ڔ��[6?|�X�Z1�n�
�4��5�e[��L���0^�N�0c�Qu�ܟ�<?5Eػ�b9C%	��{P����F3�rO��ʍZ Cd�Y��A���PȈ�6rU��i�����:vXǅ�T�ޙ��j^��ڱ�����'�����*Xvl�M�_\[�u'�)m|�x\��dN�b>�*�?1�X��"<p��gf�U���Lu�=�Û`|F5���3a�����&*
IƱ�Z��ާ���0�b
�|�hcܲ�P����we�T�E��� L�cydriy+MK?¤���"��;��a-f��oQ�2Fv\�r��j9�O����s�IUS�wI�.?�i;��'Af�?�i����詈�H��R�0j�+IQ9�[0�T��ӿZȨ6�1��H+I��e���HZ�DǊ)�,]z��hk�?o��H���K���c��ݰ���[�wƖ	��7����tBE������F)��	)�(��J�;"#5�D|ǴO�Q3�P2y�A"��#�y�I;�1����â��t>��j�(��:H�q���o�&�(,3Ljj'ITi��
[�2�2E�
�A�c�����Z]��ݎ��ʛ% p���S��y���[j�Ufe�s�g���8M�2H��"�c�c�������}##t���5����M�N����˴�����l��G$=i����Y*#	��
�޽{�G�H�4\���ǏE/O��8}{:7אdzt�Z�e��`5�*&�t5�؍���j.�ڻ�ܹs=�О={����?$)��}����<�s׮]&;Ngf�+�����Jj�̧"�"�b��G�ﱧ4�Щv���3�^�q��ZL%�l�@,e�*�����<�У+����um����̯�V�G�m ��בk@���v"��]!;���덀����	f�E(06��'��Q�jU���|�iiE�<��?<�>��ҜuKl����`t�q� �[kp���rUpi]�BfӦMa�pЙC7<o˖-�_=�Y$#B�J�"��R�QG%%�2D��ƨ�X4����Du���$��7������R��dd���OB�9Hr�!�N�O�<I��c��6��$��v�&M��s��[����/~��$��s��9�FAoC��L$m�d��._7`,�.9�6
ø�^i�J��W�_��=o�p��)��� ��DJW�j�P�ALA�^Y[[�r���/��N��g�{衇v��?�~�[�|�Yhy(B�C����;ż�d�cY�ĭ�n�)x�ˊ�턽��:oy���4}�-i~pB��4Ұ���0SA�	}Z_<x�S������R"�Y�.DR���͛�Ǯ��Z���?��[n]���zB�$�QC��>t���Ç+��Wk ��ܕ�;�u"�8�x+���){�}�z,��;0�pV��ߦw��e��/
9��Aw�iC����F?�ttt8�+�lY������d���H� �8��7�".�L�K�6�z���C
�>��:������������F���}����Sˌ'N�-p�NNL�=3Aw�o�Ų��%�#ƈ�;�U#Y^i������Uz4��O~�/��&�����C�&��72�X�޾>����&��9y�K��_M��i.#4Q&�E�"�X:K�{���cc�৑�i��]t�?��K���L��?��-qYA0�g<�*Xb*"I5C���`�ʄ#�\�1
‫+B��"�W'ek��j�1��"(�B�d�&��N��U�C�ʩ���9/Ht)�L���Q�U�~.Y\�HIϐӯ��'F]#H)T4�O��(EYv��aSB&x�/PĄ^�Pg$�P5*-�DL�$�����H��M9	��I�,l�$m#D����J�T� �Y�H�.W��IH���dƼo������ɖ�P˄�$8z�i۱O;���uz��)�*M�]-Y�,!d�"�S
b��Y�kkc$��7�7I6Ѻ��Ԭ�M�,6��E�1�h�.�,��!Ս��4��V��4Ah�(z��i��c�]d(X:��(k��R�PMꃼ�
&�2P���e��g�t�$�-_c��W�'�j �̀1\x�l�@��Dg��}t�ff	D�=eȄ��N}�I
2@�9Edr����I���jK�3����i;6O�L�)|�v4�S�6o�nO�"���i��zj�DP8j��N*@u���#��.��Ť����jpF�r��懨�ꖆzz��v��z���4�+u0F�F�e��:x�]�����+����0�t`` !��ػE*��u�+*9쾛�~��("���zRo���|q�M7כbzzzbr���N[�k[+����RB?S9O�25h��B&�S�b��,sZ������C�l�2V:y2�-�*?�۟��g����<R�Ho&m���z�t��<T6G�;-����TC�� ��PAh���UM�h�������ZSH��e�؊̴�� vr��"� ��%��uǾ��C���_q�5E'=�QtFFF�U��Zp��ǾK$i@�ȱ{��
�1�YiHr�WW���u�}����I�Y�W�_.�,#DmTx���m-q�y<��wb��6�+x��;���ۆ�R�I��&����ް����\,5�0i���YN>'y���L$*�gMS������S'�{�ȍ7�x��?^X��qo175]��[���n�Ʒ�M�\$�Ա�(lz�_t���tAF��J5��F�Zxt?5#��`ǀ���� �Rñh��2���AR3�EI�L�T������޵��G?�1�eg'��m�;��z�ؙA���62>>����篫����{��(!)���D��A�3��-L�s&���N�(�y��\�]m4u����/{����>)�Lc�AIH��R��R�d���f�*�GD��4=�Z]�A�j���z���#�\A`��w�w��C��^R��kbْn�l������� y���N�],c��{�68�SV�@g{Jp��XIwJ ��E���kj���(��/.Oш;C��w����|��@�u��ܲ�i�T��i���tnmի���猞�rsL$�=�L?������ۗϟ�
c#��&O�>n9�C�-p*�Jd*����2>14x��9zP�D���	.a��S�L���	D����"����2B�JE7�ypvv��l=���Uk�\��ys���5i�����6���`{�툆[S"%�0y�(?\�jJ��N��W� i���jV��$�'!I�0~`NE�:��A�F�u��V��\��@"p��/}���qz��-�~�.z͵啩3gO�=�ꃃ� ���[H�Ѻ�����"m;QhE(m�&ɾ��l%�nf[��N?rSϝ=�it������Ӹ@ގ���E��_]X�4�*Ύ�3��;�!�&6i'�+9k���zuye!�Ŝk�,��d>!�OIs	�� C�֫�*Z � ��Ĉ��%2�Ze_;,�}o��I��ʆ��B�J�'���O�z�_=���k_B����juLB�ӻ^�N��WF�?s����Hc�@5I�^!= !Y���mO����g\*Q�����CI7ԳQ����
���W|e�:���N�l�^*V�@ ��'�녀��Ĝ�!)�42�>� ����u�W��1s�^	T,��1�C�V���A�u7�'E����jf����Q6�$��D�b-ӭH����sr�QHP"��$�Gj�fQ�(�K"��vadmx�M��M;�q�)�ʖ�°ԘC>8.1i~�踠��r��h�Fຖ��4_$�@�d?������Ӑ-�(��,C-C&��� ��fd'i�?�]�ʐ�sˍ���q��ef�Kn�u��Q�1H|�^%?t�k��e@T�� ����D[dr�8u��y��t���}^3��E*)(4aR�d!k�pb]fX��9�M��m�u��������v�{)�C�Zi�����:e�Y�d]�V���d�t��>ƫ����η=꺶���۷'�>��aD�� =r����&J������n����ǎC� >%v�\e�v�jވ;v�q��~�Q�!Ow��\���i��Z�qP֫_��~spnn��Y.�K}��-[v��I����LNN*KM�E�w�!�@7�%b�kri�0�k�ɣqyN����V���}�"0�裏=z��s뭷"˶����Qz��� ݧ壚��'�C�@g.��a�tf#�E��,���%F��TW�)A�C��2�kɐN�K}.݆����%K��D/�{�n:ߚ<w���~�+�e,K�eJ�͵C�5��\w�֭���2�m���ˑekʞ={rJz����Ǡ���K21y�ڎec���\�Aʥ�PzP-����#����p�jνx�"A����w��4�tҶ����Z^2����굯}�o^YY"�^Y]�v]�/�<� *\����{\��v�g������c&3
��:|��㠖מ����׫�����޽{_�җ�w�}333��*y/��D�yzz���	���k,����n�Z�1r��h���$��d�)<�������.-���@w��2�S�N	�x�(���I�\Sy[�ǲ�+��4�gf���'O�<Ty���ؾ�_G�[_\|����9n��͵ZM��uH��K�����A/��w~Р�~�4�ؓ�j��W
�2�搶W(ȯ�v����s���@ˊs��eH��ܷo����/��T<�ZBo���ր�p��'�c�9]p���߲�*��ep��7�Idۖ���Rʹ7��/P:���hl
SZkt7�y�3������;���C��i|�m��6N�ЬT�A�;x� ���#G����~����[�ҝ��k��pj��qҾB}8<2B�I�>U��s��Z�133O���M+ ��Y�.��� F�AB��V0Q�Xe���޳ށ~��s���ڡ����^��ۍ�m�פɉ��kx�2"��u�]BC��Ӕ�&�=��-�_3�!�ʄ�1�f���b|�*�绶mE,�~[r�����R�2��j�DG���cg �n�IuH������Oԓ̞!��E��Z?�Cy�j�T5@���ݭD�&�S��G��!��{�!?�k�G�u<��F���x8���"�� ��%bӎ�yIӫ�f�*U��	B f#F�q�$��ε<�B�Ȧ6r7D�">�-�n%��D����s�B�:H�(@_� �N3�=W*�1�[�D��:V��rȥ�� G���ӗ<$	�<�T�n�+f)5�@U"Y&#]�ьز�8D�=��8	]D�&��,�
%ޢbX3H!�M��!��tMD�A���L���g(	��	J0�H�2��'$�#P�NTA#S}����ݍSKd�T��d��(��.mq7��~u�!s�᠋ڕ�Ӭ͓�\{\g*mG�q�d�¥�n4|�`N�Pu�T4�XE$4N)G<gW�I�4��,u5��1y�3�a��K��TΚP\�Z�i���x�zy�r��<����[���#;A��ΥB�]��7�����J�&r�j�����FFn��@Qfgg]��9���
T"�7��G�Z�@o�2'&&�z��Ĝ]�{�6F
/�*��u�a�Wi�:`Y9BGA�Ҏ��^˘�ׄ�^�4��)�s��%E����X_���\hL]� ����J�S(S{,G��փ��N>��ޞ�4�b��6h~'��ҳ(d� �.�Y�˲ᡡ������|�+����IWسmǦM�zJe�]e�"uc
I� 5�����(L����8�{b��Z���q�Z�e+����k����^0�CJ���y�2��)�Y�܏"��IIU�8F�v��S����R��������������G7�����Z��"l8I�u�II��PC��A]����?>�!���0�s�����M���o\<��{���+W�V��:�P�=Ң5�
�0uH����,�g^�i�D�ę��!��m�V�V�yz����H�"�|�h��߿�ﾓ��g����(�}�{�2��!M�`���ԗ�4���k���`�ș���.�L�	�)��p%��fx�4��y@˒�ũ*1 �_��44����($1kY��l��c����be�r�7���H�ܹk�㓧��Nj�{����o��	�h��pĒ)�ኼa�iI����8mC7]�z�[�k�B���!ݝ�"���(��+�K�fi+��Iy�����a�(���zu����f&
��BG6�&�
�F��W�D�8y3Igg��!ekoO3V���w�����C��}�T�:����n�����Y\�B͙�����ٵ����[��*�Y���)2����JUT�cwh��e(K��Z��53q��[(���ŉ	��QY���F_��5M=2����!���kh>?�0E�|xt�i��hrr�Q��J)�-C5Z�k� �ʈ3�����2��?w�Buf��P�Z�������a�¥��{������[mV��ޭWX�]<��/��!"��7ۮ��ܖ��]X�&z�ˮ���m�/ս�~�����կ�[�Re���}�ϝ�榫����Rړ�_�җ�Ϟ�t�yw���W��Z����羀xW!ƶo߲��?���5|��5W�t㭄�f�P���l,I*MS5-$�r�8�=T1�����H�g!�(G������R�835y�ĉ����/�>-�W�}5ͨ����z��0����}���Dhs˖��ϟo4���Qz-�^�q0g�	KW]�e�jU�$�����[�M��۟������Z�ך�YI+�={�7\�R�P��������B���@o�ǂP�'0�&��[Jc�~?��~�����t<QgI}6l�����m���ׄ�z�6,:Fm!ď1$��ZY��0/�e!����z&=�M�|�K<WF~�����/W�2i�~� ���%S�X�AO�'$�E[kg�[T�c��I�T݁���IN5.B�[|I�T�bҏ�X��q���|�I"�.(�m������4K��jcE��z���,�v=Q�R�	�(Į!lQ%�>Fq'a]�
G$3��C�<�43"
K�I[�A�+Lt@%iF���ȧ��fS�N�<��|�t&�'��Cj )�m�	��E$�#�0#F>I��冼�ʥ��ȼ��+�.�e���'GM�Vfy=�I���=�9W��c�=�PP܉k�B��ؐ�o&ͣ|>����c�d�&R�~v�D�f��&8%��V�qsqB�|(S#�~5d�`����r="��P'y;��"���3��~]m�	����C��X��-e��{v�	0�L��)�v�v�9Z���IdӾ�������+��z�����C��Z7���\.w���$ُ]��}ZO�ܵ5Ժi4[@�p]sמ��cG�=p� � G�[�j��&e&@����eڧ�zN�:e5}�x�m=��#3��33s�����w~����k����S��?���{�ػwg�	�=5�4��RY�&"�5J������H]����]w�u7�p���Jم-ܱ�ߕ/d�n�^/���'�C�'ox�]�h��"�����nt��� 9ʂ�c�
&�1$٣���!�.fM��1=������3g����n��w�Nj�>:T���Y���YX��tϐ��3�~L�2���g"�X3*��%,��w_upǎ��=��cHg*��:��!�(FʗmWOi#�r��?S�`w2w��d��*�/����8A��j���7��U�$-�i�ww��k��2���LX*�я~����)D����c�v�5}I|�b_���u�4��=op�_�F�-� 挅�$�D�	s|��4 $��d�Tm�B+�w߽<=}��?N�����q��h擄��?�����K��(F>�e�5�&�q2�lpppme^i� t�mzZ��-[6�������2�2H���gз�8xp�K�
˫���\{���|Y�Tٲed�2Ο���>M�~^l���]�������o��?8;-0_"�;* ������հ� T�t�I4e���Ltye�}.�"a��$C���������/\�0?3C������[0ODYK�8u=ziy�.���K��":��!���衄�?�� ��6��م]C#���." ��J��Ço
�Ҷ��W�I+���x��;���.�9Gm�\F�&A5�3���ݻ�W����Z'�7���D�Z ��U?s/]������sI��ȑ#���_�»ﾛd掝8Hқ֚-p������}���p��{�w��-M0��},�r�`b:o��Z���D[�����%�U�R���z��4��Ν����9���t���L�ݹ�Hc��@�A�H&5����j��|�#$�h��S���*T�\�+|f��#���\�l4����7�K3��}�CO�6>D};q���������]w�v��y��0��F�#������z���ڍ7����o ��8}������%�G�Ў��k�����<�
�Z/��2�.��9Ӿ�Ce��8	��k�h#L��{��<$.������{^�\]���k��-)Ӛ^
����z�S��H�S����i��0���
}Us�x�,qm�8���rm7��U~�	c|���(tu�CrQ����%D�mu��3���)��$A�T�OL�u�L:��++��r���Z�$�e�|�2u	vѥ~� �#P�����Y��p\IEP�5?��H7"%R�i��k�f�Q�D�G�0BtS*� V��2��j�Xt�D�b��PB5�4�OO<ڿ���2E��MDT`�8�p�p�چ�p��<י'M�$O�}~_hMqD���F� 5R�t߃���p�E[��&X�4V����$uL=N@u�X�ӥ�R3&xl4Ć~�F�0&��/u���k�����������%*��qF�9a�p���3�F��l���f]���w�3��gyd���.�sg�`
(:�It�tV+��ip��������W���93�FJ!ά-��HݶbMY}]���_fd����83� �p֚���4ѫ���z�9���u];Wp�0^衽9����X�B�qm3gk�v�Z��GH�;~�dA]�YY ��R��8��n����eڶ�#��Z�n������T� %wR�T]C��/�U��Vj�U�֡Q<�6�F��H��߶m��ZY�S�Z�ZK}������׫H��V�a(�BJ,����J\)挔��1��0i?���q�3N	ɐ�Omb&�(#=���Pc��_]�z�w��C���J�}o�?~�t�>5w�ة��ʈ�_R�Fk %����;1�'��[Up!�Y��u�;��
�Q5ז�C߻og���r��w��rm�r��ڪ� [F�y�	�t�d�L/��]�A�\�-�^�t7Z,�p�yM�h�s(ܣ � 1�j�h��MX��Z�iZ[^���@��e�~�ę��Z}lll�֭�|~����w�=Џ��TS��4�H�ǰaA���	�t������,��.����[�t-6Z�0r���J�^^5�r�Ҩ�s�9�^]]���0}�P ����������̙S'i�ڱc������I5[۹c����4�fŵH�L�h�!A"RӛjZ�)a����V���ru�$�W�W��S�ں��6I'�DU倦h9�30�9Z3$ �@����;��A�*��c���S�u%��/o�A¤s����d����ܙj�ZQ`�h5C�)29s�A=���@���b���`�XZ��д1�1۰�+Q���ql*g�1�O�	��$Tu%�Q �D�3�c/�@���������|�]sD�PbyD��@�0_��r���l�-| �̒&ɥ��Uk����7�a�Q���5ׂ��|9�zG1�/���feu�k��)_2��!!���]7\����jDIs��ej�ɇNmp׎�K_���<�0�Dc����{�M�%H6�w�z��?>F�}�(��kՙzehx�C�-{�w����ٿ�J�v���No)ҕ@����}���������W��W�3����=����8a�_�h�J�7�s�%���� �:l �٩YT��H/�-8j���x��i��XA�k^�R�ɉi0�6�Ǿ�f���[_|{�3��̉S���i��.������4�V��rmu���o���;��GP�+�\y啳�&	�=����}ˍ�G?�p��9�<���E%=ct@��]���d�����e��#�ǖ��Oޗ)\P�͏���Ý7�%fo�zs���~��ñ�����>�k��)��~(�����=9K�G��4A��S]К༄yha;��r���NO�T���ۣ��Q�w��YJv��'�œ�$��pA�g$V���)�]�ϔK�0i����ʫ�#��m�}�� �M�Ad((���tԴ��a��8�m�����[s|b���П(�C��|/��%؁���@�D�������O2�+yZQFɨ%���6U�M��4"O���^3�R��qw٨�$%9�X1�0@��G�T�9X8�*Cy�A.G���0��>�Qo��9ኀL�*�3�C �_�����0p�CI��ò�	P\����[��V��n%��<��d<�C #-KVXn?B���肒��l����9'%5>�#Ww�ყ@�9���Qک��t�!��]K���8���3�#e��DDQl�	/?�%��a��k�yYҵ����[���f�ϗ�f��B�ۖ-[��"a-�	A{`���^���A��kyv�ȸ&�@x����B�%;�i�����W��+���>&����]��eR�4Eǜ}d�xii�Zm�J� +2YXXF��%���/Ӵ�x�ݎ����1:�l2Q++��S��H�������͛AsN6U��>�IWH�\�&����W&��hx'�c������z٨��J������4�s�K֓6��.2�;�d�t�:11/�tf��mԆ�3�G��&�+�7�mq^q�'� ����O���R�]�c�:�z���±c��r�,U�꜑$��k�Y�n��˺_}�)���Q�4y�C��=͐3KU�d�3D&���3Yo��K�eI2YPKNf���KȪ蒵߆%.�~E96��.?�~�]\�0�+�d���z������%���A�eV$!v�2%K����&�6y�>����,xA�h��J����X�J����>d��fr5I�[�wƞ��g�����/����^b=L��Z�$�1%hړޟ�
����
�p-j;����Lt^�\�����>� ��]�K_��~'��/mu��vIr�r?1I�~ŮS�Y�c�ɼSD�?��XU��t��ŝ,-�	�%I���eR�/^��5[ԇ333�i��L�/�,Y���nni	,���O!'c��ے�P�̰$56��t^���A�<���M�z����ђM:QI�r�aE���Z]����=��跄��۫�����	4��˙,��~Bߞ={�}\���]~�v�!�O:+W��0�
��ޜ�h�����5�����ݻE�)�s�]������ D0���2���4�[�p<��6u��/|��������9L]�bIY� :���(C�Z �u��i)��j�h1X�U�4�:��ΧN���n޿����ym���ȑ�<~��%j�X�L��^�DLc���]��*p��!7��� �3����&)yDWGRdV��&�\,~����CG��H�T4�e��W��q`w�lsi�0	�Ө8�|1J��G�K�F0u�Q2��Ht �)t'0�!�,V5׋BB&
��Ւ#�q�Äm98S�|���*�$S,S�Q2��
YY,�̃^�1ݜ�z���*�4O�
�
�"��jj��i&�S�r���"���
}W��4#�W�*bc�4L9	[��(q����rv���H�j�M��\/Y��"M-z�rZ��(1�@�S#�cPc��z�H`�e�B���9�����d��/�����%"�o�� *��� �7��{Pf��o��%	V^��B~�V�*I���@*�+�a?Ef�l��	UԚ+�\^��y0��B�z[	H��sj1Uc����Yb8�)t�Q�kyr��E�3K���ܹ�3]���#S1�:f{6�8�Fȥ�S�f%'r�/~�3w�q���~)).�f���-R�IFi�Y�W��4O�u�͵��q�{)٬����`܎A"�]7�_�i��QN;41�Wv=�fmzn���&��
g�������Y��^�Z�3���K0[�e��h�oh��@հ�����}E;�sn=�v�s��j��5I�S$[�����K��pav.��_�����I������6��8܈���l/��ճ�Bj��^�rj@!���?���N6���9y)��2o((����&�AX`�A����l�2�����Y���z�*�!��Ҙ�	���׽�3G>�75^KB�Qv�n��˯5��,/33�D�;M���:P��e-ևv�<6Z�u���h�"�K��TWTz�F�5����v���H�~WFV<��'�]��P6��һuɞ$a��7N�qz�u	���+e�z��)X[Y���{gN����u/�)�z�D�P�u�������-8?�\+�RQ��V�F+���G#���G��)�*�t�߀)����г���"�d����O�eYD������2�)j�I]����պ�j-�rCԓA�W~���O||׮]?�ʗ���c'��߼k�ɓ'�NS/ΗM�?WD4q��Jd�@OU�"l��0� �� dM7�����
��gp��ؕ�ڱ�s�8ND^��VΦu1{�8��w�|��9��tv M��p�*-5փM/UVD3.��Vfn���u��
�O���.�醝�w���kQwi���l�U����6��z��v̜;؃�k�[� c�V9�����؅QFF�؁e-��km�
f+-�D�i1�XMd�m�h��
��ƕ�A����x��,��D���!��LÁၝ������cX_�җ&O;q�I9�a8�V���==n��bF0���J���W,e��&z߇��h���f�Vq�}7ggZ��\r
[��NC�X.��IS�����uE�E|���ݻ�t�O��e���?(�^�4�r��Û\��1�bn�������pvb����96�}������,��,�,�,J!�wtX���Ӌ�Օ�����@������c^u�tL�C��~���;Rl���/`�����ѵ��<sl�۵-���mYڱ�O���N!F��-�\/zы�:t�����V���al�����2����Q���(c##�;�v��MT|��ue�*��hO�<n�u��յ��}�;�x^��+`ir�CCm��^�������[��~�ߌ�_{��;��ps��UN��RV�U��@���j����F�=��xE��J	�dLM��	^����'9�t	�� �4�ҷkCk�Y��������9)��ҳ�|-79�Y 6�@n̻�wK����%�ХQ�z,�ץ�����k�'������^��`~��Q&�O:t������?'1Ȼ��F�XH�o���|�^�ʗ����m����E'��|�������y����)��\�ַ�뮻�N���=p�5���Ʈ۶�j� �l�R=�Ν{���?��?����{��h��+b؆����bw�����uB�Й�.cN-�dˤ��E
�ؖ����������ݯa���V]y�u��]@����t��_��W��go�������C���w�M��UB�<�	F�������x˞O|��y�{���w��#Hg
a�v� 6<�J�8�2[�d��t��+͟2B�M��%�%�H[2<����j��do���L*�( �7(��/�����%K��TS��|߇���?so3�]��<���o{�;��_�s��W�	���{�����[w^w͡����I������_����,��*U������}�Ih&0�ǈZ��Z�S��syʓ�=�L�!�O|�:%n��4���F��PB'���R$������rӕ�r�,)��lsW1�3��2�4�����c�y�,k��!�����A0�m[jW1��l����!.��N�K���
2!P�:��+I?&X�l�O8jg�m۶9�u��ŕ��i�&ˀ
 �c�e�~522B���cg���eVX��B�:eLR�v�H)s?��g��ʚl(f�ӣs�#�Zl�)�T��S���&;g��Y=���}���}5ru-�K�dzg��%�491�~�np�8}��-4[(D�C�R?���J?^�'a�A�����<�l�8��'s�ud� ^�mrQ�7Zw��P�,T�m5k����t�-�3uU9�g�H�.՞�M��`Gc�Y&sq��O�M��mj7��xJ�!���\���e0HS�墮�.ԫ���x�,�g��4͖U;G�+��R��}���)$���5��Y��p�Z�tgI_Y�XD�6oe
W�2��K8LBi�¤R���u�[��Y&"Z2@ �iQ4C���"ݡ)��h��â������X�8Q����'����E�*�?H��h�vm9�p�*��p�1l��n���oy����#�N�E���N���S(#��+S��Q�KfB��
��E�Ę�ր��K\�����	Ƌ���ZH,,
$1�������N*E�48���{n^�R�z�����<J��y�����B���V�7�]R���Sg�4��f�W��d�Ы�_I����Q��[&&q��j�K���XF%H)
�F�:�>�&9�h�ށ!��#����@ؿIM��I!�\Wz�B/$�%+�K���g56V�s[�Uz)o5��6�<Q��. %6�D�k׮��q��� ����ǳ8:�zG&�{�������V�dV0�_�ô�D���O,�z��@����:3%�׾�޿��|���ǽ���c����"�SZ��7|pim�W�����4u�0�ρvyB�_����<�صW�D��8H�B�ZA�����a�vE�𛒹��g�����oxͯ������Gy(�%�4	[`oVE�ekV>�����=��������k^�(���} ������~�$�+_��8�m��I�[i�@�A�K*Y�f��׿~y��i�T�T����-Z[�.`!��#OL������e���]�����{^��)_�V��������/.����k*�7��g?�������ַ�հ�]: G��Je�)[��&6�^I��,[.��X�N٠��]��/o.�6yM�^l(�%��徥Ȥ|��G�f�@�#cX[�]���0�7���_�B�ۡd(����І��׽��o.>vqV+�%ɹߨ����O|�ѷ��뮹J�;�l���-��]%���O�
!*x�Ґz`hz����g�
����/�|���%�
�D�6h�� U��0�� �&����Ε�H�D��LK�i~A�q�r*����(��0%�$o;�FsnzF����ᑱ�~��:�u�Z�6"?�v�:�\�U��A�~X��+aa�6�J*HGA��t�w�,R�D;C,�b�P%�#�U7�0 �?�|	�׳���7�
8<��k�:ME�t��KAr&~hӸ��g��V"<��V�éI���:+�"�Q�6���_����W����Bd�)�f�2�Ν����yOβIW(Y��9M�y�"�v�pv!���)-Ԑ�� `N�0M`)�o��^�Y�n�m�OM�\[%�!zK8�\0R���'7?�T���͛7��ǩm�V}��ԏzJ��<�,��N�8�8s
��זkEX��4�	����A�W��4��MÇ�ZXɬ\��o~�m?�җ���|������tw���HX��F�1��ϱ�W��7�qb���n�;/�,�J�Q�V�D���j@?�%�3}w��ٿ��ioy�-ǎ�WWW{Z�_�R]_��ٌ�XB��;H-��]3
I��@�I�mhg���� �GJ.JӐ�h�� "rP��@b9�A��)Ǣ	�5��QV��`K�-�=#Y��61[��w�<���?�i��;w��8=drǎ�JC��[��	��ZB��V�B�M�,Ԑ�Z3�k8�:H�Z�Qo��-5jnn�ڨ��T$U^IP�Ba<��-�l~S�]mԓz%V�wG��R��{{�v휘�����oƩ��%e�zů5#Zx18�-�Ѡ�z���eZ��}�%Ҽ3CK4��m�b禑�F��"��9��2a����f��6g��-ۥ-�p\ݲ�J��k!��PI�Oi��F���g����u~;�Q�PrUW��͡rg����DK� � 	0�M4�@��`3�q"�ό����g6X� ��QH�� BY��V�:U����w�*5&��Zo���r�Tu�����v��U'�J�0bQ�+{#���|����ںfL��x��Հ+}�um(�mh�+vq0�$�-��=388X,���h7މi�킇Xwt3<G��ݺ�G�hѢ�zv��
P͌IӶ�����>�~KABI�r�o���_�8u�K��@{L�9�'��i�����������E���c|�!)�::'ut�s�����J$;���`!�U~4�k�.S�f͜�p��=��/�Y�r�e��ö�V8k���Հ�=�F��e�̢�a��^Ƙ�|���}�Q�H�C�h/\��������0杭#��ej� ˎ���s�����C1v�ڶ��>���^yE[�3�.lm�H�4~b��v��9қ�y��.	��L�� ze��ܺ��	����9|�m��
�"����&�fG,Yx�Yg�<��G�����.c_Sv����3�!Ҙ�A���?�ż>UuV{9�X��0O/;��~�r±��8��\Am)a�!�2h|�,�~?���M}�k±$�}葅S���CM��1�jq�&���y�=���`NT�!��5�`}�u�,�1�	c8��x�$j:\��G���?�X�'�i��읯�F�^d���M���	�~��A9vE�ـ�}��Ēڨ�:���#�ܳ	9��*"NZ�P�UrT>�h�ؐ6��Ddi�U�p��F��񴰃���CbhX���BȋSQ�(o�c���ִv�ڃ㭭$��y��<�i��q�Ę~�
��P����'��zP#�;��ԦM�M�-Pm�PY��������k��~����={TEv�v䬔D]��'/������q���9&����`ٌ�l�5��+�d�p��˗ױ/X `ܡ�����_��c�
�LD�A���\sM�����^w�u�(T���_p��O?��/}i��Ջ/noo��g�ق��4nԍ�B���GA��2��������)��Zt4�����1Epl��&�5��q��ƾ��ۏ	a�/U�Ě�]tF��a����"�<yW�����'/;.�����?2iI޽k��G=::zꩧ�Y�&AT�8N�w���~�����cD?
y�6�Ts�	�SҴ�o��3範=!*�'���=���}�W�L��
�t�������%�:�T5$��^��Zݲ�����?{13��u��i��\|	�j�vBm��
Ls�8�'	�b�ҚS��ͪ{ֹwF	T�x�<.)a���+�O��F0t�v�t2Ѝ�uEY;9�����R��@�'}L�'>0��r���8ř]��"���M���hy�%����2�$�5C�QȉHl�a@��R�<Cm����j����{�?QE̙���E�(���#Dp�*�Z<�v��iӧO�qrH6B3ϡ+Ĩ�"i�#�a-��@>�D[�7�L��<R�fϞ�-�c޼y/���݉N3�4���C_��k�+��} ��A=t�1�'��b�k�  ��e��\E��D�����ӎՅ@��8��kA������qI5��*M���5���p7�Z��s¦J/��9@aR_ ��9s �{8��FGBP���sePY��UAĥ>�j�8��4��)��������w�Z�B���r(����ؼ[�aH���g��[�Y��pM��l�"N���AS��������ǉ���aj�¢P|C'�c/�����c��L���'2$<��5�~�p����}vc@�����qh�����������݋u��
���<7�0o�Hv_� _)z�$¶9l1sh�+�'�� ��G��<�5I���F@Y���� TcSp��l�pb�;�݂���^��$��`����*0��G�܂u>s�̸�ř{w�� k�A������:b1��2���>3�ku�"�󈏧p�$�lj��7��+���&u�/�y�B�O�О]*��l�����i��nD��j3{�*Zc
	�R֑ 	I#ð���ź(�a$pW�yx�L%�\�%P|�Z�~`D%�ߐ=t����G�Y��j��gC����1�UpQ��
�q��������
�Muԇ��	nս�c�&�!��jŖ�d�ҕ�D[7@8�+D�=+1�P����.bdH��N�l�t0�<$~��u}���^�Fu�U/�b�`��V��b,Z�ޕ|���|Y��d���ደ���5"��q�
Ϊ�U��[���=̺��+�F���$Ww(��:H�Lά�V�5�Jq�K����*v��+� �[B�(�V�S.�B҇u=�+Z�@B=��L�)	.f�7gZ����7���W_x��Ϟ��廦n
�p`o��ϭ=��O'�q����&خ'�`G`�D���]G���Ͼ���K�.	����@�,;��� ��\�Q���f�,cw����77��S�XW܄��'��c��?�o���\�����8�t Ⱥ*}���n�՟ֿ���C�Y�4}��=����X���(�.�����+M��^���^Y��T#�>jњ�*���&�-%R5U۲���Es�7�j�\w��w]]]�6�:RnohXy����r�Kϼ|��Ow�(��ԅݻwO��/�t��S��;,�O����,=k��~��w�z�S�1OЍ�H���S����Z]u ����Q��_��RM#� �i[�����%C�<R�C5gX��x�%p�?�Z����%����W����uo����z���Ӷp�eۚꙪ�`����x��uo-]z�"~�v�"	fB��� aQ�H��׊J\tU~��>{�1�=����_�bE�� �K��,�߁\D�%P1:59;����{�F��f��yC��?�,S��N�[�@oo>_��ƛâ����I��r%p=�r��\Sg[f��F%���C���d:>C
3�����ֶT*]r<�B�����$�ҙ\8��`pc���C;���b���t.�֌iB膜-�$M���F%ݖJw4����pT��QP<�ȏB���z#��:L����R����	�Sq�ac��s.�ע���jhQ��%ANcf|{��m��%�	1�H!�'���$"P!�����F�q�8k1�'N�0�Lx�b~�%i3T"���8�q�u}9�&�%(�N�=�K1�N�̺E���j�5يV�(K�=��"���1�4�x�J`5G����k�ݪ8���KQ��Vـo�}��"�F�Lp<�)4A�u���Pg�+Ws{Fu?"Lh��A|8a��/�Ǿ��S�lCb�L$�tI14E�WR���i��N�](���%kdd$	�8�u�	%ŉ4E����I�4�6�##�1���١����1v����#�7�i���Ut�ӨưV!@''% ���=����$���ha��ݕk5/��������ETq+�ԛ˅�kl*;����I�Q�Ǝ�<.�N�8�P�zl_�dM�F�F�E����F��'RB7��v	|A��Ј0a��bmh0(׵�������v�j~�d�y��l>H�0�; ��J�$j�&�y�������_���WF����G�31�3�J�'�vݕc��K\U�4�r��Q�5:��74q��x:�ѣ�~��Xؼy�_)��͒#�;I�C�r1%�.	V1yf̌{�H����{'pL��[��ӳs����mmSMz����Wu$CN8���7�'��ۓFj��`!s#�R�gvc�ĉ����Y�N���=�b���/����ι���1i2X�� ��1n��GFa�A�
�ʂ���^����T7���\���'���w�.�R��"E��~�.Pe};wW`s��_{j<�.S����k��克�%��?݋�{+VL����ݫ^{�թS�V,g۶m`��`ErB��	��S)?�RHd��O���SQuL7%�#"X�q�;��\�b��*�b5��q@J(���E�͏lظ��c���r�={[[[3�4�gXČb�]�6��֘������R��ZLC'��/{��L� n}w��k0����m�@/	���yr�#0��,<;(,^:.��K.�E����~;�,�GB ܞX��_;AE���ls�A	⊎Q1��*:q�h�04�݊F6���ރpOE�` !:ӥ>qdM9��:y1:�ٸ�
��i׋d�串�11�q�T�-���밊�<��pX}��*JQ��; ��S8����a�P�6���t!����V��kf|�`~�%��0L
B��C��%�@dO��D�
��q-�LD��Jl=�����j`�
�2��lI.���E@��� �g��lPEh�09as�Sj�%D@Z�iLa�&(��r���hD�~0����a/P����I��c��d����(���n�5R/x��}�s?���{�g���H�	KE"A_\�v-��׿���YF/r��t9<� _��~��dc���?N�â�;5��P� �ٯ�k��SO=U@�YE�Ї�V�X����o����/���� M���?���cժU����R�s֬YS�Tn�����A`;�L�UD.e�ڶ��׭[����`������n�
������P��x|��O����.����e�}�ݷ��#w>�%K�����p��~�� ! ���Gg�u֕W^�ʺ׎9z)|��G�ʻ=�����aw�0�[�b=6R�/,إb�zO��Ɏ�j1����}�u<��<����C߾�G��~:�X�w�(�}0��#e�O�|�ٳg��k�Lz�^{�W^	���?�9����s��Y�\3#c�j���<A~���.^�������8Z��*ڢp	�E����z�^�)�H�ɲ�
z��ߏl�x���V;�vww���8Ś��0!����ح�p���� �p����71�)�������+��ArQ~l�|���� ���f"�L�!��*�e���7����W�p���=�c�J�`�D��ň�R�����.@"�����֥��#�<P;�T<',�B�Jĩ�"o���ɱ�K��ь�8� �=���W�G��/�(�=�z���ل�����f
�� ��x�K� ��q�(5�9/��@�i��K��mnn���C.��J��t:]��1� E�3�?)`��������Wj'S���1#3�ҷ$0L
�:�g	�x���� ��yVy�Y#�����"�)��u':�r�kǿ��@���m]���Ev�jU�*��kq{��'��tV�>|�_KY�(�G�p��E��#K�;���#Z�M,.�T�q0DP*����E�`���1%�q�Hm�yM�����l�^��)�B�>�{����غ���y�`̓:���&����ZT����0�vTK���ٙjn���H75�?^&��_��X#�;w�t|��7��rІ��j��daʢ���p�s��|.�A�VH��O+�s,�5Z�..u33)x�Ef�x����_�
U�k	{��ˁ��^�arLYSi֜�܁�I�`T�B��ffd4��������P�zr��䇅�Q��X5]�8����ly�Y�E��l����&K� Ju�
T	��N�ó��ϲא0�kyID� �N	�,Z5Q%��2m`���n��ޔ�0i<�"F�^VW5Gu�Yb9����_�H=�[{��y�T����+��p��={�517���*����2Hg��ݮ����Z�q6Z�O�8l%�&�H�K�58qz���磏�I#��W���V�E�f�z��3�ZgQ�b����� ���u=�[�Ѡ���#����W:��r>}j�:3�4���5f]�3|/�.� 1NEa�*���yW�S	�.̘Z��Պ�,��J/FkepW Z���0�L��\��U���ki4VP�`#�^�:^l�A���7	I��z̶,#��$�f�f�3����>��.!�<H�Ų�:	"����l��_�14r�_U�`�V����-�禍&��f)s�uMߴ~�S#��ͧ�Itr���S��t�]��#L_�,]
���r �'Kتk�ܮ����W��5O>~�Ej��
p9�i� j��BIUL7�'�i��[��\���t2��z 7z�X��p�}g��O�Y��.�ͨ`�.y��%�:�׭}��o �i�I�w�<�ȓ�g͛9c��ٳ��8�Mr�������(+Nɪ��4h�����`� t�������6m�y�I˚[Ǜ�={���2/=����pCCC������?>8�k��Y�r��K�t��G����{v��EGa�:��!��B��j�(��FF���<
����|ذ�uAݸ����ά�����HW��u���s�]�mK���O;�4���LU����=���!�&fϙ����Xg/�'
�fͺ�替|�O>����9_����L���|A��[�D�R�.�d��!~�7��,]�pՋϏ�	��&l��o\��#N�oIȩ�w�R�M���qQ�,9��y���벪���zS:=*�N	B�HȘq%]��]�*��X��i��W6nLT�`�Y��`A!�����ݸ�s
��U)~șHxy0���!B+[ ���im5 ���d���� ��
"�IY̕�x\l��8eJs��]*����� �^�6�C$��{�u\8�T�#�x�hJ��<?f�-��+Y	6���u]�$ ����*g"�<4R�a7k�y�R��u�s(���]�`P��z�RL��h���z<z�d���9h��N01��%�'�WA{�6�=}J�0�gxt���`[�`��ԛ�#X����=b��(�tp�*n��� �C�T��s\�T5�l�{����ww777)������!766��:
[#Mõh/�����XB������A�V3d(�壢��x.�\c���Q�e�G*,�F�����((c\UWS�B6_%�hr�ȕ5��,�<�
f\�I��/�#�֎3�tA��n�P�� ��b��
$�WT��.���ٔ�كЉWP��ޕ~�<�T3v"�H<������������b$�?�rK����Ų�=GI�sʶDi�u�aqU|
߷�@W�:!p_2U�}C�!$װ�V���i���T�4�Z\J��d:pr�#��R�rYဋ`��
��Y-Q��02hh��Y�oaB���%F$�v��|�r9�v4��mFHQ�&/	�ȁ/��֥-����:g�:��c� �0a2�1����H�$ �Pӫ�!xE�vʦ�h��+���nVL�r*�oٶc�{%]�ݓ1��[.�%��\�Z#�qŌ5��7wUQ6�����S�ZMJ!��<锎��J��T2�G��B������s3�÷3��f����Q����H�MK(MM�����5!�I�Z2����
�LS�d����V<�{�c[�(J%�㒍�r�2�+Hy�(�P��/UF���Q��0Ml���e������@�(�wJHaV��m�0ĪCL�2d��(��c3]�bq�f���I�rt_P+v$)1Mƌn�p�O��d��B��6�N�2eʛ[�iZ9��^��wb`��뒬�F��"�����@Ҩ1i�k���F��x2��>�T�4���7J�`H�y�n�)�v��7�Y���:@�r&}J̣�L��j���(
��W�R��bM��m�]��,�L&ӌ�0�b��Ћ;4��	�R��@��*�%L��1�F:GͲ�gH�˕"�7 ���Gv�� �Frn"�_��:��q�0C�*�‛��Ph�r٢^Ƙ���!�*,g�\=�k�Q:h(�Ժ,�׻^$�3�h�!t��;0�U�5L�j8_	�ҏ�%�@`@k�Q�����N����o�����6�s:@&���%
��$Ҋ(�ݵ���֛��ߟ}�Y��#���y�57�����7��z�<�8�*6lX�|�i��v߽��瞫�v5<�I'/{��$; *�*"�˴i��v������]�j
���ٳ���1q�k׮M&���.���տ��"0���Oh�b��p�W]u�k��v�gX�M��z��������/-�'�3�?,�.x��������W�:q�R��d���Yv��)��iL�E����[`�.]�$�\)�z7��v]����?��A\���o�
H���o���+._�~�����)�������?w�����F ���8�l�<��+�sN<� %�t�5+hxg@�(ͺ�Q�?�4�}����������믿��+_}��+V`C�XlӺu�>���?�	��j�`�>��tvv.\��G�ַ�b�iz��.��B�'z%�H����qkL-�G]�#�b�
������^}�p�6��_�����W5���+��N���Ѩ�혂E�`?�L�}�,]��r t(���sυu��/y�3�T�1�H�iq�z�q#�Qk�ĩV��o��L��_�����%��p�Oꑮzz��e�� ��S�b$r_)Q��^##Xg%!�Y���}}}\?�yǎ�UZ�`��ɳfϞ=k�T�d� X;�R�!�N�0	[`'ͽ{�nݺu߾}`�aOdr�s���tL���(l����#�<������2����,`):ՙ�Ɓ�w-Z�Ā��W^�ᇪSl���}����&x����wͅOv���D�u�`�����̀h�Xp8Pn�a�'3f�iUI���C�z"U�*��P�aU�[Vu��Ύ�^�NP���XKƟ�r�p/����}�Vu�a@� ̲l�E8��]��ϥ:%���K����������f�W�L���p���\��N���̓���#�%�}��X?��@c�.Ԃ��z_p�̜���E�j���I\?�s�Ny{[kDu�� "}�ј��}�Zi��JI5��8i$��Ҋ���?�P��@�w�\��B��
��ku���Tx?<2�L�p*�L���@xx$�B�0M���Ar_nH�&O����[��ß�lm��c�6S��
$)Q'�:�>q�u���f�X\022���ڐȀ 4?���v������b�ϗ�d��䇩j�d�.��Oq϶m�8!��Ղ�B�b��H�3u�u;�9�s��w��S���԰���;���"�Vk��	&Z�+4@nM�n`*�A�Z��H0������fj�� Ft���aT&��0�%X(�)I~:.<��:HT!�����Ǻb�G�����x��/^�iDbw�^�^9#Y�L2�U�}�̶"VY1��QG��P���aKKK�{jc#o��r�A����)�Yj��r�+���@1S�0\xS5[�X�ðʣ�G�é�FB8�s�ˢe���z�k����`��}�K%�J�jx�X,�yR�i�&�ZWW(pfRxQe[1&�E�"-
̒�Q�<+�X5�
E<0˚�
������4�7cz��̪U��ٳg�@Oss�SB�x ��I��C�l��o�p��o���+����}/P���p��g�͛��w���+�O�����v6RP���^E6Xba~�Ϛ+���ϣ�}C78S�l���|f ��������W���1����2�{�4�q���/��O~rᅟ��J	�e��p�ݗ]vW��\y���z9@O���G�J����[�4o�LTO5�s`��-c�bC������;���2�������L=?�ZpH<�!{]�W\��i����>Wx����g�y���9�s��m��Y3c��I�F���~�i�:�{o����0�^�]A�����K�Z� ���_F�M����$bh�b��K:�Z����ӳdɒ2v�����۷�7D�3ٸ��_��ӂ���*� �vh�
j���������3V������>�3��4 QCҢ0��S.D��Tn�y���_���?��/��W�������F
&��*�='	+��b�*I��s�~�vL��{A�LT�Z���l��a�ƛ�|��3����%GT�0��oc9�_v�QM)uժ{N?�TAp%�w�# �'/[�c3a���v��ny�`���Lk����'H���.�TCq\��C��F� �����/~���������Ϝ녠�G��勛S�w�~Ιg��敼{�}4K-=�(�=�A5/?:�nl�kά���p6[l��:�~E�H-66'�Ά��Tk���^Q-:�Ňs�iꄘ���M8&����_���T�GX�u˦���I�x�I��㍫��/��²�HhXy���>��
�J�m<
5��o��5�_~�-����k���X �ٙ�Ԅ�C?��}�*�@�9�M��H���:�an��0�r�Z�鿟�ԅa��(T�:�j {���Q �Sm3�/�p:+����c�W� �pHHrLT� ~����_yF�X2#�9�n��`>y�Қ�ۻ�b���\�����k�42�=�۟�Z��� �z=B�C͕�D_�-�+#��q��Ƅ�7�2�'̞^�]{��%�n��;�53%e4F�����5#b�yK�1@��B���d���:�rs8�D[pL� �z�
���rLJ�&���)ݡ�?�eM4U����Fׇ�{��$uz�E62N�	%��@0D'45�����􅩓B��CGkd%p�$O�(�*�ty������[om��#��%!�#7M�n��e��h}U4�E	v� ��T�Uو�M�鎩S��@������ڐ0�˅t&�>�S� hѰ�����F5�	~&�:�:�>�)[���(4���0:d�M"qL�n�0�<�w�N��S��Y�4x�H�*^ G�0�E�t��]!�/�CC�R1��B׌�N��uN_A3B]A˧�����p���ѯ�,6�cC�AIDL�z`�(hWCVqV`���\i2��`Le(erqiN
�:t��ۍnJ���8,�ev��ŒF"�K�
��L:�g�Xo°@� ����ˤ*���+�"�rkmt��د���Yy%8� c��!��h*)��o�4�)����oʙL�H6W
,'��5!W-x0S�)Z�IGx�G�)�bz6��h��h��9i"���>/�L���mw˶�(ҩ�#��rP��
X<�İo,�
4OT �f�l���cO��Y��8��Ǭ]y�X԰�	I�s�q��I	Hht�!�:�75![fO��7�"�Y<����	,K��2��Y�X�� �`�y�`�
g�M�A��1TpO�����A3aE ։t"�%�-JC��(���U*X ��aa�\E�q�T��	�q3�ܨ&��ebZ�d�u
�����9�s��?@>��hat$��l�*V��BF�a�l+�ZN�?�L�X�qV��e�r��9���U%9ilϭ�#��'"7M@}�e�29�_�C��F.H �Uݴ]��`S&�X�6N��b�� Q��Zp��L���m��f\��u�pvЋ��]PoU;H�+n( ;�����(�����z�m��N�_�%�0{���T��O�+�h��+��r���)�(������LK����F�X��E?6�Kc�1�35���y4������s��t�>j�K/�Lr_߁t:�mF5����~.@�����;;;_yy�y�C-�K�"E�e0=�D8���o�v�W�Ʈ ZH#���=��̵��ލ7ހaU|�`���Q㓯|���������*;�����-��&������SO�\y��?L%3�G0�^U�z�S�jqW���Qe���-7�c3W��_YӍ����_��\�k��ԉ#i!�݊��yр��J�XB��������.AEս 0%�+_��]�����n;�G\�d2�?��ׯ��i��w�عs��K���w�	(h��� ��*3M����Y���;�W׭��GW|����ֳ�r�������U��L���^}u6����ݍ7�:G 6T�5��{�*Q�R۔���?�9�ċz$����б?�H}�O:�{�x짶I����ի�Ν��[�ְ䰱�G@�#��'`h���?��W\#g�xtNٚ�I���Gl/��u�V���NY�Y
��3:,����y�pq����Z��J�SN���'A_d:��ªU�fϞC����
^�) ͞'���K��Ƕ�����}ւ�9֚�b+�X��JJ�D����򕯜q��]mA���x� ��>��^zi�@���(Rx����E��	��tK���(�Ah����>������>�ӂ�X�p㬺�7�{�cr�
\_��C�,؝̱��F\�1����/�����]�2j$)�+�TLphE;AN����+�/\�袋`5�_�|2D�18�oPM#Li�@S�N�RɆ���yʃ��i粇�~&
��bTs�V�����y�)�+~���$����������Y����W����?��T��:����і�QXb>�ko�=88�ޖ���n���b*�/�1¨�]��OlG����6Q��gΜ�2�q�ҥ��2e�?t�~�=�`#I���w�>��=��3[e\hɑ��R=jᖊ���#�q\lƌ�����r'\�*_+.�'�SG��^�Łֶ�6���?0��Ha,b�7��T�{var�zD��{�Z<Q�BT��8���K2Q�+a9?\��}����:�^�"`�O>��gyh߾}vo/μ�>9?�B�+��E�"+��b���_����ܵk�z`���~f%�����ӽ[�z��g��=i�$r�ZJ$�~�+�qUE}
ȏ�J&�VA�u���j�`����K-��#ix�a�
�&�VPB`�0�M�6��៸����'O�8q���Ⱦ�^�uGGh��=p��ӧ�*c@�0`��-��@T@��:H����}�x���q�����������`6'N��Qc8k@Gs#0Kp}��(��'?���۽�l&8w�;J����1�܂M��;�̀�x�
0`S�����s�N��K�,��=vt�ܫ�`��� �n߾�4��t��el����sx��V�2�We��n���J�����1.rf����w� ���c(Κ5k���m۶%Z�`���"u�C�K>����d��ǌ	�'x�0@H����}�%À���4�>?���ႆ�%�q�zvw�}��4U�
u,�h��G����a�`��~�]m<�5�'/_��ug\�'y�*Q-�|�R�i1�A�FK�c�:�#^g��|
�C��L�&��{y�[��r˭���`8�a��t{�7F��E��Ѐ��cF�t*σ1�]$:�`<��
=�=`���0	˕ \T\�:��`/#+ �� �]�R ���A��6z�=ʛ���!V$w@k��W���\O$�7��IQJ����,�{l�X �1���ϰ�@��;c����-�#TM�+ 1�$��!��0�|�pBGH���	`?t���Ջ��p�4��&�2Z����ع�l���b1uo��*�ć9�n*��U �Q�'�,bY�K|E��/"]�$��%[)`+�|�2�Rg�y�e���@��y�c@�Aa��⋦^�	��t�%��u����w���n���?��}����Ψ�����bY�ں�~�*����?�u�@�"a�D������:��O�Ǌ��L�u�L<QM�Ø��ޜW׿|�m��Ǒ��!�m�&N����{����p�i ��x�ڈ�'D�qW5�R!�
���;��NTVCD��d��8�W�R�� � ��+p�G�?�m<���K�f��Ǧ�j^���]��z�ua#�np뭷������##��A���y�z͍�v���ݻa�}�_X�f��1��9}��w�az�1��dBîսe��ӟ k��|<q�bD��+�t��r��]�x�7��uT&&|ڴiO>�d�PL$c�������R|"d4�z�\~_PY���O?s�CO��ʳ�j��ݷ^�8��+�lL�hX|U�	2�đ��"�dˊ@K.��~�7������__���d��D��a,�GA�&rR���\� ��R\A��P��K�zd��%3v�ٟFV�0�(B�C1.�qO�>���>�Ď瞙y��;���=�=���H�u7
���k����b��!��~�����A+��[񕊂��FQӱP����b�*�(�������_���߻�DR�� �J 6����²s�y�5��}b��nܸn���9_l�T0���C�<���������c�������¦�4��+�+�b����[�1>��Fc�V�[|.�j�*��2r1�௘+M%�7��5�ȁR&ΜVY�r��}p*��C��z�e�}���m	̝��9��=Dtq�TB�$�� �o|�?|ҿ��+��ҷW��XxZ d��E͵A���p��Fp?�/��?�s�$�Փ�Z/�W�>��a����`k�܄p������b�$Te�W��0�+�4�a�����Gf�(��V�PE޵����j�K,%�)|����\Q�F�Jp�e'_�D���Hɶ���р���MX��I)?02���֍�n?v�@���K�垃�VmO>�tC�����ؾs��0�����5f���2���G��W_}�ٗ�z�� j �*Jy�h�����e�� $ GQ�t�r*�����4'5��D=*��р����.R�1�����זJ7L�6��pk�T<xPSP�� �d=dt
�*E�a	�T�(��£�@M� +���nc������gI��a�z��n ����(n�D�k��jaN�S��q��V=4�oP>��HH�JL����+б,�@�|с��<�#�� ��;����G&6�2�+6���8}����7+i�.f�2�h"�?�V�B�bP� D���Y�h�MLQ/9eQ*b{�jo.)��-!y�E�|1wOf��"!�Q�̳:��/d�V$t�o9��������s4����̜}�i�VY�a��]�}�so����;v��1g�y��A���u���}��F~�{���)S��;����w7��_�;������S�v��J����9�DM$�����Z&���O����#�;��K�����ƙ]�u��}{�'L���3�M�6����5��O��پ�iYKN?-n����Ԕiӎ9��l�w7�:��+6����?ϙ:}s_�_��?�DE3���F�+�N8���?hc��G�Zan`83e֜9s��J��첥GM�6,�7{�'�7�أ�͛�{o��9G� ��]S&w���e����)�;�=�͑�]'��ڸt��w�+��YsSI���͂j���dF�^���f���g'F����K'���ZEے���c�����K�qyV*�(�;���):�O>��a�.:���=2��:��z�bQ��/#�&�$O�+I,�P	����e�ۻ��c��a�ϋ�M���M�~	��\���&�m��o�5�
Q��1������{p�Lc읬kr��RCc�UD��!����ɘ%�E�;!��Y�(��`f�;�t�E��I}S� e��,�QdI�C�f$*ر��Zj�e��V�)��m$�!�omP���D{T�,Kqݐ��=ۧ�=�/b�11͢A�z��h-��zx��S��Ed��u,K��`%���ˮXn���Tc��]W;:&&��W֭��u$A3L��	:3_*
�2�b�37o��@$�F<�!?���CN6,_-�*v�9o��Ra�q�Vqr��-ۀ���h2�.����$-���l�\,
.���biɨ �� ��eK\����G�t������.l�ઑ�5[�'�av1 �*[�\_UO��/|�iC��K_��e���~��w>�l)fAU��&w���;��y�-�m9jA���,����NL6�
 ����t۶m�?��RS1E����b�E%­,[t�KϿ�է7��J�G
r�B7��{_�ʗ_t��]r�1}i#�]k��WO<�T-�/=�o��Y�T85bfl�G�,�'^y�lW.��n\�̒%K���g}�<QQA�ꊇhT1"P��~Ql�}�Ҙ6�<C��ÄR��;���
�A��_�7h�����!V��`����cz�'cD3XU�}0`/{���l� �P�
v�<s~�J�H�����]�(o�vw�O�~h^���͝7}����Fvf�5������/9�I���U�BY�*�NXt܉ϼ�ryh�hjҴ�TO�����V���\�/��� #����[�o�@�,���(` T_�x��=	He6���	Ē�[��p�����>g(;3jyX'�xb&c�)���^��T�+_�J�S�sO�*XPpC:�eJ�.\x�9���G?�<��My���Fo"8V�]G\XͧGҍ�uA���uO9�����;R�S��j�w\&�����O?�G}T��+���tvK�����
@�ש<Q���UX*նk����j�\6�iK�����O��?�s�g>�*�=�N���'������^x��a���W]u
�&1o)l�|�!�C�<c�<?�ǐ�F�����$�Q�$���uw~�"��+О�� �yd�/=�&��!��^j��,ˏ�
�;�%��O<��ܹs��55ݳ0���2���wQ��F��@�zX�c�>��'���h�wX��3�����,R�;r�{
�w�U�-<��@����Cs�5v����

�VH6�6�_|q��u��c�01Sh���r�\�W��E�%�'V��,�J2��E6�}�aS-�]�6��罦��F������ڴf�loR���5͘>}zy�*��H���o���K6�#��#�[�-�&S#�噼���7c$���������A�LS]|�aȥ>���$��F�}g��\+��Ì2�8���☉%�B8w�b�6m�4��a���Ř��<~�x�I'��d�t��/�u�K466
6"U��V�/�����O=88�c�mu���9���=����<���|��LTt���gCT�tbvJ�w��)`�J:��t�W\kC�-p��1y�"��5�?��8
��#�&���_a�aݙ�`| ~޼y�L@�8ΞXk�-�|�gҜ9ң�r�����gO7X<F{;�БG	�i�������-TL�`��ݻw�)��1��\!݊5� �3gΜ=>,�.�t�R��G/�gZWב>��3��v��3��B�4cƌy��"3�V�<y2fv���� �	*��'�1��۰fc����Z��0!K�-��z
�x�����;v�:u�1�l���p��/+P�I���O8���~�W@1~��ӟ{�}}�0��S'����n�t�Ygy�
7����G�1��l�Q���˕���������f�d`h�����=b��hi&\'gY\s{�]w���G���O#�F~7�/�w�C���'|O�S,^*�����`9���X����N�s�U�k0��e!���a�D2�-� =f2=��MT[�ы�9|8;��#�@̖�a�������z���.�l?a<��b16��NՂ�jYlu���ӏ�ݨ?)z~�j'�:�Gū�^r��y�*k�X�i��)+7B�U���
��vw�K�h�ۧX�={vC"Ϯ	���Xq�2��EF�[�`"Js�����⣈�Rw��|�bɗ�a{�e�*;��H�;B���>l�a��̓;�@����7�|�X����V=���U����皏r��!�*��L�x�q�/JN��������ޏ~�-���f�!v$3���o������"Ej�}�;Hu�b�.z����i��L��l���?���뮛5k�8�U�:�
bX���~v�����������г�����ww?��Oo��RTq-�u`�-X0����5RiS�q���'}����|Sk�򂤡�l�T[%�O�����_!��ik�l��������*����z�H,�6 � �L">M� �+!�Vx&(��ڋ�s��nUv�ы��p��)r��W�R�3�8��E����/��,�a����5����s�9�<�������P�����;�-[F�*$Z��V�+f{��p#�cnڴi�ʕ�Ev_��xq���m=/E�rͪǳ�M�<�˯���[����;V�rbc*����at�M��ov��u�/*V��/��������/��N��.�_��\�O��_7�����Wvl�0~+H ���B�޵/�<�/���]����J)�V&M���+o����w�u�+�iUĎxa��t��Ȉ�ܻ��9[��O5$A"s�"pw��3̪��.��[���ͷ���W�<�� �2�d�Z2t��(f͜u�E�Z������=|��'577IHV���t͐L��Ǔ����ӧI���*�������)v��ݎu��ݢ�I���?6��o\�)�i�Q�t���v�H�J�d뀃���}�����7�0g����;�<�.�j�8^��H���9��꺬
H��5�h��_�`ԟ��?k��n8)t<�ʬPq�p�8H_���ۮs��b(
�R@��Z�H����L��)��1�X-�9���EĞ-웎���EA�����K��p�Lj�������yϡJ�/�*=����G�G8�G�_!g>�ଂ+'b������#u��^�݃�eP*�`%`۷0�2���}�l�B��#M��v��j'�0tP��3�/Ga���a��0�b�4�����2����+jJ�T �yJ%�����
A�\-AD����H�L��j��ћ�|V���FB͹S�>��`�}���gTSi��`���l�t�����;�hlHL�ݑ���֭���\�� JDX�O�b	;�V膘��✓�g�fK�o�g�*����ך3X/�D���$p<�WhH�Hhy��u�;��R,݌�ݲ��` �ib�;l/��*�E�%=".c��ۈ.(	���]|K�t;�(��7��v��)�I9].�F^UJ��S�0BX~0�˲6h{V<S�^�9��y7��ڨ$��F9�G��PJq͋�>�\�)V��¼.�����Ak*rr��4�.�.g�quX�{�#Ÿ4��	;�F%�K���a`���hv��@�qJ0	�S	�PSmE��S;���s�J���V��[*4Z�����A�K�Jꈠx�^4�BQWC-����Z2�~l�#��TV��0�.��IfQhH`*t�@��TJN&�7�Er�ϷGaH
�x����yvc&#��GNeX��r�3����6���d ��T,PO��x�*�b`��R�����2��8�e���BBB�C�.[��W���N���3f��yv����o߰q�	M�X^>p`�����֦�[����x�'�������2�s�R9��:V)ݐ�d�v��5L�h� ԥ��[�1}��l�P�TC��֒w��iy�m*�޳gB[;��~䏔
���D����!�-ɘ�H�U�+��7j)�.in����cV��r�𱱔�:R�D
ɑ�N� 4�.����3u�MK��%��[��X$(�pbI��zC����]"N	��HFv�Y�%�t�>E�"�S�D���r9 !U�`�3+�B��)�j�g�1�����׿��N=�c�=�}���
 ��܈��b�ؚ�5{6�_���ＳN׭�푧.$*��C+Ls}�g��:�=C0ڎ	��ɶ����%��ss2>��C�G}t��}0���"%�;�[�VD�GB$������Lw��CJ��!V�ŵ	[�lihH��l9(P2>�O�4C �{��W_z9�I��T*��z���KlX�O��ݻL#
|0O�u���,��[ޅG��Y��g�#M��I�Gӕw�lA�v	+���10Q�&tI���N� ѷw��H��u�����0�iL�:�����{��ۺ�����TT�zuR�:�3+�q�X���>�ՀE5�$|�:dR�]@})k�$`=�`���J���f`0R�%%�w����ּp�)����)�;Z����_����Ey���̞�8�y�g�N����3k.���o)�|����2��1B8�Ba��'�Lu���.:�<�*�7n|e�8����������$_�XV,��q��i��M���@����WK��űx_�H����*��;=��M� ��t�- $FGG�=�\���؀�@ς�P�j㛲��!�m䦌��@s���_�җn��EJ-��<��D�
������5kV�Pػw/�5`��1�+{z<� �;�p LE1��E�8o��f�g?�Y��@��f�62�V�X��17,S&����`9GW��
Ƶ��{�w��������s�? ���F����D��>���^��(��/$��PP��=����5k�L��)E�|� S�^wl�N�}3�%�w���R�im8l%���m�e�������j8����s�*Q�:`r�r&�܀�m�x���/<�S��?��_{�5Y@�3eʔ������{\� �nXo�A���^x�o�K�A�ڎ+����T�\����O�>��O�E����,�z��Z�9���p,��%6���o�4���R�<�"L%S�Ye����������03����s^>6�մ�i��{�9Y�₧���Tk���]��q-�����'�+�\.��,�>y��2K#���N�#)\���?e������lDEB�F�3��Q<T�P�]ٲ���5� F��_G��z�1.��䋴1o
���6m�dd��?�xӌM�4iӖ-�f�;v�G��b�����@�a��U�;�d�^=2 x�jdd����������m�Mx��7����罂[(�DlȾF�tH�2�h�cd��Q��<��d�uXRi#s@��|��\=z�p��5�M$��5����PU ���7w�6�q�`�
9�A*�}H-���`,�-.P����^n��c�O�_a� b�Q���y� N(ɾsoZ[[ND�R��͠<S	P%�N�'===�o�t�{�>|�?�w�׾}�ؿ�	�#��?w����3��{Ӎ5�/����:g�-`H0����p�o �����ܹ�������Ë�ٶm�OA$��{��
��� �E!*��c����ܲeK,������ 'LȲ�0�---X�W.����c�ϕH!u۫�o=�H�'V���sܴip��|�3�ׯ�汛��ŋa{'N��{|ߩ3в���AQXT"�-����6e*��Q�	�Ti$���o� �������C��*��:8��MA�Sixh�����Փ�1u"�5�<�0�̷���J��ڡV��C�@Tʹ�ڸ�C���)�N�3A��Qx8��ʧ*G̸��EFu�/�{D�T�,�[L�~�p6����/��g��u��]��.�*��eL̵k����[�0��(h$��D"PD��:Ւ�2����[@��_|�'�-T���eJ����wn߰a���(W����=��s����7uɲ%w[�{	6%c���7	�qor�� nx	���gHxI ��o6`ScSBlc�H���t$�~v_}���1��gK��C��B��Zs�2昣��X�%fw6��L�8�|9�����l��=&,������D�X��	���
��
����m����� DA��	��4��q����җn��&l(��j�(���4����"����O�,�J.�����b��뉖8^���J�����O(vǍ�I�����L��:>:�*dTA~����̩u�uBS�C]$�s��p��zQ�|dd�v��e�DZ�_�����ob
!� � �(UF��n)8}.���SS�V[���}�k��+��w�9���رC���y?�0�}���]|��z����ۿ��/`��;�<�cd i�Y.}��Rr]�I�۷oӛ�����|�N"��'L��Kx�D�b�;e9@��i����m������^(�/{鋱`PzI�	~G5�\1VD��>���8UMh����p��v0��ߺ�s����X7mǏb^������C���U���z��? ��(Q�|��nm߹�.:�6�w�!��B���V�k~��m���������^t�ʕN���k:��QPYqa<Z��8��UҘ_,��E���a����韧�z��.#*^HqJ��d�pЖJ�|ޅ���tƖ���?z�;q�\�m+��r�j�6�gC������v��w��e�!IS�KD����m��nrSI=J
�RVP�����`B�S���):f23���_�_%\eKv�ٽ+����ņ�\&׭(�#���kN!��^|���2���L\S����Tf'y������0�c��aO[������a���}��w�/T�(,P�Mj:�Cw뭯�ݓ]��pJ����~wh�<3��E���2kE�Y�Eo��|�����O�V��_�'C�9yT�d����+��l���f��T$Ԗ0HҼ�Ku#g��I�N�&X�6�B��B�1��F�����X5H�c��Y��Y*;���*U ܴiSi����v�a��m�CtZ�
��]~^(�~ٺ@�3`_h�IP�}�S&�4�+H��͡�P,4�l'�4��+V�^!�{��U�N�~n׮g�p���avO�1eu�@Z�^�$'F�꿪jIt�(Uʵf�_���+v�Z�rrr�{���OOT�0d;"��>=̓]���aSQ�J[���
���w��~�����}��o;�5w��=6����j��*1X,�7b�5��YQ���I-H��
�!�D�9���]��Z?��td�	��5��59/Mқ&+Mwh����>wS)%p��+��T(�P#�f]Q�/,N��Xl4�����^��X�NכMÝ��#������@94Ӛ�%���L��B/Ċ���k��O�v,�`��
�酥\��t�^��(�Re���8q��՛f�4So���B����t�f����I�J�F���iV+�0t�r�q�N5�;Vo���ax�U[QZ*�-�\g�o )��_�R�H7���i�{;�NS���a�F�R�F�RZ�k;�T�U�>iY-�lh�B��[X�j��t&Lʉ-��<P��Y��,7.�����t�ϥ�������l+�o�{�.T����ycߑ���A�6��6[��!4�bu�R.�9%%E.�M�L���u��Q�Xo�!r"��H�S�Z��{�֬���?������>��U�rק?eG�E�pؿ)�*�a���jR$���(���95�;pt�E/�t�u/�-ؔ�D±�
�!��sZb�\��,T�PU}`��ܳ{���[.Zo�0���Z��� x/���\Z\��k����3��F�եV�1_�����S�v�>�t�s��.�qA=�rge�G]�R:�FT���ؠj�Yە-��Ԩ �`���d	��y��D�4T��b��R-�c,��P@S@�T����Ic�-TMC���kQ-f?��y�u�k׮�/,��xÛ�x/Jk��ݻ!��/<xO�K?e %���BZ��&y�L�<1�{�����-,�����-��f͚�
�k����,M�T��ڱgjv�t�br)k��m��s��I�dd7��2 R
!�dȯ�ϻL>ɤ��|��ʋ�v�ڵn�:���SRF�a����[��f�Sji5���믿����-*��3��[o�]7l5q�):�f��3s����?�E'c��D��Q3(���?���6Z�Y
o�K1�Dh�fjz��}ַ��(se��c2�u�����7% ljh	e:� ͙V��}��J&�C�I�&{zr���k��K�ʥxƕô&��+��?�"%%�Q�9M&<	λßl1a���c�[�����ŵq����M=�����֛�О��l>���q�%Z�?J��3������o�vi��������qU:����&��������cSG�����{�~�e�\�z������&R[QL<ۈ��:Z�����w�񒗼��x'&�i�=�T�Rz}�_*זq�W�R�ḯT��W~������(v��"�ݤy��Д���o`�8>��� 28�7�w�ׯ�{���7�����q^�{�S$�ԍ7�x�w�>�s�#�� 
k��8=��q�tRd�*�eJ�4��믿�������^q͵�$�M���'qP��v��j�v�4Hʉck�p�SO=u��|έ�=������Y/a8=���$��я|��/~�䊉f���sALȇ&�;�\7x��ӈy�����A9�'�C��ｎ�S`G�<�ZS�g}BS��sz��vWyӨ�D�=*$J�	/#fZ��P����g��N��7��|��/օT�R������|���)�-�.I�bo�"��\�0f��Ї~�7���UUN9�k�wʺ�׷������wK}�~
��_s�.G�����3!��Դ�܀�C��s�$0�S�+*�ui�'y�R ���,g�I��D?��Tm��Y��k�O�v�0��mSfN6mH�T+�$��R��"M(�KD��%��fDA��L��H�.�*��{i-�	��6 g@zK�8kss��C#C`�R2!/��l|^Zp.G�m��[�~�� ���uh�[�n�O��֓��b�Vcrr��գ�
u�5Oy2)���
ӢJ;j'�y�D������i�&�r5\s�LP���(@���]����&}�#Rt�������/`��˥2���9ºI����
��F���u'X[�N�u�-��	Z��7�۷ﹽ{*�
u�T�W����l۶���~�K/�����/m޼�����@)]�b�'lq��g�V���%�\�
e�RU@M]�j��=:�6���3Z�� E|��*�gb�&&&��C6������匭Z�s�N<������$��v��	�����и$x���Q��>K%3~ !v�W�>P�3'nC�8�7�Lń���c�.2���m�o�1�"X6���~(�OI�2)6�ό>���y;;�M�S!2첌c��18�i`������w�໘�6�{�s3(���1HR"%�A�WK���`�s촴-m�ʡ/�pg��<�%��Yvx� �-X���M�Iơ677�i�%��w"���݆���rN�N�W�,���k�B��r���h���ݿ��*�&�c|�Ǉک;+]�]�G�XOȽ�YiǞHg���\���=[>O;�]Rݒmұŕ�TM�S� JRf��G*;��~!]<��c�%��||����%�W�_�r%�R�V�[P2�u�謔�y_���B�.>�g�3��r��x�޽��(�>���,Z�۷g?�uJщ(��觝�rB:�P�YX'p���ϧE�u"�RW��w����8��T���3�(�4O�dNy��Ӓ��~�Pc��'�� �ش����~!��صlɎ${d�(�����O̓!^)�J��J�9�8��R�)TS	Ԯ�͗*�j��p�P3D��2⠒�q@*�=�ӳ��,/�����1�09���ޟʥfـi~P��R�x=M�	���U�g��������x�������I����'�Z �q���w��ݷ���.�r��%Z,fℜ0p��"�����>_s�5�r��wߖ�OS}��ߟ0_-�����G�C����}�s��;��G�G�~�;%�#iݼ:��C{�L��e�Y,)5��#Q3/�t���?�����G@�M?RuKW50��o�r
��9PM+�dS1�N�x�{������pC�Gn��o|��P��]�LUMc���[x�8�o����o?�����w��ݔi�*��������M�	5°�ۤځ���b�7ur�y�������4U�b��a����Soְ�q�ؖ-�XC5F�o{�����~��u�*�B�m���'���vz���aLS��'�ƅ�Fmf��>����Q���n�k��<�<�53���|ߵ/����ޔƊI�l�$���7�L���V�J��B
YH�tl��t������HfK�
wڤpR�nw��c� �y@DٜH��c�v�j&��>�q�9�Dq`�ؓ���I$� r�#u�������?�s�*%�bi&�wX�׽��׼�f�.��o����o��>�_���P*�:W �(5	\G�)T�:C�R��/?�|-YY���lҎ+e�,C�Q�����xk�R�|�T��[8[.������f���G�aBx�B��d�Qm-z�Q��Nj2h~D��:�f��Z�I��9��'"/��3�C2Ʊ<f�q� KՖ�"tL�G��V�8�;��ť�K&嶂IZ	"�!�x��q�x�p"#%I�嘝:$:�&����V{`��!}&�Ԭ�&��´�C�l�����#[մ���5Z��ǺIƳ<�mO���bu��su�=�E��Fȗ�0GedE i����G�bY3��׈y	�KS�IW�f� ����R�.��5�!iM�k���
d�z}���SH J� �t�������"dȂ�n`U� ,��P_yt���@��U��vv�B��D��Wy�M��<+�-��s'ˮB��i�F�uhّ�6Bʍ^������y�44���g�kW\um;T��?2�BwL��f�iCC��O}~zi|xrdp�k&"T�VQMMCuZ�0g�5���Z#���v�P(��-�N!�W�^]]j�U1j�&N�j�������]O��]�.�� �m�446��(��+���\[޽?6L�T.�M��5�h�����g����̝��+�S,��/I���+V����������j�Um�������#�j���odR�
��7Ce`x��?��9�,T�b�S����֌�\m�y�v��ƏL/�-6��V��u�W��F��#�c�+�|\qr���/���C?2�CC����6�����o�X�fpr҅ƒ�mٲR��"Е�:T�'}�L����V�f}��c0Y�L[6��\}|h�`�53W��K�κpi���;>�����o�����VY�:8t�^[�6�Y��Ha;�4Vm�2������������^9���u+�"Hjnq1g}C#A��ȃ�BE��s�] ����A���}�G�'Wl<mS9�.�L�(���jC�3���R#�ɲ�D�iY���-���KP�Fa�^+O=p �[���m(���`݄ؾ�fx�c��P��a@F�*�dγb�qD ~5R�����,�B�Q$�3p-�Y�!k���bVH��`�T�)�(�����@�cq�����'��U���֫V�p�R2!���\�w.--�E0���g��4� V���]�-�vG�ʹn.'4��%%�H"��K$	��,.��l�'=�V�?:����a������o���lC�´bW���!���֧� �F	�}T�U ���jڤo��{�D��N1U��e�%���)��aQ���ڵk��կ6�Uw�$���_������H�T�޳g�ŗ\-&L(���^��������ȰǊ�0+����F���o�6�Ē��DI�~��G�x��m��TD��n[S��{����cOL�8C���zx�R1br&:a�F$�R�NC� [^W[©c�a ȘFX
%�*8L�<iY��L9	��'�z�][�ё6�S9��L�PEV:D�F�K\0V-�Z�!���̆IY0�i�3I]7����/�x��5��ۻG5�W��5�(�k��:�^}�kj_����%�կ~��>$I�k��0LM_16~٥������w��?|���/y���Q5�V�9:W)u��o�����������zիb69ᤍ�+Ք��� "�ޙ�)�?��P���ZV��'O�J��Y�l�R�ka��,�b��dCF�b��n6�y����$��dH'"Ѩz����ET�5�׭_�m�a��q��S�|����XL��14 ��N����ȼp��d�U�g@�̜k5[�����b`Д�dN�r�z\aeZ��mhG�< À��ƶ���v��Hv$'����J�ʛJ���=��x��x�4i��y�+�������7	�Q�j@�e������݀��avl�!���;�����NhJ�ڭ;.��\'��d2�4=�c�2zY*�v2�7z*�L#���se�P�����@jq�m6c��ǬH�%�>{�T��1���K-/�s��xh٠� ,�&���s�8��߳����l���;��>�|R�����\8�"����3�
T�����G�Q��0T�N�p��jH����b�dLJn��Lac;O�.J��5y-��L�v��s-[��Ȇ]��,��5��c�� ��b%)G�f)4u���P�5Q�oj2%�N�zO�qw��N�D/����Ev?K��ً+���`
�4�~9��"!04P:���yH�j�SD�WL>d!Ò%:*��)4.r�(���u-�rtl�Х%O���X"�ۑ�a�A��<����/ĳ��~*�~�p844g�ԥ'YlK�B:0�d����W ǵO�:f_IfoJ������)���̌�\�a�\�O=�d8r�q��L���sss�#��*���g�AI<F*����~ZV��m�#x
ZXX���Sh�<�|�B�0�W|8x�j���4ӱc�T�Z�#{��=Ɨ���~�{:�����Z-|��_���a�)|?>4�.��}��a�齍�����aܠ2�!i6��C�!^�?��W\�a�EX�����V�7������裏�y晠v<�}�vY/�z��ЦL�u]�F�ߓO>�Ed�@W��%ȃ}{楢���Y��~Oz�,�ө�D�1��{&s.%�m�.�{h�{�y��_>1>~dϞû�ė�L�ڜ�>H� T���E�y�ƍj��9�z�!�憆�f�Kxi�T!���yl�:�\�j��K^��A��\�
��{���#$R�Z���4\,W�g�}��՘���ai��%�:�4AxG�Y�jU4��{S"�)J'�*�N�jZ�np�;���ɡB|�93����W���J�G�J�\��lxm�%�Ic6�u.��ט�Dz�w�ak���8m���I���$#�j�����e
.I*3l)"��������1�_-[��X��#q\18�C���)���X��"���N[U*RQ�d��K%3�V���,y"�א�@�u�p�e*�ea��j*/��fx���A�|�_<������q����DCSmڌ�E�X���'���l�[q3�yu���x�+��+��ַθ�"���� �����퀰�����\��R(O*e���b�ؠy0�:0ly*U��>�E�@3����O蘋L�U:*VG�O9\z}S][�tEJEK��ʿ�J���p�������p�D&Wp�	Р��e�'�4Nx���N;m�Ν�>��������$��H�:� Ӷ�\W�����Ͽ�k������?�я��[^�� �2�_n�������G?��Ͼ�U��-�Z�c�F��)�XJ�;E�S��R���'C4�t��@bd����1�)�-VD���\��P�(��%-\%�=#mA�������j�1煙Fj��Q*աI�}࣫7o�����w��=x�ts���׺鐱J�t�o�Z�WB�C����@BY^Ǯ�;F̲� \��� BW�ΐ�GRe!�nt]hb1�F�n�8LJZrm�J;:�4CJT��E�-'�!Q�
���E����(�Sp[��W?v�'^��_��� �����˙f����N��	(�ɖ�dͭ[�/K���Ө��ދ@�l�X猻��*J��*c>�	�-(���۔IutC��FVKUS4���ִ	M[�UPiB�Y%8a�(�9��S����R7�gp��:;[�Z̮-�d�>��¦6��^�r(�/�IU؁�K,,vh��*�4#X%>�҈x�Ρ�ޛlcL��04J� J�:����YI����R�*d"��!��e���r�N=\]�a��y��G�5���D眻ep�������Tr�b?О&E��NU��A�9�X�a�#�9��򎋿Vr�����0TJg5F�!I�aN����=���H)gI��8o��ZL�F3�AG���6�3�}C�����4���y.��ӢY|Q "��6��F(�L�H��!�g��ڳ�-�<j#�HM�H�$-ͱs�\�� C,KjN�ȏ�V�B����YN A��OEN��,X����*ڬ؃C}�J�v�N%Y4���Z���Q3P�j�z��W]{��mlUm���^�z՚_��E���/��|�؎�U6�\�a��3�LY��5g���̍�{6�nX���s���[.:�_w<���FV����/���|��sΟ�xƙ�.�l��+��X�b�gA�p�y�����+6���yr��ի&����i�����|���Ͻ�3�:��7?��c�2Դ�ӷ�����Wl<��f��}������^��Б�<1:���._���+��̳/\�n���;��6m9shl������X�~�/�z׮]�=�ܹ�o�`��3���Y�r᪵ݶ��Y�^42�:U���-g_X�͗��F6l8��h�D���k�}1�|�x�[�=g?�Ñ�+����k>9[5��.�`�V��V���x�׿u_��6�F�dnX	=���X��өL��2r8� ��ڬ����z��T�Ei��0��Wԯ����e�*Zx�+_�ѽ��6�SDs��3�fBh.z��v����&,I��TL�����4�F���ɧ����Rɍ�z}�qxs%,�MY|�Q�pt'���$�8i�ʹC�삦:QĄ��צ~�Q��v��27l���)g��:EOx~<̂��ꇏXãi�i��e[!9(>����\���lcϞC`67�M����s�\A�F�� ���f�����
�zS�Ӷ�M���ʺe�:
�<4@�e�,ժ�r�jA���'��Ì}��8�m��S"֠�b/������2��b/�T��Z���H������%���ap�(�v�V�Izo�����!�66h�I��b�5L�e��6�0��B�"> L�V4ʙFG�:��Nj�Z��q���B� gSmK��6����F1N��,˒���a�Op�����:�9�2Ou�j�,�r��~�|�q��-7�tU��yG�	�
d�T��<LI�'<r�A��'A�b��C
�I�)/%��I�j��[n��?��|�ϯ��e�.��\�LE@��~�۽g�������o��oP�W5T�(� �Yj���fh�н�Qn��}�c��ڹu�Vi�>:;�����_}���.�JQ6�DP�4�ʫ@-t8PH�uU��Ry�w�
�S}X����X�l�;�����mD�@����Z)�A2��V�j&	D	PU�#���u5 `:�WS��5�dlA�9ɒ�+.�Х��k^��x�6n]xы�*�Xt��@�_{���+�NMM���I��~bٺ��T�zD��wK���5�R���M7��-GIE)�6� T��|����G?��σT���)����]�x��_��!����S�A�(#��Țu���'i��?�-���`!z�Qծ��5�O��/{������_}}C3$�	��E�k������y���������G�(��2��8�L+��bY'l�����iMQ׶�)2�-��R:�p�ł�)����Q��O���o�]
��@��(���|��]C]��r\������� �u����K�1'���o?n]Nݱ�i��ojOv	�$��R�Pd8/�D���t���g8G��x2�LUz��Oe/���:�X�K�?����O׍�L�ϊ�m9$XzhNR#Ң	�USf�A֙�C�~\&g�2[�a�5�6IWO!����[j���������ô��]8�]�<���]'n�uGFF|�I�g���$w�􂱱1	&-��U���{f�A�Cv4������А���DsYkK~�������ǝ�|~ժU3���&�+H��VS6�I�T�gR@�8~E�֬Y1]fs�[�c�_M������ԲЎ�㺲Z4��\�lܸ���i2�@R��͛���/�ȶm�����Gp�T��&&'!8�\��` x#ڧĪBa||b��c�/ŋ��'�x�^r�%(���JeӦMx���虚6���s��r�LX^Ga��سt�Yg�ݻ�R�FG׮]�.m�{tE�+m��T;	�l,�$869s�~����f���:�"�7u��3R/�S�|	�!�����Jr�A!�&��ٓc�[n�lr�BzV�)��TK.թ��ǯ��n���|1���)y�	�ȗJ��z�pH���:Vص"�m4ƿ�X>�\���,��/�,cm`�i�СCx5�����ǟ�j�.�����eP�J��ey��)�X��9
�b�y�Z����3YŘ��.W����)'ʶȱZ�x,.-�y�c��$1�h����Z/��/����� Ur*tSIक़(Y)Qa�Iz�R�D.��,�,+��`:�֑��N� ��E��̽)�f��6)��0� $}�q���B��Y�	���UR��,���|�����n�Ї>��
�u�[\����â���v*���:f'��1՗����L� W���
�*��/���+���%/y�W��865z��~���D�Y�w�M���-3�/�%W�3�?�FSا����_�e��H������k&�Rhi���NB�I����+�cf�=s���g�,wS����J�{)2��l��=�1V���>���$�ơ%S�ibe]8���.�T�Ė�+�(ĔI�-�L{�� �SEץ�I��a����������:�Ƞ2��@ȥ�[l��s�9���}�. �Ů�9l!rٛ��&�}�{�H�z뭄B�RP(*��N/�]�T�<��2d�H�K�X�
�Y�X�w��AV|JS!2���>�%��e�)��2�i��"���Ěʵ�d�/5(�XsL����3�8
U���2��.��+���^I�GWL�-� �8��.��&N�R�ϓ�O��*O�Ơ[�2���^�}�ͯ���0HMS�bױc0��f���gB>?q�Y��X.�)�)\�DR	��u%��̼a�<Z�(J�P:h����+�m����j��?z��5W�K��!t��t{�N��Gh�`%J�B��Xʔ��v�\������9�cL�N�F������@�[溵�\)�f�}d
Cl)��|(vz�ڗ��ZȚ5�C����^I�v}GҪ"L�b��s(���(,H�V�T�C/���U�Iil�|��|i��L�^ozZ޴ۂ~A'\���'�8ȟF)l:�&p.�����h�j��ڲ��<SN62N��$m�hoI��@��̑���J�x���	�4M�bc�Y��T��,�@S"�fjX�bڄ��~:#U�	R�*Q�� @3K��$���Fu\b���b�M����%��OOǕB9��0hn�-SP�!r��o�4[I�[]��jd����z+)U,* V���j���6	�V�I���یc_�^�4����v�4cr�����a-	jQ{!jO{��4�E��i-����E�L�f-��a)�]ª(��H�Z�4baa#B����Р\����4Hh�U�m'i��0v�WtP'��H���V�7�� �,zŖ�OՖ*b�ـ��=ҍ�j�r);P�zx�M����R��SF�L�B��H�H(7_��P�5�ԩ��{�ՂZ��6K�B#�<��v�3��.�\��Gqm��q8v��(qT)�!�����S��s*E�t�����Y��/P�H�`۰k�fmGJ����H9�8D��M)f�(!��
k���g+��Q���n�*�v�p�]�L� 	Cq��T�#?n�J)ƾ��O���P!vS�E����‘rN1��Zԗ�n�T���	�,�?K�)J��\���t�A���ah����$��ȣ��M�)J�5B2��h1�>J�*�9B�8hlޢ�T]�JL�1'7F,z�qz�5\I���F+r�v���t��4j�A�o��S&	k����`�7����֪�{�<ӠHW�2�\j�˶��P�ݲ���+��~L��,Q,c�)����' 3
�R$[ҙ@�T��K�A���XIZ�a[Q*]��6�`$���ji��C"�A5�I3&7T�ڠ* �꘥8�w���B{�-#�R�r�M��m�x���A�bs��۾`���]���	_�!B���"�M>��^���]C���t��l�������e�]�}�����f c��r�(�}�]�J�|f~D�ad2�iX��
�)��簾m/����P��al������+�~鷾����'�D��>�h��������,|lA�6�AU�˭��%"N
nN�69�n���.8��xٽ_������W��W]sͭ��L	�a�d��?u-�>�rDAW=�
���e0�H��d���ډl1���o���]���P�&z�Z[����Ȕ��д���1�M5J)��`Tr'A���[k���DD,���`r1�v<�������w݋��wsA�1!Z��182<4PF�7�^�����f�LuL��n�
�|+�f�z����o�ʯ\Y(H]l;�kG��Ӎ>85uT%e�*�bc���ك��J�Uズ���I�/�F^��3�����z�WRz�|O?(e�҈�_�>>�ş圞�`�k��1�4ԑ���ԡ��Ⱄ�Ǝ'��"�|�v����O���ka��_*�d�jo���,&k��S��?����\[����ARHX���S�O�&z��lO�bO
�o�Ļ��������jnϲ�F��v�%��D�e�܄&d�\�(�\��\'|Y�gÆ+'V<��;w�P;ٺ������lۓ���-��+?��w~��tֈ~U2��ʿK�*�B��25:�Ґφ$��N5S��h
!��:�R}.7M��F�A�Y�X�p~Bʌ������!q~q�J��b�FV��E���	LR$d��(��?5�&u�y�O(��������W�p����[�V?���ʵ��u�]���v�����?��
����g�z�)�Ps�~�������|������;����v���� a|��_߻w/޻z�J��������X�rdd�駟�ۿ��/a��~��/����}�k�ChmNMM�~�̓~��ܱc�W���+V|�S�:|������?n�)1݃��o?�!�Y\\ĝP�z�!��!=zt]�a���P&�ǌ}�_\�r%���`�O>�$z���5L������0�+���/|�G04R�W����]���;7mڄq�W�}�+X�=ޮ1��Ν;w��5}�ȑ#G������|�W�c�u8Gu�f9_�I	m2n�P�[��gU�r�ʅ2��
����T�jan�܃ymB�Ǽ�hb��nJ=�ƨ-����|��uQ\}+��7rf���f�1
)B������۷�HP�ձp��АLk���&ʤM�7�h>ʛқJQs���~[*�ħ3MtR�*3��Qv�<�b
�E;��+�
���!/]�~�ƍ)�niԈ��l޼�֊�����w�$:��g�}6�90u3p-�������c�@���g) �@��*	rhqev��ef�XD��u*V)�e����b�ڵ偾5k�,�AճGg�:�+���cT����[�+���$i�<�ٓ).]"�E�xBU�*d�_����N����.�T.1Q��ch��JG�Wd�vޥ����!!���c�Y�0��Ӟ�g��|�*u�m۶�el��/���)$��o����>	�,�D&�A�!����Ҩ�/:Nʐ�G��������$���~����n���i�"JR�Cٰ:�����H��9V�����?����ˤp�?|�����g�F������z����=��<"�saZQ�����+Ib�I�(� s�l��(/�s�h\��pMr>e��?����wvA23yy �C��[�S�0�&C3"l��7U��o�������[^�Y �:qJ��
*zf:z4 `%(甈E`��=v�y�CQ��J��-��r뭷EI�y1F�7�x��o��lF�_z饘t�d~�E%q����Y/��f�vH`��Ne�W�	��x{��"h�K�Е�8
9�@���kg�?�ݛest�*��-"�K$�7�A�����d��n�*��Xz0X�N�nMEd=[3Ef������e�d}����ۗ㯔�����8}���i�/�H� JUA�7��2���bT�RVLC���ĝQ�u3O����S���'Vd��Ϲ"������Zd��
�g��t���Z"�H�(�)}�2��o�5�L���Ȥ��ʨ�d���Ǣ�SB�y���4�i������}(���7�Ӈ�=by6%#a���&�F�r<��T��D6(�D��:u|O����/+L)[N����&�g���&=>�l�eò� o��̠^�� !�s�$;���I;U.�J�)���N[�qc�Q��[u%��#d1*SB64�/��u�P����c|V<�LM��ݩ�n�h�7���$�2�Q�3����R�I��Qady�:�F�OQi?%�4(�E{Y�=�҄
R@0�%jf�eRx�O�j��b�K
��T��À"�Truj:e/�~�8m(�8��Gɱ�1xE�P��4�k��PH�����q4i�{h�F�[�G1f�V8S��a�Sl�%f���Z�f���xzn��ܑj�%ē�����>83��s9����b= ���>�8w���W]:6;���1���ꍦ���T��:6ut�vs�zcvq���|+�<*�_\j������������RU*𧣳s��~&�����櫵�O���t�o��y���1���o��L����;X�?}d��0�j�.�9v��@D��n��ߵ{�^���+�:Z�mό�3�S�s>�.U�=�?2ĢWO,uϑCxp�^��ĩ�J� ���~Ʃ����$��r��������;V�c|�5��0�O�~N/I\��]�텬tf~znqvf��,-����G�<R]j�F~o[�Y  ��IDAT��=���e�^.���F��l�� �1�|�
���)=���C�+g��%z�"I��;�7!��4�.�Ìvd�F����9�3r=��%,V����jn�r���kNO㶒��ib�l}w7�������B��ʰƿ�Iup��-?�CK���Eٛ�b:8�4����p�ĎfP1�(qt�����p�4XB�{�=���n���hB�����[6�MN��9\9�dsanj*��2S\\(>�t�Ȝp����𚕡��{�3���fup�t��M��왰]k6FG�םs6Y4�yo�R��0��dg�l$$c\\����SN)5*W&D�@~��V,�9��?�o�`1~��=q4�fԊ�Gr���b�6Z�>H�;AB������O�0LO�`Ղ���`��;�|��rihfD�Ρ7��	!5�eb�MP]�t��>�n��7<�����@�v������@�"�&�P�9u���2�b��9h9.�OF�a� Ls�G�c.K69P>����[�p���Dd�*Y9��OS��K��'w<NX��<H�nx�/o��_����c�!�Z�S�oa)9[�ھ��Ǽ�Q����r���
�G%����s�������y�G>�#�h�^�X��9I#"W��Ys3��UƝJ���\�cT:�$��9�x��J��zi�����htN�%0����hݺ[J�*��c�q�m���<2$�5t.\@��L}-Z.!p�js�U��X�����U��#6Q��I�R�0G�A��p�v��p�E��a$r�&k~:�M9ܐ ���Z�j�^�K۲�u)d�l�aՀ�	�UWOh�Ku�ү��e�z�z���,�W|?�a���T����_Y��+F���T?�N(/�g����x6��:����鞫�Și�QBA�%��S���Z�/�u��s�ڛ��p�9��Ҿ��Sp)�I{��-�D�l��H�^�XG���J�7���d(]?X�YFEGg�Ϟj精|0n��.��D~�N��y��E.P�����=�\l��̧���S)���4�*R!�!�����ST	^�p��Oe'���ãx�� :� 9��(�9��\H�L�o �G>D�����#��Jxh^@.�Ȥ���Sj��Tm��B����-SƎW�B҂%��NH�
W+�P�h9����$'�O�.�H}k�\�+��p�����ࠓ*������뮠Q��	ԟ(�Q��O%���k�B��������|��2�Y�o������֭��p�زez�5ճ�:kvvv��ݘ��[����{��ʇC"t���j���=Y�*�σ00��N;-HO������~����c�ti�ƍ�J��'�Dp��>˴.��g��@V�^�o~���Kccc�	�(�����G��g����>�,�422�{���0Ҿ�><��'��eYtq����Շ~X���g��k�Y�7`�>��|>��s�{L�p 6���۷���R��9��� *��1'�xt���$8;��T���*�$aK�t��G�����^?g��I�!�*����e	/t��|�����C��.�6����C�� ;v__EZ��ۚj� v���x�ʵ�����c8�M�O9�PV#��6��4Kk��|��22���H�]��n�,��%�RN�O�y�V�~��_]O���^���x�g>���_m�s�=睹��~����� ?L�%�\�������h�ꫯm��A�.���������������X���������h����'r�X읖xQ�-WL��5�������i���_Iq�+FHܶmF�w�;RA�g�=��ș�J��m8:Kw8�-b�,g�1�����mR���`���9���c;�:�F������ԇ���E�˶nI_q�� �m[�W�����޿磌�Z59��?���D!�K�j'�w9^�%�92�BpA�&3� y�gqmU�_d��d0$�&�,9�b�hFU��2�$tB�2��TSX0�1v��V���R�t�\�I�0�#ıO�˚��IL�]�͟@��E*�@&a��Ō�0d�N�Yu�ި��Y&JFV�!���褈gZV�ٰ�$j�t��q��\��Ů�K��0{��ɭ�Ri�C���T4���4����O�����d�U�ʳ��10&8Bّ��	"!x䣁�R�<eX��s�Z�2��Cjd�/���:n��,�	��'�p�E�ec�uIK�B�t<U�>+U�����3aȼD*)ņ^�8����~qD�S]�qⓐ�Z\1��z�sx8kg�{٨�tIQF�z�׻Oe 	lH��tB�S����
G����	����̇&�/;�w�zF��5��J�v��[���ܕ���
��0Ď҉(	�(u�B^�I�o��c�h��_<���uh2B{�����ɩ7D7b-[�&�����<D���Z�\IN�ɳ�9�d���$&���$�7�a�2�#^~�b/?�3�+R���p�sF��^f��l1��ҹ�ά�Sz�ȱ�QNJ�Kh쑒$�����	V�x�bN#3��$�]"sqeڑ.s��hs!0��C/X�H��9*wgpiUjM�S.��w**z%�Y:K�
�]�BG��(D��;MUE���j0w������+�	�,�RN�$ª�n1@v=�Α����N.ܓ�%}t'���e1^"fy���̵����Vv�q�t!B�6cj��cZ]�좡'�xud�
zS1�UM���Ks����r��3�34�;a���f�r�TJ��r��e*n+4RT6ݠtfr)Ym�D&�1�g��"]-�yho�J��H�sa[ANsWk#�G}?/twd�m5�L�4�o� ��в��\��R�+��y�k;H�FWT�ב�r�[�b%e�[���D~�ZNi 5(��)�ll,Ҕ�����|qp��Cc^@A/F����'��>�$���	J�)Ay�P�	���J,����W��[2}�Xż�1�j�jix��-���:G�d�5�GG�/�GF���n�ʀ�
�FK�,�#iGnB��a__Yp �^��7
 k?�F0'm/  ;�����O>���e?H
�>�C%�Lwl|%����u<�h���������-�%����}:����ba`p�VL7�rA�l�~�����w�n��Fa49�(�L9�R�i<D��f���lj�AG:d��jŁH�;2�F,(�(Ms��8������i�݈D\t����1v� ��!�F��ՕJ���O"3礖��L�\j.��f�Մ����o7�Z_k��o�e\7���a�2�[�j�����qT�(A��MϏ�("�m��@�1��Z1�ֆ�6<2VZ�b����������@�1g��k�{��c{����Wsvd�5��Ss3K�ULK9̛G��CO�@�ç�+M�Ǉ���R�ޱ�����`_#����(��|�R�U9�?M	i���}A	R8�Y^�^��r��CO3��R�RIL���y�~����D���� �ݼ�� _<��@C�$]|)o��}]3-J3��'�R�Y�F�s�U�V��*L��?�WQ8X.h!��:�����F�$x��|�zљg%}���paxķt����5�o�K~��))�6%��	c\�LQ"�?va��؈�vY�('�0E@hv���W飃,!\A����b�oim\Q�ry ryqr��իԡ2�T���H��L�&g;a���`����Тt�-&O�N�g�(� 9I�O��eXf̎G/��T��-|B�8^.HÜ�ם���R�!XY�L
s0M��6��M��.$ui��9~*G��'�VD��c#K\%�SĲ�;��8Z��>lU���� ������I_EƓh�rtu��"�l%��92S7�f�Ƽ�a,K?SH g~3�n�+�f���~ z�4=5��mC�ʛ(�f�r��&@��B��m�-(T����a�j��	����0%�����vDu/rv_VO��6��<�C06�-�aaĪ��/�1=���+��r��	n
�c`���'��2��#�w*�jݖ��)��v]��O"˵#�8��_X-ֲ�(Lu���.�D��U�0�7!��{�	�>��b��}�\�7�.{�j����%~�I�L�Y�����j'ϧk"��.�.�{y�[���+{J�I�ˎ���ٽJfR���,�Hɐ٢���l��	N$˙�v1ǲ!tF��9#���o�����k]]KJ{R�0����)JqT�Dx���+W�v�m�j��e�xn�>���s�)[�bNC"���R�㮳�翻e���ls�y�d}�-�T����ԱDZ[ٌ%��g����g�uV��B�#�A�̇m���Z:�jn�1�[���R�n��=������0ŭ�9u!����FS�c������nU)���W�������Sš���h���8Hf
W�':�h�ng�����b��Ż���1Dn�h�J3\,���2#��
%��a�I�@��###��*+A��g?�F!d�����$=D�	˜�"���8��W��+R*��}T}�U���aBsC�"e(1�T(2���2��}�P��J;g;�Մ�m����L�������`ҵ0d����H�kL��_�����F�wQZ��8���''��/�a���h�V(�n�4F�x*	���)���s�Ek�FySҪ��Zǎ�x�hJ�dS9}��!�v���Q� �ZD@�}����o�606����ŏ�1���B�T0MY���L��kq` �T�P�2t`ݺuG�7;X����#=��������#G���G5y�,�k��7"5�L�$��U+�^�j�h�W�ܿyr�b�s}��֓�N����C]]�z��]��o|���O�q��glڷo��ͦM����c+�|�}���@`��2_X��;��z�/��n݊Σ}l"��҉'�ڡ��r��CP�ɵ�l.����1!�1�:�_$����ؕ�l[�jպ+gxB��Ֆ@۠d�ƈ��;w>�����<@m�3]2%LQ��7յ�K.�d�ڕ�~���(.<�B����/΃��;gffv<E�ᡡA�-�y^�]s�52+��s��+��U,/��4^,��Ó9�wm��Ξ�(�lV�I�W4?���C����9'��Tz���G#��_�B�x$�b�d��P
�u�j�[�|�B 9���*j���t�uN1/�<"9Fi����O%��u��QD�S�Dٷ�x4z�ҁ��M�0&ǋ�NH��(��W9]J����2�Oo����������׋�؍'$Z���nI�/��:�Z��b^p��<�n���&	�����"�ͰА	�]i�%�\i��h7�.E(���[Mۤ��%�I4;�D �AXb_s�
�a��1��"��B�R���k�ȱxqL�T��9��DTs�+�	M��_�e؝L�J�����;WǇ��|��2�r}�΄,�#�p\ޥ�������*��4�7��V����}�8p����3 -�F3���q=����?�-�x�2���M]n(KY!J�N�b.F`��BN���#���!b9��4{"C��<QΜ�t'Oj���C-�r��=Ԣ�d���V��E���岆^8�-������ҷ)�>U�bR�P����$	9aVĂ��:�;+Ƚ�Ȅ��Nu<F<�D��H__Ĺ� :ȃ�� ��=IPvj�����`ۑk[Q��Y��~�jA�(�2kI��J��wCYqR�\zx��F�kL��;&�(�=J�Ժ3C�tK\ʁC��m+��=���-ټ'Sǎ��^���9���-�bH��H2�Y���R��4���L8�ҩG�f%X�{�WN]�{E�\�)�ݤ7(�(/�qy��Z����Jȹ��O_�[*�j�T���G������ŷ��ذ>P�-�\����y��SFuA!����*}9�N��􅐴[�?Wkb��6EI)�.�M� ��ȋk����J���NӹƢ��o��1�ЪIX]"���GMgع�p�%�r�ڄ�B��c�o�/����Y=R�)=W����5=��P㌑eСո$%[$�7!�2n�HQ�I��JU<J�b���t�p�F���XV-��������F�
���p}7��`�m��`��ZJ'�DҶ�-ۍ3�r�|�k�6�� 9�"����i�g"�\�ѱ)�j���dN��i����������j4��7�x�M�ݞK	�(kn��5Kx,�&�c�c��6��i�V���a��U�vtF2h	n��G��/�ڴ%�sG�Vi���e�@;�i.6lg��ݐK��57O1��ܬEy����A��n��Nް�%6����J=� Ee�5�el��.�ਈ�REPD d/%����Kg�K>�jR�ha��Iؤ�`Au�b�GiѴ�X�;��J�!mBq9-����DWI�QY�omw����x�Y5�zb2��\�o���\���~��ÊU@,�*�A�&TJ�u-��n%"͗��+"�,]bp�Jmk�{��l��ۚ�[����70(.*�;`xc���!�����p�P�Oc+R��������A|T�*dV�l����
))�}U`�q�)*�ˀ�0��V��G�9Âv�ӭ���i6�/{onYY��y���g�Suj�
�@��P5�"�,p 5C��ƴ�mǎ��Mn҉z����H�� �q����
�<��3�{�k^������gW��	I-y����{���������ld��FF#�<I��`fh��ȑ#��E����~������b���Й뭦���63��$gg4��d�	�e]�4ޥ�%(����{�����P�d�
�U�5�|,sӐ�'K�	~�Ɋ����F�HU,%Utp�maQ��c�ʆ&,��x+��w�%�!r�J�G�ndPC�ʞ���K�����Be[I�VǱ�̽V�ea�bC^��+B��X�l�\�b�O���==�*<L�Ɛ:�HnDK[���#�^!ha=��"�"Ԋ.����cW8A|�k���R��(�*� 0����Pc;"(q���F
�`|�F0�"�i�T�,('�J�]�b�5\������]�n���;���Lf(K������uw��&CWB���z�eg齮�]��!�C惐rpt�A�FCF�O��X��M���N�ze1{U��/�������׿��x����������k��?�<g<�V�.�dZµ��,b;l�#P���M��U��D���*̓Du��n������8���/A�j+ۆw(#�	'���_Lo��طo���<����dȪ���|R��z�� \�3c�P��]̰�0R�K��{����Lߋ�b��Y.��kN�F��B��"���\ʨBb7�!���x�Qڿ��w3�m��H1 r"!��A'F�F��w�<f�mV*�����6v>3ƶ�����1�i�>p�=��`�F�AC'(�Pۦ��nT�[vl�H8j|�D7B�%�v���sA@�Ғ�7.��P�VE��wBz�sTZ�o�b-�l#��*�w~gD�M���Dt��m(��������<j�M���NJ�S��V3��Lא�V��8��Q��>t�L����Cu��
���c��ePJ�e��a��q�i��w	�Q�9�����ET���H&7>>�����ZN�0� �E�צyE�;,�ũ?] [z��"]s�dصkWÖG�@|Lm��x�+���>p�@�Z�Z.D\-�"���·e���N�6�ʺu��6��4Q�w�Wl��*T��<���B�jqq�>5�v&��"�.�r7�/q.��O�XD�'��O�0PPmf$,�aB1���В�;�B ���ʔK�)TPi�j����c�-LO��,-��k�:�Ê�2�h���âY���؆�	w���n, ��Nْ�f�H�i�/���o�Ѓm[�w��[$�?�����QcvC�a&�ԅ}}}4�ǎ;yj�OO��X��gηKvl�!�����ܹ����<� }�v\N�02r>�����t�_~���}){�YqStN�ĭ*?��9�U�'��L$���L���䎍=C��,{�y���aL |�@�i��5P�{�g�6}�q��%ޛ�0�eQ�`��(�>0t���-�mQl�}U&�8D5���r��V�-�P)��d|+�ucWDՅ����߹���b�`Y�$w�A�=��뺈r�v�KE(�D����t���ϸ��Sᯚ*q 8a:�0P��LQ�j4�!^F-�{�M@�لNn�"���d�8!��/U[�*H�ՠ��ki��<z
�P6 I���	N�4I�'�槩����f$�3�	'���_�t��u<���o�<�oA��E��S���iE�q�У�:Q2p7�程D����EN�:u�g}U�Y��غ���� eѢM����`�ڱRi%HPx�Ri�g����rpK��>G>J��l�k�p��2��I�
ا��rZm+������>�)���t�d��,���i_����s�s�M�6IaҮ5b9���CԱ�$W��g�覒S��Z�3��-F�0d��>L�B�D����XK�J��űV�ע��ѭ �aچV��f�V��ӆz��`NӚs3��&mc�N��3��X9.�a���׿�#�ݬV ��e5�����������t,���	�DK�x|�ڡ��c����&�4QY:4;�gMr
����?�f�Z�4�{�|5{�ؾٙ��Lx�2��lɛ���Z�{�t��h����Y�ʵZaƍ$���C�nH�4��ɧ��A3����_R7G(��F&M� ���(�#3���'�:��)^I�I��V�qD*��E'��p�3�`̢���{�:~���iN8I{H�a]�ܲ�_O۷ر;Z�hY�� @QM�A�B[!��=�i`�����|�����\{���HUV�n,"8�W�H��O�zE��Fsrv���fӉ�L�%rDP<�l�j��hr��gk�YY9~�x�E��ɚF�WІ����<ѿyS�h����K�w��]�|U�sY�hQ���\��Z�֒&�I��!�5#���6�)̈ }E�׬���;�̸�?:=�:Jd[�a�vN���v�E�q0��A��CESB9�t���@��frv,E�@��B�4C�X���#���c!�����`M /��ı�v�U�z՚��۹�kU���J��?��S_���F�N�������)%�7�ϩFsq%����w�M�~5���w:t����nت�Z9�We���s�&�ɚqCJ�Ǒ�x%�|�9���`�U�E�B.W�����Q�x�y���.�U]Z���{���̇�ɧq����	3���e/�Y�gٙL~j�dƄ�鄰��icy�K�S�p�\�4�?�v@+��񉙙� BA����>����)^u�UY[+������g�P{C�[��KA#��y}����4���Ff'����
A)u�u��D�e�/�x��@CD��3�C�-Z��*j���H�z���1G���GP�r3Y���m��P-�uKgUg���bT'�S�~�
� ��,7�cofA�+f	Ĵ�y�5U� ԡ��nH�rRIa@WU�Ţ��%{�a'ҙ۹(H�X'�&�H�SQ���2����u����䮮q� �PBt�Ƅg<I�x��4�w
��8	�$�D!@&�(ȘF�b�%rq�����	i�w�����6�)�]��`��ل~���o"u����=r�6"FP��b� �j���t)��&LK�k�Ü�T�)�!=A�i������� s��J��������{�/����ő<��(�Ij����pz��~�CN���ș����8��
r����ț����<*sS���-��˦�"Tt~��F�8�ҖF��$-Eb�HS�؈@{nj����B4f�_H����Ct6:-�jta;w����EKB9Dȹ)���I��LQ~!U�KM���D�0�I����h��Y���u��eU\���"�M2h�ݗ�FݴI*��9��Ap+GJ�����]t��5��yL�%���������b��N�>=��@^���^~��;׮������V�k��.�6� ��/��ر�44@'����j�tDe�@�D��~��c�=V��j��	�^z:G�L�e8;��r\J��k)մQ{��nݠp�D5�Ȗĝ���9��ts\"c&�0���]M:��˸wj�f�����x�H5|%�����n���O��;�rG}A���{�X�R�4����@���.��@�<љ�]�ܒ�aCx-d�ez�EC&�&��~��c��F��d�����l�]1[���-�VV�\u-4�m��D�r#���Z�P�\"�U �gc�Ab�H(��
��.�K��.�����pzi	�m�AK�6�ݭ4Zt;1�.��3:*�<�-�Bߠ�8�PU?-U���������iёe4�d3t�����֌�q)��S�8@��h���dh�֯_��k6�]~� @����s�_�������d��m�$�B��ѩDv�w��������N�<{y��\�ۊ�� y�4&�K��h��:y�$��)�}!�J#o�:��5c�x��dOM���O�������5��H��9>�v�Զ����1�\01�����Χ{�{��ƍ�p�����)��G��s�2����_����tׄ�L�����S$��G��'w���"����(l zD������a�0h��,X(��J`d �U�F�u}�C�	k��E���*i������z!!��:��u̨�11���l0"2�4�BhF�i��*r�Iz�H 0�F��_�1�K��;	+�[p����lb3b�͊;��Ң���~L}��CqU��)�%��;�T�����fƥ۷-�1��f�\��j�����gz:�lh)�FZb�A�0Q��(Ss'BIR�ǒ��n"8g�タ������b�f�K��>o��3�/8B�z����2���sX�>~�Ϲ�п�C�&��8�����hE��TD���/�ɷ�ʞ'��>�(�zw�,r\R�N6�q��H�-H�uBD�̌�/��Bkx�)�6o����~�Z�F�U�L�?��,x�m�J�ZZZB6�s.����R�,��� ����DƱУ&)v��{ʓl�zŋ_q��k�;B�N�CP.�Po,Wȣ<�p;�/IN�i[V�nt1�w������%2�]2K=y��ފ/�-��1"�<��@�z���T,{�oe��ظ��m;��⊂�'/�s������rWn�	z�"/r\S�I�Te��K/}�u/�%���4룙<�a�UH�*}�+��z|�F3�����Mj��/�-���WBBys�֭#CC[.��.�bhH�I��[;�P%�����믖GF|<Wa��9��y���i�:{TY�D&\7=�L�]�k��ۋ��䟝>�7�7:��̴��V[)��w%F4S_z��n��E�Q�yP�db[�;��i@�ӛ2�r�!�A�)svQ�`6�aE�'�tQ^��·�a�V'%�9�"Q�ع~��3e���Z�d��h֫C���]^]&ZJ���*I���:���3�3�ip�A~��� w�y�ʑ�S�s��4I� �����F������[�|������g}�B�a-D@��o|C}nqM��3l��'�9z��]���կ{�_�\C��74O�j��M�^(�VѴ2v�ݚ��#����A�uY����v&�Eᣇ�a��r������}��sӐ?6�l�=��}?��v`e�M/ؙ}���7ۈ#��i���|7h5��P�V��3}�����C_�\�8���u�j؆�I���4�9<ک/ʑf�qd�����:<:J֩�8?�0�$����Ņ��A�,,�m�ֵ�iOO�42Y�,1�o�s���с��-3KK�6U}�[���~�z�E�&ÕZ"�#�����J�0s,���1i�Zv.8����6uslt�\�z��V,����Yy�9��|7�VZw~�s/���&�%u�\65��c�#Gb�>?lK�G�q�� ��C��ǏL<x2c[kG�ˋ�"��|�:?9qj�py��X�� IxI��O@b�i~{y�(9�������ŝ[6��q�57[ֵ�.�Ԓ��S�Ⱥ)=!�	�短��9�ܳ����i��ʺ����E ��iP�R=/0��n�CR���*HС��F��8��kY 7,4Z6D�tA@� f$JPB��M��C�D�����(�xJZ+�ft�uۚ�*�3q��9dHrv>�t�"T�dh|B��� �7/H���tטt������c��\�|�D�L���pK��Y���i����}�H:��e[o���ʦ���d�~�A#�x2�IYd��-XJ{MShYGH��d��(������֡-[��"�	�����5�Y�	��)`gQi�7h�Z�AD��: ��Ph��g2��W��KC�/Z1�tV��G��8���玟�8+��W�4Z/�bpu���������]R�z�(��6	2p䝟��ڰaJz|�KW ������-��؎��m!���ߏ����]�Ve�O.|�z�W{f�Of�Y���� �k�Z��(8�L:W�����s��Iܮ#<�8�+���Q^��	wDԛ�]� 7�[~ӛ�TqQ������������1�m6�"�f���ozqvv�QgV-��&{����l�3L/-�hd���$����Ź��_t�������N�Mәk!*sQLWE!d����קGC�S��O?��l�!f�����.[��J�r��Az�H_?}{�G/~�Þ����i�޶nH�ٝ�DN�AR"��JG�3��t��.֊{���B;�~�v�ԥ��P�_1�q洀ԓ+SeMj!@�ɢ���Ժ-��D�R�^��dD�9�\V=��ŜC�%i5�f*���'���d���z�@��.�Ģ=+؂�Q�	}�h��ۭB��������~��N�J�ڷ�NAش�\@���-�ir�J4UDb֋b�K��������[}}}��ĩ��r���>��d�h	p��sv���B;+i�d챱1�~���E�>���K/�e͞8�q�+��-K��;wx�*�(W�Ыu����
�j�:M���!/O��l�����H�bJ�|�i��ށQ*�e�Y4��e�>�GV�X�Z8}zq�ֱ�'O�?t�\�r��*#a���~��_���h	�KFw���n�]��rmtt0�W:���m����u��\���*���k$�n]���B�K4lh�[:J�"ϡQE����h仸��~�T	i��ހ8*�4�־H´����.CwҶDg]�H"A!��l�k��IY�����8"��z�c����42�K{n�?��ā��>-���iT�q&��_��=�MDϕ�aP����n�@K��-x���@O�몦ES���W�ؘ0(�C�ƟN�$&�Hӡ<E�\� *o�A�>�A�Li�p�p�ƌ�d�|�g	0�	�K++�������h�RW�1�kRz�CwL�#&=	^Y]嫎��U1ӝ���v��� ��{���5�eM&`	#aQ��GIt���8�."��̘�$���Ǿ͚���L���"Q��>+�NIX��o��$n�
m��O�����vh�0�*3^�"I .�� ��%�g>�sX��q��)���82ؚ^Ā=L5҉�(���>����W}.�b�"d?�sV���u��.s;n��f�IJtzE�8?D`T�B�	 �˙��"�e˖B.O�@s�s�]��lĩ����:�L��������%��=
���G�#3�43m� �[�&p�h�+'�X3$�͒~��|��>6�hr��&��F`vy.�����B���sI��R�GQ�t=#��i�w*����i�!���ɥ��Py���d+!�.��v~����aCV*Q���Q��H���|��4���4�h�]/�u��vj-.���R	pf�K�B�ї���©	YU�"xJ#'���o�L����ԏ���ѩ��5<p60bg|K^�^��'����3]\��檝�W-3C �}��~{�BeK����O%���|1�����s�)�͗hb��4ms9���+�.+�,Bl���{��u�7"Fgot� 	s4�!�
;Q[�6��H3����.=
Gn�8�p�������/�
b]>�W>��K����'6�$�:��B�M\g��:�iS���TV{�E�9ad�t|,��]�x�U��)�$��q�Y�otX�T�.�C����sV6G����O=��_>����r� ?�N�.�^�:�U��E�2�^63ք��U_�ɖ�v�8�O�j �_7�K^+_�����I�s��h��D��j d���ꭅj#(�̿���Ҽ:Q]!<0�y}��˒�g(,� ��깶�t��o��!��=�X,Ӳe�o�l���/z�ڋ.@!k$9m� +2{�:8r�@�%�0� ����n����p�Ӌ�@Š��e�ق�_�m���D!V�%|QZ�]�%���[�fg��lY�f���J&��Rq[n���o��v��X!����9J���>�����G�'���4E��VTe#ڶ���AA��;��b"�H�U4]#AoW����#�#�����r�V"Y>T��Ֆ��7K���3����#�<�n�:�n�:���/��8�|p�����D޼4?7۬:�굚ӕZ6���8tUKյ���|\N���D3袇�˺"��Q���	�H��䁽4��s����ЎWPj��qy�c9]��:|N@�Vt�T�-Nk��t6���C+bb���j6C�I��\�NkWRE$��7�@�+�	҇�O�mp/	�x:\LM[����>�O������4��&Q��E���L=A�<���"C~	�x����0{q��;�j��*j&���I�"�Ld՛ђ�ī\	��a�][���K��-s�{���(a���I�n 4j�OO�>9d
-E���;��w�9�����rn@�)�}�����E��������g�����Ӱ48H1������_�y�]���D�G��cG^H{��/}���������������.��7����OE*۲�Dm����YH5����G�;��� 1�O�.�	�u����'��r3�}�/M�h�v'��<;�a�sǹ�>dyu+6Q\�L����9y��Un�X��J"��ɡ�˂H������/�ɉ7��0���������Z���u��E��2��x��7DƊs�"�̾D��'N�h�L9�PLr��k��f�ر ���J&K���^~[�p$��cih�� ��;w�|��7���xE�Р_����e:0"��I,���YC/fzzq�N�1>�|��_��4����!<��SSO=��W�@��Y�˙,*�B�;�k{��Ѳ�q%=o9)��(���E��F#y���[�ւ���k(���ׯe�����?��%��9�h��x�̊t*���@�l&z���Q���:�x�Ӕ(I"x�@�@\	�4�33I+d��C�r���ԉ�ҡk#+�y�'�b�}V�Uz����L�]&���:*H�wh�VM�<XiA�d��hK�a�q��L��CQ�z��?�z �:0�3���2b���Nr��HP�	��3���޽{��
��f������@���L�[&��̌3���O�md�h�0םs뭷nހ�F?"c�4U����t�g�,�<�ת�2��F�J����2��ׯ����o��9u����qN�+65^��fH#l�d� ��kZA�h��ΦM��l�@Xk�ΏA��D���W���ۨd��3d�S��. �+�	���G���<B_�����r���-a��6�v��J5�4C�����c������@s�D&r����
Q�$�!��B���0����$g�8�ʏ��0z�,�&�i�D�T��_��M�K"�Y|r�y*l4ٳ����"S�� �m5��pdgfk�4seZ�b�T�K*�ɓ�A6f�Ș&}�r�����!��wb��Də��s����9�ٙ1�r�����}�� �kȨ���>��o�1��>%C���o��=�yx>h�Yas2)�m��s�4 
�aTɒ��?�p�/ぃ(a���Yy�M7��?�c	�R�7�����K�N�H�!�%A�ꭷ��}��G�}����-���"�@�Y>���B��[�6
x�z��EJ"G���JŲzژ��V����'Y��(���1��xA���ee�Eb�i����-�o����z�[���O��_MMMa-x������7��:?��{��ڵ�V4�uk��֢Y��*80�}�k�2��$� 汥�����f T����""���������y���d� �\����ֹ���Ǫ�� ,�瑣A�v�@4P!_e�uK��$�a�1Y?aE�T�E�T��*TAb�آ8�z6$���k��3Vd��A�GE�eg5��A����Q�6��'Oq/)�h O���(w�LMVT��4��)�zq����9l�[��S��B�*�r_,,%A��0i�w�-E1mN�Uk2_U��J�cS'�"l�dd�$��U�0�jئ��nҲ�{�&�Y��Ik9�ld�y6����n����k�8�|�XԾ�z��o۠��vJ�6S6H�"�%7��f\���J&�
=�W6݌.�~,�V�	�-n�4P��~@_F{�����º�SSO7��'��`�E�}��AH
��[�
�R��2J;��f۔��I����u9�A���͂Rq���~��A��'䅴\5�a����{�-42snp�y��m�Z�L
�m��l<~p�ᱱ7�t�jZ����s�ȧ>�)! ��&+3��ey`I�DD���#�`�|H����n��#M��4�(�Ԕ�j2*���|7 ��-�0�;"3�|��fL����������|Az�~_\\޼y3�B��I�(E"��"� �#�RV'G҉a�\D���5Y
�G�s�,��v�A��|nU3��lB��q�B!�2�ť�u�0N���/�5c�c�b�B��M\Bκ�e��bx+��[�ޖi�ѳCā;�g��ʳ�8�N#Iޏ��B��믧�ap��ť�F��c��r_�������	([�XGK#k2}�s���Fn��V�9�c�+��a�#%J�}����[�䒝t٧g*�����o���!����e�kF�,2Æ��<)ncma$�k��m�2ql�>�8_���^�;57}��*�y�%^46ҷ�B_�N�W2�A�5 ��b�'�M;��%�^�I�S�2�������ΙCF��MU���	 M���Je��v� =P��S'q�dMK��R��'2-���@e~1��ټ0��Ǥ�aUx"��8�]3V����9\e�nK�d���,q\���3К�j����AB�5�� R��o���2VV��C��\p�y�Z�^�+��ƌ
t@�����v��@2*���'�Q*eGF�6Ȍ�Wۀ�mD��&�	��s�n�f�;w�,]���'�Aj��n)�L#�Y"x99��X]�TE���Z�㘈
FO3�	f�/��Y��C���Eg&&2DE7�� �J���<�^���:@H���ZO=�ԕW�b���nĢ��mo���}rr��Y3C8A
�Q�h�C���4����>��e����Lo���TµA5� �Z�뮻���_U9%2H�j�M65�C�����$�$�[��5�\�w����w��m_��w��	����D�E�5�'���A�C%�p�t�,�N�G�M��v��nٶ�������u4�Dik��a2|J��m�ta�?�O��-oȚY۝%���������_?����_)���Ck��½���_��/ɑK�����S��������ĉ�;ο o�)����Ǐ�zܲe�"�u]v�%�������7��z��<[?��ƾv�W2��뺓 ����e��7���o|�%�i�3�QG���:w�;���q�ƶa1�BMC�\/���Gҡ��ZO����N�,�k#\�y�q5Iva�T�p�A�z�\�t!�(N ���P^MY��{>�,�@f>nz��r8��m@aU��=P`Y��~�io[XX�g�t�����_r�n�FF�?k,#�3w��c�=>d(���y�Z�"��1Z�[�*x�!z�ځ�����ȅ7op���Rߕhݔ
k׮}���ޱc�2�6��P���!a])%�Įw�D�P����L>1���-�f�^���;v�'��#Ȗ5�����&�l8!D@�l�-��0�*����H%�S���*U�fz�R��Ǐ'����6l��Ɓ����ly�^�2tY��
�����`�v}qB��p���BI�7r/��޹X]��TP��
=C��t��'��t�=ķ��c((˧�t�b&�!�L�O\�Db�3�+Ú�h𣉭$��"u�m��GP�#���(�Q��yw��dY>k�v3*I���aOK���D��%�@%���?###k�3'�.�͚T1������y���ѓzӛ_�m�9>�A�5Z5�}}CCC�O�F�ޤ�6�A^Y0��I��*榧�������-,o�	J]200@��5Ӹ8R˜J�۰��pbb�����y�{�[�q�,�1�) �OV~���GO���\��J�FN�����Kw����/4ņJ���n#!j>Z��]���n�(���'N��Px@�P��?}�S�h�����T��%�Q�t��4�����|�\�5��[�	��I غHT��Q�������:�ȶI����,wԉR	IdwÀF#�YJ���>?=E�Yk"��\��ܔ����|���_���qH72R.������	�<�	������[��HR�j���:9sb~��~��Ν;5;K����Ȗ�z�w%a�?K5V���'?�X!<��״��|��_�2�*�y�k���/�;ȣ�5���	������>����,��H��3�y�[n6E������?�_>�g�������$6/❺�EX�(ץ/"�E/�p���{�)������������y�ƛo�Y���?�~�x���Ç��|�ּ��|��_��{n��Ƅ����M�������s�k��?�A.�T��^�J�j��2�t����G>r`��w�󝩙����+������>NI�^�P�<o|����/�y睿|�/�^}�����~���Ͽ袋$#�`�]wݞ�w�����u�yE.c�w�0S�ݻwbb�7~�W>���&6;���Ӧg���\C3��+�~���Q�����C�
o+���8���玟�P�(&��z�;YDB�Yv.BW5IU8�ⱖ|$�a5I:}D"��JY����ѥ�:�[dk$���\�i#�׍�1:�b��z�����B��G�"�W�7��Qi���ek��y��&]Ik�t>�;E䴯�?)����h#�mt�u:����C=D����׽��=��K=r��1T+�/ؾ�����/��~��hr��\N�H����u�I���r���-#��aB�J�s\�>n匼M=�зK�Ʃ��j��u�ظa�ƍJ���$E7��y�0
dM"d�t����C^$�"z�|V#��ɨ�V6���Z���?���{�������� �^_�[�q�q���d[74?Ȣ'7�5�r4ڒ�L��ڝ?P{)�t7J_��>��sR2���;��ʲ�+U*��F�<l˲��}�qQ����]1�a��CUm.����(��/;4����4.�I�Tx�.�B�IL4Y�V	�G�pзS���rp�GueiyAȶfݸ�)���~tv+r��?PDL`n I��A���r���	͍I$X1�-�)�K���%��x�\Q ��H��j�s�T�v�}I=]�E�R%��y''�}��I����\Q��8���%,����c(�lr�"Ў�@7�>MS��@�Y$#��ɧ5���F�Nc8��\����=h%�T���Vb0�$�����: ���lX7r��;����/��V���0�D�3�qm�GJb�\j��&��p��"e��6]����^�$5jRX�֒jؚ6$��j�k6O}�ˋ��b��7do>/�A�6mtpU�Tb���,�R�u��3�Η	�uzja��ڭ�-����eӔ�X}�e�?;LC:;3㹮��~�\�R�l���a�MX-v<�4˥��1��Z�j����%������n6|�_[�n]�W�-z^NEc��6׸CA)�	:���'3��� ��pMMV#�f��+��
��qW�@±��oڙ�{�V[�X�t�����3����������\D�#�}�΃�H`�@D�Bq�:�T��Ã�|_M���4.TC�⩅�hv�<h]�����Mv3ӗ_�Z��݊=7r9�b��%ĵ��w�lE�"�HT0�����~F?C-�`�:ֺ�-"J��"5�-7�J��/���m�ݖx� 1m3NµkF�gg�|�/�{�{�=�.�E>:2�
�vWdht�'��G��O�~���+��ôJm3C�ﴚdyhUJrt�;ߡ�㮸�n��xz��c���~�Wv���+��k/{����굿���|V}z�>���s-��z�ۄ���ޛn�I���^r�����u���p��v6�������t�A��:u���B)TL쳮�uӶ�>�}]�dI۲e˃>x��5#����uϽ;_����v��>;5SY�����M�O��U׿J&W��(dբd�������|�٬�ȝ�2���/ܫ*�+�����)Q%s��G?�a������7~㉶�D����\I����8������!D�/r��k���!�ݝ�sN�҈}P`����5I7���>yw^l�~KU�=ݾ}��M�4�Ggm�aoE>G��m��hY��Q
�����je����?�[5T�{plI�d'��<����M�/�cY��v�ڕ�����R]xᅻw�&��w�!��p�\��[oݹv��SKK���v�z�������NIz��������B�i�X�Z�4�	�ۗ�6i�]x��»����-[��Y	�@� Cc��ڄO"�[GL�4BS�t�$�-��_%��u����Y�۶П�<q��:g�"��(u�)�Lsnnn@��ر#+�O<�� "�fi$��:V9T�)&�Đ
�}Q�#s���AwT�):���pee�0�eW�,�?���g���{쉃��'�fs���~�߄� �Y�1�H F�))����N.�w#xBv�(5�i��`�B< 1��!�H�5���x���� �Ĕ��?D�h�	�"��M7�,��v�������6�#�+�=~�a�"F u:�%M��T�K&|����ȝ����_`-II�,E~O���Q(��?s,1LW*$bĔ �����DS��ƥRi$\155511��\)3�V�F�P%:�E�m��n�8q"�'''�)�4p�=4�d��=033��׾z���3�������%t�;�ɓ'K�׌��`B�q����L��oȽ_3�O��Ϋ�=~����S"s�^B4u�;���aZˊfЧ����_\���<jA��� m���Zb@�V�---�ِbB��)8<_z���>��㜛���� �Se�Ƅ�Xa�1��Z�>Ex	��G3�X,�Uktצ�C*���Dʑ�$�IG^��_�m����E\��U��(7f�%L��3��c�E$��u�:?����o۶x۲�򖷜>}��>�30\X�T�Ї~;�QpɕW��}�������`�����h�^���"�~��F��ٳ��{�x��)�R\)�l�Hv�����;.���_�2�1����|ӫ<.�3�Ҝ��e2j���g��~�x���N�Ȗ�#""����i��4�I���v	�sZE�nl޼�P�� 50V��ȋ�u��9�������J�uˊ��k���~�o���?��?���D8����/9Ҥ��qG1)��߼e�]���*mi*=����g�{������e�1����&�x�W�x㍟��?������r��=Z?���������n��w�~٢Bn;�� 1� ���L4-Kv@#��o��?��7�|�Љn���׽�ud���js�rB��G�B�;�)iW�9�s���P��ֿ�#~nZ�G�t���'�(�OEJ8����!Y�h)�K�l�1ycR���x��;�Y ����qvU!V&���'��Xi��Q7�ܿ�<��:zb�24I�薺�q�u4�/�MxiGD�)��:+������lf@��Uk����o]p啲�׿���a.Wk^�oP6�7�]�Zo�]��n��
rs�� F��*)�;x����Y�V��"���mI����,qU��������Z ky��@q�3��7�04�.�eK��_�A��C�i���Jb��b1{x$�I�B��Kz7��j�O�|5pm���0�45�3���Uo�[�]������r=̵֖L�0�D*��:�~�KJ�ud~*X�:��Z��noX�j�Z��c��+��Թ�3�x4�9`=蒕Y;04V�oa[J/VWbU�Z��y�3�Y�fϑ����7�������d54D�Rw���@�&lW�t�|��j�g@Dr�bli�9�@(��la�M>����Վf]W�=3❊�0��џ�,�&G�������iY��!�A�:*0�Yq��c$&�d�Z���J1��K�j�j��R��!����[D���@h��l��D��
m-U%����0�J�e-��:Zdt��9&oFu�[�0L/�]*[�lnh`0�����CB˯|����$��6������V)��O~���ypR��Z�:Z*�Q�&g�m����w�8]���c���L��C�J|����/@T��(�Hr��V7]|�.Z	�=Ǐ*e#��`���c���Z�<=��<Y�U?�W*O�=��{�T�h�|s�����4����	פ��)h"�}9��Z�z���v�fb�P.�	����Je�ݨ�%q�^
@kA�޲�EQ������s��i�j�2��Q����Y?@j�V�^��L��� �Nz!���
��:���CZH}JJG�2����D��L| y�����͒���RP�'��>Z��z�>���8P���O?��ͷނZ��E�,c�֝���W�� ����
�%�w2U-v�ÉӳE;;5=o)F�X��[	���<Ff���	���M��7o$/�Vi�8xliv����#���AN�Q�������x�b_㬗*���B� /�3w�TG�97J��iK0I�2/�P'�)JN;Ngӛ��23'�?6/O�t�ݴ3�k^|ͷ��-\��IHD�d�'C��2_��id��f�4�r�����7t2ྒMh�<�G����k��O���1�@
�-C7hw}�˯*�JG�Q%#��\�`薝Ց�����"Bʺ��}�� PqʹQ(I=s~���3��Z]���}�C��X��j`*6,I"'B�6M\��j='��>m������}嫯}�k��Y�]����@�ɽ?_K�����}�%���������/��b��?z�I3�y�+_��L���:�^zJ�|�K�9��{�~��7����8:9���F/�u�f�j���v������� �큦׉h�	���g1w���8������K^��!}9YZm�����/�3��PdE����gz3�oH�HA��K����٩���6�O��Cx�S]G U��H&���K���.qZ��N��C1�pa[����b�кH �$�����a��H��7�*�"�7??O�p�ƍ�����h4$��*���S�J�>N�A&�M]^^�1���E�@:{u���i�Ng��t�x5:���Ţ��!�5C�_~��-[_����J[h��O"��|7��1Դ|�4�@���,�GKJ����?P�+$��֭۽{7��j2�c��Ǩ�H06˃� ,�.��2��I�R�o�묷����יe�Dw
��Cbe�,XD!����Uk���v6KN�޹y�8a-B#�͛�k+t�s�s��&9�,���(E��E]\� w��𙛛���!JҖ-[p�b�P�Y�1�8]���*�5EeA-��SԦ���MU���ل8/gx��g�軀g"e�ZMxY���t�R	Jk�B.���:C��ɪ�g���kA�t!�����,�j�B�?���SX;�`�����`,��#F�2��11D]�;q��F�C�ʋe
K�V�K^�뮻npp�^�����:E޳�,;Z�M��T@5�ɕ�t}���X3D�~��qz��ˣh]�͖�B���Gj6��5�so��]�Ν;��O�*�N��$�@��'���o�l1���u�k�s���7�믿��4K����B��o�X���Q�����~4����C��E��_���4��W������Kg���86���)�� ��V$������/�J֭�]�ւ:����E�.����6YY(d=+Ѯ�H�I-a�;8-%�:�}���/dN���J,������ҽ0z�D��o|��׏����}�׿��Эa�U���Bz���w��=X��瞞�����/��Ӌ�k׮ݺ~3Y�z�J��[�\JE�o���^Z*����ᾯ}���{��E'�j?�?�謠��g��J���r����ׯO����d������Ʋ�t��i1��q�(�T �h�����tｯ��z�6���@�M�2�ߎ=J'$-�Ob�3�'�BZE���fO�<IS���cǎ-,T�d	��4���������00(G&]�?��	J�D����cY2�I�1�n��v�=��x�H����P�����77��۶ӌ���@ݸ�|�󟧏����A���c�=&J�i��mۆ8�aj�3��SJ�Is�f>-�5��4�i-_u�U4�"�MO*��Ѻ�D��k��=`���XQ%����sX��q���G7�-Hx�Y8�AO˼� �Z��F���V��g��,��JJ��I��B��?��0b-#�.�7i�s�|����֑���seN/t1�ܡ���F.B������U�����#2��ޭn!����"��*2����Z�(�V��C7	'ЎY��Q����?||�;�-��§����#�,?z���Bry�����Ld���FɏI�F��&1봐���)��<���Z������/~��~��G���6߰sA�I���0y��sϥ�a�9���`Cy▜؊d�s�"�<Sjx��IYGix��/ؼ~���b�k5m'F��\򴴌�d �8������i̶lr��Su�T��/D�<�A@��)�È;�������rSӛ!��	���/7�yU%/�#�h�+f
�X��=ʊ�֛�ߢs꺩��� �*�WH�r��r�&�J��)�c����t5�=���OE���84đh��]H�5�����J�<��(�糢�Q�S�dQa�K�Dx����8�)r<Wk5u��JU+E2x�;���9���?�PV�Ģ؇e��^8��(�H:G�v" qg���b��S|���lcn{rp5���h��󖩫 挂$��?�� �D}�(s?�2�W�{&'�a�}#��;�/���G���Z�F�"��hV�irA�f͚��JI!cҙ�
i��J��m-//5c��p� uѹF��-κUx�I�r�f�� ��%XU�ԅ0�;�����6l�X �Q{�<HGXo�qŐN۴��,ͯ,ٷo�X\{��k�sˋ����
|O�в��~����4��Ǣ�4e2�)g샾r�����"�S�L�&����!�n�h���c�nj�mʲ��ur!�K��*qH+�XȪ�Mн����M�E�X�(�cdK ɰ�H��$/V$U�~z��ޡJ��2��f{�0زG�l0���9^��DL%��K������������o��<���9B�v�xbr�_��<��^�TRm�ar�b9��u$%v�VWB��|�����鹗���׼�,#y��Y���������}w}�ȱtk�霉��|�P�®�������`�D��Uۄ�H]�؇�����+$�h�4t�!E����C�7���س �������
ˬx	�����ᮻ�W�9���y��B&F�|tE3/��[��?H[I�,���BT��ޮ=�o��͛�\��%����0��>=t3c�ֶ����j�9�v��������5�}��m3����?+ZfL�u�E������`�h����-�e�n�k��&���e�l�iI-�"�ά���^v��|�����nrv4o~�����~rߓ/�����N�`���Dj�����O|��Ҡu��=��w�3�#�Z��)	�VYS���7���oϟ�X72����}��^�7<|db�o��2m;tZK�F� C,�*@W����|���&��s�5V�ҌsX��q��)���i RM�f!���?�n>3�.�rW�EB�4�ǈ˷� 87a���,���L��~���� �B����B�H�FȺY,�C�wVW��CO���x�;����-+��HAܽ~q%ǏG�^7e�ب[j�>ܘ��Ն2��y|� Aک����T7�cJ7��	,���nݾ}���y���:7t�PK�v1sp�o���*�<�BYK�B�^���Fx
tZ��|���	��f���V����%� T_\"�8al,�bț�R�tǥ��\`tH#���,(����b7��1"�����~�� d�c�����c�@E�
ݣh��R���߯ 	x[L����Բ�F��3�=ψ���]s�8f*G��M	��eM!nROoMp{J��E�P	9�I��!���5��:Nsb����0�=�z��Hg�ϚZ�y�4������]�b�ۦ��&˔i"QKU&<#n��s�S%�T��\J�n�`	2������E�{)@e��DN���KYh�No�}v�V��.Rߐe�����RđlvmC8�x.���;	�	��+��.}����
����<X4��I�*|�et<������.䤸�9�L�=��d���7���]�,�%F�UsEdh�ׇ�G�
�zD����R%��FgK<b�A]��W*�$5k�X�a�P�	B�h�R��U������3uww�U�u�_�A$ǂ����9E�1j7W���-+�|���#Gh>�=D���f�!���<|�^�^	���U�;|�&�	U.Y��a0�G�a�dsh�+�U`�o;���h�M!��s�Ή��س���-I��b�]ϵLr�M7.����G夥d�������[��b+�M��N����@�����Ix����{��V^�fPa!���)��.�lbb�C?R�D��Ҍ���C��V��f���`__���o���;���'��M��+���7����/�BK!�	�Z���?��1Y�gy��%HX՝�qh0���nz#�T��.V��=9]7c�Ν��W���|����P.'|��[�������%_^�w
g@vZ�l�[�s��WӋ_��W/�b���>J��o}+�_���>Ҭ�s��A�;�@q(���gPU�i����wp�sWn����,��h�i�� �m#.E�2�
�6����}�u�.m	��2Z���-��b�閣�_���-z?(u�����a� �V�CL�Vɵ���A1�P�"�&*+8�^d�ݕ�D#+��Pk���/�>�����&kF�BD�%�?�����x%N������{ht~�G���Ӯ�D��$q��5�}K��9|ī�㉑�J���E�fX����q/p54�e{��B��I����ť�����e)�=�P5TT�s$K���l�:�ich�3�e�`o�4����ю �
I�"�v�n� ���L�I
�!�T�@�+L��D����qm�:kEx����ϵU��&T(��rP�5�vʹ2�%����R���K�r_�V�9֞����#�Q�Wִ�B��622��
y��\�4��H!�&���̠�A6��,f�����7�b!�lG�8�ʁn�a�޽����q.�h�\\�@�R&��Xf DB�'�9�\d�S� 0� |�FCyO�4Kny���8�웖��
m5-n��E�k�_��׾I?��<tx��	��BnJ�82����M��u�7J���S��� �>Vظq�h���^6$��=¥%�t!��7����h���3�pgi�k��]�vm��*z}:
FGG������~)�v�ځ��k������ػ��g?�YI�"?����Q��p=�Mz�������s��+fl�6�h-��gJ�R�ڙvv1�`L�B�9��R���
R�Q4(	�Ȭ)�ai�i���"T}��J���pH��v�UY^�%*�}j�a�0hX�9����Ţ�0Kb�k��%�-�5(њ��W̸�Ԣ�Չ���l�#�}�(k[\���5Ơ�љ�n��"ā�x-GUL��F�O�B %E�?.Z$�kWڵ�##�^{�/��*��=�4����������2gG!JK`�#�H�67<<����{��q*��qS���\���V냃��Q,}Ţ�޿h�P&�3�Q�@�-�Y�(��ؾy�5:J�|��,�}��{��>�.T��FQ�b�q�l��,��}�������t�M�����@
i��s��l+��+�f���ů65��9�X�Q�Cl"�����VNO-�<���Gf@6��������L_KW�P� �>0Bs�V��u4ihj��7it�8���m�P�u�9;�ɄMA)ZB�*��t�NZd%hB�ZmY�>U���2��u�{��5����{h���\��P���};�h�
�	�(�1`�apx��f����Fx���c�F�I���Pl�R��չ��X�⩓����:}��`l�Y:Һ���	����.V��Ћ5� '3PǗ���]4��X�Jj�ܞ�K�Pq�4Zq�^m:����¾}��n�Iw� \�U�Y�Dc��:�ũ�ТJ[�]�kYID�z-���\Y���S��{�Q	��n�Ȝ��� W��z�oz+$ۢ���]�u�/r��F�9s�v�ĭ1����)p�M,�n��j	0bD:�/�k���X���Q��Ii	e��MR��G!i?���ӷ���;�>�w����h�i�7��7��m��U���.��|��Ts�B�!��$�뮿N�d&��
�+��"�U������{���{���~����N}��52ut��߼k�֭�	m�q����O���Z���]��7�|�����[ٶy̴���֗�*:�朔sנ�ߑ��a� ��"����p��&A%�==ӛ����Y�g�Շ0DB
�
��0���ˌ�ٚf̡\�ԛ*��0�6	 ј@��*D�9'���sv��K�}��$��׾��(%����+� �u�W�1��]��\�T�fk5T�v[�s���_���n�����?����z��^s�5d+q�[�����jq�@�k>m�( 'Y\.�Y4�`":��ϛ\���_�'<8��ˆ�����Yod'�B�����Z�w��|���P��.i	��l��l厄�٣32���j K��	��Jri�!��Ù��	_�It�����Y�v��{�i��;}oHJ��b�J��X��-�M������J��J�`��I��z��:�dB�r<[��GϿ��C�L�GO\����f4P��mh:��4�Z�Ӑ^\ZX�6����Q�|q�Y~(A���X2�!٧Z�K�ăU�'�I+�J�{ �MZ�[=KȜF��C?G\���2����T�H��mP�F�x������Ϧ0	b����U��ډ�≘�>��(6��
��|&R�p��F�y$RqX���Np$�H�!Tp��(nܶm�� �*j6�B���y�{��2t\|�T ��u�6���{���K(N6��T�4#���A�q��fq�QEVGu���L�S!-����r?�pJ[(d���`W�a��k�Űє�%^�$%�'*w�
y�$�p��A�B-����Rp�J>0�ZmyE��
t��J\4m=Þ,-�n����_:\9�Q�>��v�Se�V�	�,]ý��Ӭە8�ѣ3HW�7`ҍ�
�}w��Ϙu�"�(k	����M���TH�	f,���Z���`����A�?�*#&ڂy��a��m@��L���e�����*���v4%k�e�)ȉP��@ׄ��^�	4qCCC���C/2�fV�T �d��4��ZYX��A�ö$6�1i���J��S��4ϯ�8��D~$Y)z��Ih%���ю��>QR���T>��h��u��-=����C�ݳ�ԃ�a2�"�Emv�N%���N�l4�-C��ccc�Y�7�lE���7�t�b�h\�o���MҮ),�4>m�	{hFi�kdT�R��crKw�����<��t;�1:]��xF���]`k�/c��K�T�`}�q�%Y>�횇]�VÎ޸i�HQ���(OgC�Ǫ�*D˨1k�$�9�C����V\w2G}�R�4����S�����e�U�uh~����ʙؘ#q��櫊��e�ܧaܱc	������un��6L �V�%BU
�i8$m�i=�XN�vt��Y}2ǋE�������[���o���
*�:9yY3t�]�v��$�1����=���v� Gr��7�q��?
L?�!�}�-.�XW�iR�&��Y���C_���v4;�6��%�Y��H!��P%�/�[氱��DJEn�D&kp���P`\_��^)���C��YbV�Jo1�d�i�{���Q}Æ���w||�� ���^�:�6aXe��D��e��l�o|��7~����w�񖷾9�QԒ��?3��Rt�	�n�4�IZ����x������l�i��z 4Tl�9X�A���f��F=�B�E!vTi��MNH�TN!��$�� WM��{��P��_�t1M���(JV� �A�[�=#`�$�_粤�� ���A�Ǜ\�s~_i�m�Ec�@~���őa6]���5��d�	�:y^�[��3���(�@0q�X��8��<�?�s���N:��o"dFP�rD<G���SD�,�kۡ��e�~����-�i�fV����Cs��b.�3��yd�)&%?0�Z���s+���I�bOi֖O��"4,�vQ���yT�pH��zJv^�R���4Z~S�+�e5R�\��$Tj����U̻$C5~Tu��na��<ey��/fuq�K�|E��j�Y�Ӽe��5�!s��o�@�KP�_�k˚��x�3�fiQ+�Rn���3(���B�k����l��[g�}�ע1t���^���_z1I��U����&ښ��!b0T0w*�el��c��a�6H�������k4JE=�҇�����V�Y��Q1\<����O���N-�\�-ڈa+���`����N���_��S����&��-[F_|���h�+�����GW�g�Ƈ�ؾ�2�Hs7���{͵V��P*䱵Q���<�pRM}��s�"�l�����Gcr���ݻw����|��f2L�`��9�k>�}}}tےY!$+��
;��5ACљѸa(nC�9�nA��Rw<��I��	ʊ��xS$��v��B�s��S�,�lv��"��8�v*�z���[M����(���5���-�����$������2:b����^~��#�Uv�l�V��Gl�������#8P�I��¼�È������GN��
�:n��o}�v����9�g�=y��5 ����W��]Zǩk��i}==f�i���c�䥴o�i�j�J�v�j�Zjse�
t�d���c����;�^�ky�R.�=�����������4+�_t�c�(KKK��25DHE=���^L:�E=�UZ��� �J����it�� ڔڸ=+J.8����?�����ܛ�E��Һ]K���Zl[�c�{�����k��3S(a%�M��B�FI�f.	A��bK��0���D01f����͋�q��gt�^o��-�˴�5(/�0^���8U,��U��m�IuFhE�T�j��T=�pL��(��v�ڹ5��b�&9(>v���}5= 7;�u�F8�9�c�zqȫ����@%k"sՆm���%}�%zSi'�f�N)�i�\5-�n�v���l҆�R��Mᰄ�5���\U�_�.=����5c?6٫��9BMv�7�ٟ�����ܾ�뮣����jyl��#τs(~K���8Т2����0��$`'m��i���o��G?��?��;�8l",1�<SSS���iv~�~K̰7�����黾�]�`����O<:7?��_}�e��� O+�L;�Pyդ��a�n)T�TފĮ�0��>q��-7�?�%��A~D>��ZA�E��b��h��H���N���A�� �jI���z0K��:Ӿ�k��~oێ�%���S �Ֆ&�֫_w�_�gqq�W��_�-l��v�@�!R�X��f���첗������cG���z�l�ٴ0ר� �W5zMJ�L����wi@B����Py��z�#}@?�@�X�
�o��4�P�")vV�#��������Y">$N,�u|\��9�ԓ��ݴXf���-*'�F醍%��]B�5y���l6Q��-�dٛ�O]�T:��NFK
�TA"���{�1�jf�E�6�G&�+��$����a`s�z��1�T���ʾA�<Aݎ�YZ�#^y.��
�Rݼ�I���oP(�rYV���nO��R" ~��s-sz��%��Dpj���B��{7���b�k6%=���iI�I���ب!R.�H��#(�/��G���:���/��!�N]��&����E����ݮ�N�P_��r�+Vӳ7��ϐ�'k`hh�g��Yg��;0 �N���d.�bD��Dk�N���v�B�rfr
��5d��+BxX�kt����FH����|�݄])ԏ0�䬑���"i@?v�X�թYB>!�d�t��H֮�}c�q�$/�ݛN)B�t3`��0�w϶ɀ0���lph�fvim����slG�:�\�u���^E�<4�s���OmFa!�֍�_]�H���tM�?k�A��в��cp(�6K��:��M�:h��1re]�V�u�C�aTU�Ħ`r��Tx'����e։|ǝ-@;�n��B�����R�Z��İ�Y_�Nf�+�R�\i���+4GҌ���t!@,<���9�+r��d�,ʜ|��p�D���~��dHe���8i�7҅��Po#�BK=�8�%v������9r�lMڪ��ꡩ�p�μ���aYY���g�ٚr��3�Kb,��@N	����j.��ұ�0"D�3#�(�=�
 ���{p ��*j���y-��H�V�D��<��
��o���#|�(\������2"�ʦX�2�Ri�1w�����9��-`5U.�Rci^��7��'�1���)�c-ܡ0�9�[�vn��kǾ�`%TY��v��9�H��\^�vnR��E҉S4����@F.��Ix�A�!P�EUO�]����2�hԿߑH�Fn��D����}��+��ŷ��.����7^���d8���W�	�Z���g��ΰ�Y7f>�nD�[`�u�[m��ԧ>��׼���Ͽ�u�}��_V��������x�4�7����岄��<���n�����I��{�W^�J7��ꪫH]��Ak9!��2"t�F5Q�Z�Zn��mɎP: �N>)�뒬J&#[U�7K��I&�b$���%յn��8o�a!�ƽ=%v�p�AUR���y��P��Z��H�LD&����g�M*�'���k�SKbC3�9N����Л�^{��'��E��i��jy��M�.��ۿu7����I�ﴋ�LE�A�f�JA7�0 /?�z�����x��z�C��Z���205��nC�!�u�� �2JM5	u���.lz
mZ?͖���Iˇ�-��۠l�(Q�J7N�alDV����)G��$"	Q�Ur2GN�r����$��Z�Hʛd��$g@A��$��D�'T"؂���!M���\�vPl=&	⸤��Y�QQ�C��b����y����j��GF�H���`>9[�D��Ka� �c����D��XaL1�+c�9}��P|��G�M���Z~hh���dr):�����
U�X b�y�� JJ��Kp�J���S���vo��������ȮUTnY� �9����Zo#g��k���b��@����hp�T�4�H�5�A��9�٪4?w�K�7��l9���m�t�E�V��5���ZS���hWP4�WX��8���~���ǹ8�K��؆i�IQ���[���_��|�����xtqi``��PX�u��B�fH[�c�J�[�$!�JV�����X[!][,�tK�V���u󓣣�j4�p�IpU?|�g��]���n�O�f��a������Xk�c�S]�R��!X��iX*ّt2���_Z^��I0g�y��՛�0��m�Uw?�����R.���s��
��n>Q�)�e%&�p�ZG��g�՗�sU�P_�җnݺu`p��γɭ�� 7�DD��#��/��Л�����#�8�{��xq5E����.ۅJ�ہ�`Z�t�j%�X��K��F��b�3
f"}S��J.���Np�W���5]��N9��
��:6�8��%�x 54u��:Q#�{y�����9H��^a��XDm��t�ע���@�)�x����P�5ɎOyCEZ���+�ͻR����[�%@��4�%�{��_~������с����r�u
���f��ovM�ť�6(��`.q@��ny�>J��幊j7j��K��MZi�W�p��=��t��ۓĮ�::3����s��{��Z�I<:2@w�� o}my����e?99AZ�<A2ձl�X6\�"r�+8
���K�`?�ݨa��,ň$�]��w�������w�t�Z���a�F�Y{�� ���Bޥq���5�����ѱ��ni����.��l�j�N��]�v��\`r5��sh/|��6�矋�Ru_^���3sÖ͖����2͗^��Ks�A�Q����\�/���q�R�jp4D83F��Y3�O����|y\̕sv.ѐ�m��=����ۏ���Q��5|· �\)�j'⮀� ���5�Q��R�\PTĿ�\ ����w���j���T}�x-�A�I+��K�AM2�[�&Y��K���l��ՔΆ��f�F04&�ڍ߭�$��z6�&3Bz��/��7�q�+_��]=�2���ɗI�x���?�����$�>�o	$�;����F$ �� g * 
���uI[_�˾q�W\q�W���D�.��7gQ������t=	�6�D�_������~�c���>�'�d�������y��$��Ԗ�ra[���j���d��X]���ʖ�mw�l2��ĲD���$��V������j(��|�K#�2`�}N��FK��.wEv�S(��#�֛��)I�ـ�/9�N��l��:s�����l�u׾6ږ[HU���d����bo�μi�F��	�zS�� ����׮�ox�n���7���B��Y�sW���|"��0�e��ѦA	<O8:Oʀ!�g��q�|��>����2Q��e����<�����n0G���j���馛���_Itt��ꕗ~���D^�ya.�M+�3�R�R�B$��t�7be��#�Bk�Ȫ_r#���ąܿ��r-��Hm�$1$��"�v�\���>NW��W����鋟��k���!�4�*I�}�}��	i_��������zRij ���z����w�Ke&G�.��'�D�s*!�C�sssS3��C(����z{K��z�w�����PS��ri���D�.��؍*�0�|����5E�zHs��$���+着�#�5�<�B&�#k�<P�*l��Q$�ɶ
ܫ���\"a<�m,zMoNMM�9�Z�zzz�n�tI�������@vYJ�d�ڤ[ �tS(���۠�;��3i��Ry�e������3ȃ���ҝ���d��t.��j�~��>5ul�^�;�P����(�)�� =�=Џ���t~lr����!�Y|\���#�<b0���R�4����P��{t��|)S��c��NȨ�o�ǎai����4Q�-_����/��k===uN��9;�щ$#�J\�H�XĬ�T���<+�+]��=�n�/޾�,Zw/�n�TRy<�F�KT�Ę��T����e��
(ɼ�N.�#Jb�J��a$YC$�8{���.���.ə��	s�l�$ݎ̜�BF%61MifB;B5��CI,sV���A�GF���)A��@��`K`��-����R�$n�L{��8E�
��U�l�b���$��ˢ5$�-��n{�EtK4��MyXڕ�ڊ$��}r]Hmq���#G����y.�svy�N>00P�L�c)Yɇ<2�������:d�Ĩ�������e��8���)�&\�ZșR'7�u,������G�Q����;Dk��}�������(p�=n�!0?*���}xK,?k�ƍ���J���ѣ��jbb��C/2+g/--�dh�'k�n�;�C
�I>�5�L$"�i䈓rvsM`�<�r��H*#ü�*���Jfzۄ�R��1�����i����U�C2x\��EZQd��4�JJ�V`��0E�| W��YF�? �%y9I����Z�����m����Ww\q$�����?"$�x:�#'��.�׳'�=L!9�j jXx]tQ���{��>��O��!^��_��/}�K�B��T�ض�N�ݴq��z�)߼�{��rNҘ97�pa3Gq¬:ZG�K�?�v{�.+�]#���y���'v��^Y~V+�=��x5$�t��R���;9�H��Q��Dǻ���t)l�Y>0�
�؂-�k�ǧ�Z.��m?�M������6Y��Ĭ��t,x7��^��ɴ����w��-�x�����ɛ�K^BZ�Fz�Է�F��_��_x���g+\ ����Ï|��ൈL	R4|�'V-g�#��O��g��c���OU���������5@�Ԍ��o�~�+��ڝw�����#�&p�(,�'��.�/s�N����@�i��@� HI�A[EĽ��g��|��lS���iS��H~Y�	�cH:} Q% ~s�E��>��O<�;����Ы�y-�QJ&3,[ j|ٕ/'�?ĴHO���;.��%�?����e��ty�O��RV�Z�p���̆T��K��_��1B��$w��Vc��M{�i�6N֓���Fl�ˆ�O+�������l�� y�d�%��*k�0(����
8���-d���H�b��T�5y��,[�ف�e�U������V����A+���
�<��F=���[�:>;ۚm>��d�z{z��k�:�o�h��{��++�
��7{�r�VUX�[���6P�zEe8\^YZU%fP�֊�^/����a����b�U$���5P�҅,�|٫�޶mہJuϑi��XOR�z��	B%��\.�dN�9/�)u��_5��"��=y7
ڞd�P/�����ʞ���w����t'�9Ču�1���ZfM��j�cǎ�ο���N4`;��`��`/� �fD�oT���xD]��f͗IC6��=E�Y�+QHI�TH�Lشe�VMOU2�5�!�0��ro���je�p�[YY�OL�Fƪ��յ
M����O<��l�}���񙩱��Ri��cǎ�璒z9�u������>��C��u=χ+����a�cߩd�EbC�m����dϿ�5�1v|��襰X\��iz�e�
�d����`.z�Q�!�d�# ��h��RG�S��t6w"����)�@rE%�9�!�Je��$��	#�貆���h{�~��/6�,;JՖ./W��Ia���N�sw��e2�&H��ahz1�h~����Ѥ�ٳ��]��@��L�o6=zg,^��@]b�� �����Z�����-�V����9�մt_��h!�����k�.�����/,�^�(3O>��׿���[�,k$�Ҩ��px���͛�\ޫ����xmE�B������}���B�w��f���1��&-T��zi��U������wD7����_!)�SF����G0�A���c���Ϲ}�鯾������P\�Z�C[��@ټu����.���=[�8k˖-�gg�����hX�:����q�V�w�w=:41v�y���W*���Կ��ٙU�Q�E�,�J%d�X�h-�r��,2j�0F�D�i����br�=�ۀ��+�+�z晁#L9��G�R�&
�4�6�p�g��ڡ-����fq -汏Ջ@���[Ur�E�9+�78`ƈ�T뭶���R/�p��)�+��}�ڜ�)8���&?�=_]���ˁ�`��o�hu��²�H, !ڨ�c]r�Ŝ� ��G������1�<�v�o}�;���2�hx�i�*���g�&t��lk���������Z,"1i����닒8[%��Ӭd�uhp$�!��A�2u��kӰ��`��c1��ϼb�'еx>i�.U�ƺ.��KpJ���T�Phi$�%�P ���E�@w�i��Y�����s�3�+Y_1����	Ր.�$��ފ��np�(ι�Oh�)hhF;h��Ȣ�
�m���2D�y����ǞPQj(�{)�Iny�d`&��0B�R�s�[�{ 	�]�7��l�U�����Ox|��'�ի���׿Nj�����H9w������;�����H$;�O�s�=��~�mo{!�╀)P�̞�4���C�Yt_xf�.Q��4�IY������IF�G���ـ�#1u��U(���K�F�v5���N��bm��(��'?Ig���?�O��}���#W��ul�?�7���m�0���r�9;ϙ=t�=�y�w������>��0�m�ЋQ�?���\nY�w��ΰ։�qh%
f�!Gett���܅��������M
`um����'jh���d�P����
�j���8���P�1G�WH�c�@d��^��B٪������׮]�x�j5�o�*j����?,/-еf-/��N7��
\��Y>A_д�Z%K��/޸q#����M�69r��Nr���U���V��h/�����T� Ӥ=|G�a���W�:��P}"}DWl0
�q����H�3:��>�$=��v���m�7�^m���G�?���N�I�0MLAh�uI���s��XlϜq�i�Q�h�ŶZC\�|-�,� �׬��R�i�����w�l+�8�[*!��uA� ݓ4hd�h~����ld�?~�6W�O��+�:�GF���̡!�d�p��a����s:��̌�� ]��V,-?���@��83��}:��$�B岴��X��m�l�d���9Ch����KZ���$^Ǽ*���z<IQ�]l�rr�#N���$lgș$�$��4�us�7E~���o��(���C�O�Լ�8���m>5�e��y���x�tM|�N���X�Q�jm����X����+�_��;<V��J]���?Lk/��C7GW�H8DlE�cߙ��� kè��������K`�>mz-�K���\4�A���aYc�Kʖh�c?�8���;X�,[�Nggg�)i�bO�;h��o���.��Yl �D��)�i��_�����Z�� -���bqG���ٲeruv�����
�Ŝ��|���x��U���3/�讻����Az�b��v��K���_��vl>��Ϋ�[���i��޽{7}���΢�yꩧ�9�x��Ӳ�'rϾ�䃝{�48�+�R;�,�a����Ib�x�F�JM�߳ca'�U����m_F8ˌ�Z����
��XȖN(h���	�;%\�Hf��'A]_� �Mo�x�7�=�k6l�����i;?��0��׿������\�yr#�ߪ��[~z���y��#.��e����Ȣ�H�̗���0�0��>܁��Da4�z�]D�8���Pn�R[!8�X�֥+�*��/�|P݀]�Yuܡ��"��,e�N)����"a��~@�Y�H��n;+��J��Tj�������&�VL>�K���
E����}��R|K�D��8�(��z�)���I��4����2S�ߪ��:�F��Eq�]]�`�썋7�콦Q��\�VF0�9�;c���:CC7��'7��"�$��C*�m��if,n���l���?^��`nXE
G5#����-��֯Nl�|׻~�K_���߹ﵯ��h3F�+7�k�U���8}���j��}���K.��K����_|�j8��Z~��lN�_IlC����!#�wrh��1{-�Y*�D���mQ���A�	�@�ӕ��/P����y�-�q�2�6��[���K/���~�������q�]oy��8�\���o��M�S���]��z�������oڳo/k���o�S�v��?'��=�0;ғ�`2DB��������H��n�v�r�%�VM'���J�A���f��웫u��L���^�Hy�u��׼F��2Kg�/��n���攙
�=A=�@~1�
H�]%��
{�-�"N�|N��#㰪=��[�&H%�������݇�V�*�3ak�U$~��HJ�@�;p(���<Rf�q0�̹�]��'��F+��b��`�������j��z�W�:����ַ��U�'�g[9?ז���=6)��M*a�	����M~c#"��]C�[��,{�Z��F�wRoV�@*#1l�i&ӵ+�*��$5�Eäs����8��v��6�ۻu�����C�����o?|�v�`hL�C��,7u��z�G`�
mY-��iZ9r�<�#��oa�C�@��a�W�W�6�|�d��n3��F}ei1iT�~H3ىe�d�FOV��1�?��_������<�^/�sEaue�l�P��f#L�����]<00���1�V�����N;�4P/��V*����gV��M�lt�d\�.׎@O/��~���ȊH�uE��}�.Kx%�!�v� K��P�/��g*,�H�tz��8�%���vs`,�9��HwN%��Bh�����A�,��z2��(C�b$�l�/�t�$b�6�Ls*�G�	M��r��� ^������']�L/��7�-tuBL
�#�՘�&aH���mZ�d�ؖ�����|en~uye�P$�A�����s�m��7�����zUI�k�S�bb�<˵J�noܼ=���ٙ����'�F=����Ռ۾�i[~{qey�n��:w>|9���ְ�zN�F�spzZ-惶GN�����h�P{ư�r_	k�KZaj�EI2 T���ݎ�b�	ٓw�+��j�Rbw��f.-,���7�ɱ��Ն��K�����}�2s�\978���\m{Ên�-��=r�����ǎ�ʱ
Ã��:���+�����}��Ka��J�Vm6J==�6�6��<E��|��n��J}�G����Yi�e�&_K���N���Q`�5�k�
߄�G�aĪv4�D@������(zFGFs�r�����Z2
��6Q�L"���!2$%nR����+��)P���̶���4�SD�YȮH���*�ּ�[H?Y�c�$*�9��*��U<1��s6҆1�b���:0`�&��Λ��`�chkf�X=0*�L�J�]��z�)��1�h�Y$_�dH�NA���P�,�I�M�
�NU8/ة�|�9�7P6΂B� p�P緸�4
�[Юt�Ab)] �T�Z^��k10"U����@i�n����az��K*�gmN�s[�$MĦ�vb�)]
)�xwVt����GP��.2�t�}rZhv�WJ�����Z�Crw0�*٧x��X<��6HA�'�1�B��a�(U�r~;�CF�	%�JE��jZ������8��[	��m�Lݐ�4��k#F��[17C&K�?�;���~��_�9���Yt^��SLݤ��������/��/_q����������b��|Og���/~q۶m��~:j?\7�������?����V��`��,�A�?�c=�9;��j�w���Y��x��҂6z5D�Z��w�/�|��7\v�e���7�x��x5٬��=|��'�x�;cdd�C(Eqt�B��̌I�9E���a?��� gCĔkT�"��8����:��#��*s��mQ�6w�ܹ��*�ʬ.R��笭�JV�l�����W_�˛�}�x�y晓�[��@F�2!-�w�^��E�⭷ުh�a���fFA�u0�傳}����6րY���۴i����}������W���jjvi���Ql,..�g1�X��-�%jv{g5�U:ϖ�a)�=����)2������7��Z�~�ߤ������C������)�"�YWn�ݻ�:#��f	�I�r�q���չ�҉)$��J��|MΉ\���E�+~������������
�7��V*�4:�D@i���˯� #�"��T�Eu��q�*UD@���s���sΡ����_y���NF���az���hGI����l�|�%f!�Bf��\��P+��駟v9���Лg�,ˤ�>
S�_c��b�E�$�3:!�9�_����$������A��Z�j�F�Yzbrz$Kq����z	�<Np���wi�1�'�O${�M4A�Պ���ʊ�^i��T�L�M/�>������-�7�ݮ�J��|u��"�u.ʩ�Py�#f�yR&������|��7�f
@�B�|-t�┅#���+������f!	�̢J��[�It�	�$�T�]z�W��U�x�+vn�N7��#�И��h��Zl�
������O.�c�:��e\ۈ��j��"���ѡ�NNN�q�9PV2���.Jg�C4:Ր�1L�+�ez���]K+M�1Z�E�Q��t+谉��,�"F�rH�����%����ee��͙�&�Ʒ����}�)��(5W�7�s�������C(�Z�t{�\s�O��gW��;�x�;H�u�V8	O!��*/����[������3==M.�˵�^K��Ɨ��e����FM�h�Z���LgH�T���+W�
*Uљ�)恭�{kֽ��zJW���	�_7Mp�*򓣣��u�C����:�5T�~��7b��4;��x+qZ>Ʋ�\�|Z-�,g�u.��4�^3E�mu�z�ȑښO��W����O|���%��رcthX �t�.���������W\x����SY���DA���DZ��T��@/B�*'DD�&yv�D�P��ؖ�Ȗ΅��G�\O��U�׋��U|(�D7+"�$�tA��+]�5��fY>I=e�w�.q��[:����ɞEA> �!*R���rmn�JΘ�RT�%�c\j��[���*3o�
�L؏�'\�wF!��~�j�6]�uL�������A���ٝˊ[dx�>ߏ|��84Ԋ��n�njJ�n������{J��ۿ���o��3����.]~.�2;;��\���K5�Q�F5���㳶m��#G����n�M�]m;�~Ù���Z�X�M���>w�g�v�͡ y�$��=��|��\��׸���\����������ec�j����]��/���u�ǿ�k���������<�)z��/�N���%�'�� �Oň���Èm��Q���b~ ��bp�����޾�R�t����b>є��
��L�Uk�	���t���槎��4�L�l�/���~c��k+j�^�T��k�~�خ�"GO"�d-ً�����w�޲S4��d�t�hj������`���_[��z������,:/U�WtE5�Y��WG��&JJLN�fizo�����Ej{�2�w�|�k�s
v�mս�!kr�v��?���\�" �mCo�#z��	�M��m:�.@^�&�Wtit	-׶ό�6zc��q��G9�oE)l>ZR��Z�!��Dq�G��ƉS*���u�Q�8�a�k�r�]4�'�����Vo.g����R�Mcj@�vrsE��֦��9e��������J���������։Mgl�0^(��ϫ�ր�z�zH��@���hmY� ��o�Iu����JX3u�㖩���*� �5��bޱ��v�N�ZhJ������q%�@�]d"�Zdz6}�>��[���>X�=���O��xV]|���D�)�;(��T�!&�Nr�x��YwJ�W�yD��^�f�HJP�UD�Wp��� `�n�B�`�u��(Tb�T( �AJ��+zO0IcP�;�e��k��B��1㑘̰����u�EO�4��w�l��"?����!�:Y*-n���u�vz�ef��S�-�df��Feiq�@>-l�v�N��s���j��n4�$�E��mv6�7h:��i���VQXE�^o���z�0Z\�y��0�d ��`�����8*�K����'A̽I݈��Z������@oO�RGw�\aqq1ܹ��u|z����A�X�n��j"[�H����2rL�P�ީ�i�MQ���Z[W�^���+[���[�}��m7:Mc+#�	�p�6p��؏U��K��������c�w�T��]8`Ǫz��Z��� i�[������S��f�y�@V<��r�=�k��{IXܳ�\3ǅ����h�c��?���mMT��3؀d�G�a����^A����`\����r��8��2��+k��J�p6��������C��5xj߽��9x��Oc@�=�F�P�����Q������[��9}]��ᙹ�MuFFF�m��y*8nUr�J�yZWO����J@z����4�4P��� _kna>&O=\����Oj�E�Z���꣋��ɴ'zv�TM��*�]��-��	s�^SN�rk\>��'z�dm��q�RR��?��J�h}�s��S�?Nr���J
�"���1�H9�op�/L��%{u;�^(���RErJ�����M�H��,�U��De��m�#�Dt�u��'C�V|���FQ��8h	�i��B6 �XZ��ޤ~/��
�!6�1��/g��H�Ph�`/a���V�K�5k���|+&^&�C���y�����2�ϙ-�O?^���0J�(U�>>s��w_q�U6�}����_��;��y���0��2b�)ò�V��C�����l%�?�X�)'�����.�u�h�Hf"Y{��{�o��o���|���>���v�5�\8P��/��СC!�b���o��_>55U̡G�kz�w��*?�T�����o~�uz��oJ��nn�w��";�'�h�h�%��g�-�[��H����Ee5�P�޽��${Q1-L·t�E�\4>>�H���?v���O�Z%�*�gD|K�Tf,�y�l�$a�\XX�j(��q�d���=�\����aE�h�K�)��+�1�
��f-��e�*���9� j'O>�dЮ��ef7��;�:<x� ��{}��Z���G�F�BJ*�R���*!;��Mr�>�w����,�q3Û��ɕ6\?�w�\��B)K�4A�����K���HZ������
7q½�8�� gɶ�*�����)��L�E���4n͞�����ۓ��|�W��4�˳�vn�B��±��vG��<=e47s���Y��bh1a�"QOZS�0�e�:(�3Y4yL�^���(��Ë�����ٿ����j��^k���5�Z����qDC���.>PF^��P�r� ��4���:���ٮӤ�湆$��1
�\�t���Һ-��N�o4D9oݬ�$���%ZonNx�۴n-נ1���y�]�m��\�<��gp`����Z�SK�Y3:=��W4Y4qjx�m��!�#���̣�(� Kl8�H�F��]+�c��xPX� N �x���}�{�=��I��>�G;z���Dr� T�k��D�$��� �tZrm���9'RFWR,�8��M��Z�|k\��ur����z���o��s�	� �u�"��V-_�#���RJ�p�����XҶ4q[P��P=�w�^��i�*}Ԡ�+��2b6l�oڹ<�mzn�Ƥ�"�X�ѣG�`rr2�? e0��i#�9I��i,W贩����a/���¾��id�;�<���7�L��q��ȓ��;���/��ANˬh0��C�hx^��"��ԙs%B	k`�Jԟ>���/�kM��y3��̂m礟}�sΡ�G�/\\4]�"���)a��~h#o޼�����Ç��u��t���5���_��W��{>p�@�< �,8�v�ڹsg�|>�:#��2�K ����ڮB�!I�T\���!6���~�������x�ɝ�N>����N���,@ �C?�<:"��l�iv�2+<�@����2��R��/�>闥"�/j��P��(��h���_i�T�)]؂��%�*$;��o���eG1,X�%/��OD
�&��K�o��}�a+Pdmd2\nx]	�`���8eɱa�)ϵN�w~�ݭ|��8,�T20�7I�~���������w��ߪ��%/>cÆ�~���/�Z(�=�駱�)i�^��v�0S��vD�n��-@Qh�z~��]�߱�&V:�J�D»��L��!�@�E������7�����/�X�������,��7����'ѕ}������?�cD��~�w~矿r�;~�_���Y����=Cp��u��r�"NC-M� �ւ�"[����T�,�L'E98��Qjr-ə�0����c���+��c��|� �o���+���1���8W�=2�P�������>z�����%�+���8��U����hAF�a��$O��Ur�ї�MԢ����b��v�m��N���s{��ٿ��K_�����VDҹ��?�����<���I&B�$���S�*�A�>�A�o�!�0���KO��������j{U�n/,��6��jC�"��顾�6��u��D�FJ�rC[i-
�������$����+�����D�k��q��9+g���]����tu)��7�K�;�	fg��+K$Ћܡ��`S�S#�XK��&���L�\�e������O�9>�W-�Q��y�W\����h'�<4*5��ߺe���{{���N&��|Tx�9��ӳ���G
%.'<��.9�͒�yι��Xd�ԯ�<�5�~�жl�bo���m�Ʉ:td���K��&�l"?����m��v|f���R�m��3�|x8��A��GO�7�3ve��q	�rw��,F�(�Z�.z����t�:Q�d���
o*z�v�R3_K�6�P�Di�$UC���!T���t>����!�̼��ڜ0+C���g�k�C�$�i�=�[Uӄ�3���k^����K�N�VST2�m�D���-��d���r���F��A+?:6 ��jRYo���Ɏ�5�[0�8��:��.����2:>mڲ�|�-�C�\�D�Q*6��%KgT�T(M�q����!�":L�z�飛�j�=�R��8��㽽�k�����P׬^z�=��B>_�Ķf���F�	�c:����11HB=FmdʬX��z�9�ۭ0lk�S[�{[\Y�w`ߠ���E���[��!�;{�+nx���u����7n�[�|��^�2�oy�rda1	|���23]��wUc�\�I���M��ms����և�����84<33��rdϾ�e�y��7��M�X�Q[Zu��˄��d�
G�������#'���'�0�H?�fݶa+��Z]R�
Ʉ�`���yp�Q���iDR�g��#ڴi����}�o.]G�_iaU��c��6 �q�L���3X,E}�j�Av���Rnxy�q�����8{���?��~�щ�Y�5###���Z�25-�i#�I4&��V���Do�PO_s�R]X��+����(F�J1�	��I��'�����g�T=	+Ȯ�*y*�8\Y7s���}GY�O�߈�����I]�N��䔲��J�����A����z*ewaU� ��3��y2���<M-�p	n��v��H��}q���������i����:W�iL��$ܳF�|B.;"���t.�I���jGAJJJ�D$|��4�	�B�c�aN&�m(/�T���o!׹b���0
�Dh�HP[a�,h�H=�w�����d���T�x^Q�픘�����sBEU*����Cd��o$�z�W*a��p������t{������.>���GR8�@[��E�+�M�Ư�C�g&[�kp�0)t� 7�|3�W^���"�@�0/$������������Ӯ�������c6�1�J�馛�����T;i��ig���8�n�������r�DEΝ|���c�Q)�~\J��U�i���K�E	��Ǐ��{%{@��066��\N@����>b.�g ��(����&Ce�m7$��u��tΕ���8Q:r���Z%�LF!S�iA�=��c���<�LrH�(B(�<X�����-�ME����u�JR�nI��4:L� ��@�l@�r�}�㠅N��B�P`
`�,�V'���r$��fQ��������_lur8�h��\�����O<|�]wYM��u����:�(:�[`�bN�y\��ӃX9����w�-�!OԽС�kQt�};v���^x��������j�)��c��au?th�V��vԨ����Aʜ�1�r8	�TY�U�;�E7��4�m>����"r>400P��k����yͱh-��E����[n�E��4��wj����!ks�������d!{�v��u���y�n��)?�}!1]c]kN���,o�� 50���R�$�Fs@�U��Pk$KE����Ν�X�D?dkK�'�br���T�����U�߫��)���Lo�FcK�Wf��Jm��4�I���rO����"
3X�Q�Y(0��M�_򒗼��?Gg{���wz���[D�PK�hoꋳ�"w�.4n �ȧ5}���Ӽ���
|��J3��Yk�4��Lcj�TѾ�Z%�r�gH�.�S�����Q2��v�����>cډ���åٴ����\�����>=|W>�V��S*��3�J�m�/юh&	�[�s�z�)mf��.(����v�s�=���A?��R��a���JW���	���i�t�w�M���)��C�H������.k�?�H�X������,T�7>���4H`����t�C����>�ГHG΃ı�ݻwW[+t�tWiD�i�ԺM/�<�99Ob�**��5y��@���V����r����$��駏�q���`���-H��C��4�$��C��kd|����M�m�gny^'R[��x��+N83���g�b�`R��ⓔ>ǃ ;�k��gOHȲ�� �$D˸������
+Y�g΂҅X�r�e�1��c;bvܤ�,O�g���U�R��y��9��j�ӏ��Ȩ�@U�^��=:�OHSK�P�.��MSgF�0R:	��S�J	\*%�%	Id���.��Y��Lo�3��я|��8Z^�T,��~�t���y��#3���7����B�̉�~+�'��W]5TrSS����%$��-�e ��hqj*Z(��j�z�y��;��f����-����sw����j�J��M\�����T��h]�l��Ͽ�0-k��'��=9�i׮G,�1-=]��Ԩ��W�k	u��h������ԋ�
�b��"$j^�
)����g��������J�ٲь�I���J%�$H����.� ��WM2��R>x���M�]Ε����׻�Z��W}�� �S+�s#C����vD�V��S����b�ܐ���hzm���^Y]���|����b�]yt���p�5��ඥq����(�z��M�/~�F��N�������:IW� ��6����f
�v��x�x��S6�&�"�I���頓]'��.%PW�� 19�NuK��v�&褁����~��Ç����
�}nn��S}�It��1C�F�bK��dbf���5��iQ�#����Ky����Q3h�ݿo��������E�f6��{G�l�822�����cw�ygZ]�;��\0sf+�����{����\M�@T+��?e����>��jU�}j��i���ke_U�R(�	����A]B���C�qln���:[�Ǧ�k5چ�v��>�JV�q�5V��c����q	e9I���.�u�{�N0"�=8e�B�0��B|L�h�WA���z?X�����$�5������+��@@�& ��NdE�uuJ�n�?�(A�<H��F)s��eiB�Q��a;C�����<���R�vA����c#�d��Н��ͯ���fzK����>�)k�V��n�b�C��fO>j��A���e�\�&�%�Pr��]�����������t�1r6?�����AQ9jί��Go�q~��j�lێ�6Z�����a��v��׽~��gL7���'�8 J�1�� qFO�vcj�8B��q6�L��q �U�)����m|#M�������ᣇ��Λ kU��[��H_�\>n�	�¡Q�0�c���v0������Bf��#�3
�*O��]S�6��z��ku�3����?� ,K�O*5Z����gv��z�������w�#4����C�x��PLM�� K�rT$$3P#&�4bS��0�Q���\��l,��yup P�O����JZ� E�L��h�߽��;�[���7;�"yM�����w|�!�t�=�Y@,�/�G��V�֖�iW�Bf]�-�Vrgf������ҫ���ٳgj��7����L%S�J��rˇ�[s�>z�6�U�������=eݼॗ��X8>3���`���g$�2�*U�O9��A�i��>#���Z�*K��q�k=���$�Q\���B2h��s��"za�(R�jr!��>Y(J
�$���k�.Q!�̈1�������)7�0v�����-"��}DM��(iǵ�$�./h�Սa��.J�l�0hH-a�p#C����^��������l��x�=RAg"��I`�l����`'��IT%7M�txa@�{z2�ɺ�p*D�g�7{��z��X(����yt��o��3���j9�S��G��߿���7m��U���4/B�tج���в#;O���-��8E�(υ!|փØ:��z�7*����l�UK��W}�o������|�����_{�-[H�~�_x�[��k#LH�=>���M�����l��ْ->R�J�X��-d{4Vj)�ِ\Iʙ.�C|�)e���
��}�AiG��5��r��#>��sc���y�5�.%�d�6l� ���o�G/�c�B�G+�Hut%fۘ�l�u�M��B�u�!%��IL4Q�PA/�#�(�� k�)�J%סb�@QO�D�tвWؔ�ՙ��LZyg��ܔ��%�{R�7YZ ��7�q�vlq�..�ȧ-��y6�ONN&~��a3۾}�Ν;�K���v���D6@T�������� ���΅go�����¡�CP@"J��Xb�k�c��kn�MnK�F4�?�kGE��A�~�C;��{�u�5���;�ZsoPD�������<�٬=�,�7����]U/DP��X�MT�ۊn"B-�N��233�β�k�nݵ�^a" #���G�`��x��#�%g��n$��$����v�N �A�*B�Ed�@��@��$7��j9�K��
����,~������v:����#�=F�VJ�.>��!�2-0B")�rt@�J�<�%�&Ms�Js�z�D�3_e��b&yUz��3��[��̟Y������D��`�	�lD����u�8�u�2^�qʵ~7f�/�3��?a,��I&�WM��p/$�k9���	����9\�@6���˗�0�lcv�&4�4��H�$����(����t z�⢟�F��Y*�3�
�HiLOK��+�LZ������,9d!�>��� ��V�U)xeŢ��%ఝd�UV8w�T\��)���0҈̟Dz� ��=v�5k�By�lqi�$���&�6Y������&c�$\X�h7���u�ݥ�mٍ��	N���w�HT�DxT橓\+��4/1z������*p8Y�N�N����!T,'�|���"�PX��h y=|&�R�-Uz]�����҃���=o_�F� ���Yޗ��Z�(\�Q��%����SOIz�\vgBI�x�f��� �߷o�Y�h�� t ����~V?e^T�ӮX@����۴lIJcǴ
n!���Z�{�=��90F�����J5�V�#�t��.{衇�.�\ј����m���ݫ��|��l����3����U��;�����׾ů:3�M+�<`���1o엚�O��1R.I���=��M�\�O��3/�ɕ��=�s�������m	�zB�
O�"['��Y�G
���Q=T^zv�&���.�ŋ�J׏�� C��+b�!ÉP%z�Y�'�I!7C�>eJwG'M�SA�|��9&�:Og��n�|�W�����b*����UI��'?����nݪ�ԢWL�֖d�_��{���_^}�K�;�6�^���|�s�6=t�QG)x�Ԓ�n�����0�T�+N�4�G�	O\��9��֧��;˥�2��KnZ��J�3��f�ͣJ���x�Y9σ"JG3{屪+� �膙%ʦ�����'��e�˖Mu:�i%�e�I�|������+n��'�xכ�Bv�������o�J�)'g�K/}Ý�=p��_>>2�Fd��ZC'��%�L&���[�wO�:��^���=� �����I�U'��d�ر�!6�u�I��&�y\E�*��(�?�`iqj�z�U��m/�?�|�^.2&�W�
U�ݽ����؈�Y�Gqu����4&���A7��j��Pͩ��-5u%�9}�
3�}�������-��ӭ���Ꝡ���rL��vtF���n��&�d���2�0#[U��h��R��t�J����8K\�$CO�l`��\��a�C&�� �x؃1���oh'��Ʀ�t��]U!cN�ό��� �GL3���#j�-�l����Π�$�͕�>]��×����ѧ~��Gx����j�֬���]v�KO>��S�ۿu���߿�ч��l{���qA��)E�m�M[P-64H?�-�5�)3�v���ٖ�v����Qn*df�ƫS���֝jܞٵ����"��;d�:�k@IM>���Z����F)M�����E�跚�F[�S#	G,�����:B�Y�-��A���Ő��a��V@�ߢ�}��K]�z��{���?�����-[!8
t�9B��g��z�EÛ�_���iY�(�g�w���ԧ����pGFF<��;n϶���H���$������~D�ȲႶ9�!U�`�L���bih�����a����8�4:��H�!;a��d����g�����^�+y��ofA�nY�L�-"4|k��YHiS�r��]�TZ�:}���<I'�gt���Fe�EN�ew�-�FV)�]9�����5�u�ߒ�֬����؂��w�[�ة/>����/:���%'�6:::6 ��Һ�u�f���w_q����NN;B=c !GCx
,�q���V)�Nu�\��ёES;��ܹ�h�g�z����#GG�d��C ,��,��b�A;��Ȉ0���4��r���8�J�4:��ۅ~�4��>�k���K�<&��G�=8p��2۪�V@�V�Tܡ�!�l��E�ߴ#ep)+�_�j�-�$�ށv[�U���S��ó�`V�I��i_v��/�,p�+]xH�Z��j�T��k7p~�e�C��G�Q��M4{�+t�$$͝�j����R�n\E�8�x'%�v�E#�S^�.��;���o���ni6��S(z�l�&+�:<�jߍ?��W��<0ڮ�>��6%�3�?	=�or�h#��ru���M7��~p�ƝT�+0�R�����7������x衇:e��:�M?���P���-`�o_����8;���O�'�p�'�uE\ʵ��9`��t��H	c��פ׺�����BD)��0c�I�Z�l��H�,�nJQ���"����J��^U���T;t�f�Z@i��K����D�1ΐ��3��)>���!華�B��\�Yy!v
���vs�`��cDx�,�t���ԲLME�p��t� QyW�8w�+R�^ Q�;T�!�b�	_V�M�`��u�Rߞ��r[N\�\�*�j�>��|����0u�s6b�a�,��-��FYh��*Q|Z�69�*�'\R�z�8��F�=�������f�a�؜��X6�C�ѴV�8N�M�ڎ������'F���40}�t��4@���^�t_ՊC�1�<_��ϛ�eEJ��G�md%��ڲ.5`<P��)��L�gr�������p����?�w����8�<��X�Q��(:��3I�_q���~�k_��/~��SOݶmۢ�ChG<�3h�������C��;rGHaY��#�o��|i�=B�^��\D�&�OI������^�t���+�<m-�k�/��/��Y�%
�s���'�p饗"�N�G�5t#cv�U�Vw�q7�|�m��v�+�������u7�t����m[~�ڦm�J���w��,@f0�8Ɵ*9��w�UA�(L�~��n(�X����*����K�9^� �f!g�e�r�U�f���5A�])�q�6�X�}�((������i�ϒT��<�|�#u ����ݱe��]�Xq<��Q���t���!�ffp5�������>�e�l��G��а�?�E�L%�}�e�}C{����}j}�o�}�Uj ��Ց��m�K�H�*�s`s2hLfgg7nܸ��n߾]�ӣ�:�T.�u�Y�Z�;�G�j]�b�	'�p���>���S�����Sra��ɫ��e�@���J�1�i��Dc�o��|:����M�!�u�bpd�Y8:_j��ג1a�&�{��0zld	�Ť���#J��T a������$3�Nw��u���te�z�]��}����g����g�ӧ�y�;߹i��/�����Ɏ.���sqDeN)e#H��F�e���̲��G���~�N��$'�8�8�J���En�q ظs�. gh�i�j�&�����Ñ�J�(����AЕ�(�S)&��O��^!Iz��g���cn�$��ɬ�6�5�A���v;�
�C�-ϖD>=��r~0Q��`2��x�@��9+"�_A�#� ח�Bx�)�\|��G��ο���N�aÆ,��k���t��P�MD�9�}����a����W�!7;9	G�S������� ��Zݻwo�G�����n��ɦ��P�X����ѝw޹k�#�8�ŧK� �&��,'��|����*>Zb,� F�Ӓ{F3n�H�W�Iz���~c�,\���g��Ah|�qPQ��E{�͜�O�D�d�[A7�3Qbv	(�҇���8O�2b�$��n~i�ΛBEN���n��g���5��62����{vl�Q�Ak��m`-wTg�	O�AŒ�S��t;�:�d�%*�r���(M�W޽{��T�󔸣"������i�S�z�	��wI���������t��8"{����AQ+}z�g��}.O�g!�˦}c�!Eha=G�/���4ԌD�+@�>���_G=m���L��f�]�!��6SH��t<Q3��������(��_1�v�-���ɿ#�Ͷc�����K���E�����(�&��$��-cJ�����k����^��W�/���yQ��,-�m./�#�,�������m��;��e�0,Y�u�6�N�t�#�ȿ|������u�EB���\�@��_����Y?_�8-8r�lK32�޻�>�寠����7���y'-�^��W�P`i�bTtڔO<��Z-������o?L됬Bz�o}�[���f���%�{�O�����MƁ�F�/iE�'{qA��x��z�C#��Y�k��O��	��^����� �/�㭭X����}׿�����_^x�'�t�ٯ8��?�iՊUQ�5�b^p��\��$!���u��3��Ht�hOIH�s�)��D?�n���6h^N&k@��<s-��y!N��[��*+V�h�>���pT�R�8N��k_�Z']�j�-�0-�v\��/y��o��ֳ���f�{��������7-˳�=����N�\beGJO���%#��<]߫��OZKY�܅��v����EKM�Kb=(�]Vu�Nh���MU=�s��Eh"2՞^��T�㈲=[��L����z�n�Ru�V���⪕G�޼qff��VG�G'�m���y�+�� �p
������n�0�����0U�[��uȄ/  Ҧ�g�oxzϞ}�!W���d}��n��FA��t��}{Mo`ph����=8Q-�:Yl�zH&c�]N@*R F��f�y���CG�lߴ�����#?rȾ	�>���£0IJ��p�7�]0w�9�ĴQ���Y_ļ���B�w�T��(d��
]A3�͛7��g�@V������ɟ�������&7�Ԃ�⥋^�֋뵙�]u�G,���^���=|��w�u׆Gu���-Z�266�6�FX9�Y��E68��Xc��~e�Bq��� ��������}���O�W�D��?R,����4�XI��K0�n΢�PQm�J������@,C�>�h�ܲ���v<ujj��mٲe����9S^�Ƚ50D6��5�[v�x��ǧj5�V7!c�D .d{����a�Y�S5Ϭ�#;J_aհ@HT�i�p����P21g}{�,W�t���z�L��m�eK]�m'�ۜ������t�H~&݋~'fb�dP�����R���iE��"o5o�+җ���K�5ҋi�:VS�U�N�F�Ѷ��ZPZ�c<8�F�:$��2_��FA��BA\�"&�S�L�P��V,I��p��C޷g;}�&�~V]���6<��Hdm�.Uj�ڈ]m6�]�: Z8\��1��������2�f�Mہ��i K��ݳ5[G�w�ٖ5���1p/[~���e�V`�t���ďY~tzΙz{����lU���,ߧ7*�ұi����j�O
"JV�XVy�j*�J�-���@��� �C�?P��&�����;)�$-���b�&
ȹn�J$�K��H���p�}cd-[@�WI�u-��A�=9�4
�$��3+=���ϐT���H��JGj=,C��IH'{<3�(Lڭn��"����ݻ���FzI7��1�5�m����A��F�����Z-Ԥ:^L6z_hw5��!ǀ���T�cm�zUG
�Ob�h���6�[�F��P0��ۘ��_7�J�b��BO�U�M�Y�����t��l4��#� q�^�A:��y�x:W{0��s���3^J�{�@rE�-�(NuT�������������J �G��W���?};)�F�U*����ͯ�]�h@-�Š	F���މ=4��`���r�a���x�t�IS�]#Ʒ^�ڋ����Ԁ�Dq���]��2RJa��ê��E��}���|�v�r���gh���"0�41P_b��J�<�%��o��^T���on0(�l0�V޵��9N�d��q^J�ّ?�	�@=�y� J�B���^p�b��\���{�=�c_���>��{z��?���EmD	����������ĆG�>�貭�ؒ��i�K/���?5c�hǴ�;�r���4��bL��mA[�p��_�ܿ��Ffx��t8f��_��_}��ߦ�2Z�?�^��|�J�bY��TK�ل���&�z��k=��*����ɧ_�d	�Bv,m{(�P�{�E��?���>�1��--��k��������俘�G��^�_���Gԫ��w&�s�G��3 ��($��m�I���owʟd�J�Z..�#
�>�/Nb*�]q�z r}�.a�A	{qy�����D��a�_�^��ŨeP���h�s��=�y�{ߛr�^���?���}�:3����$P.+�O/���l��h�;O�N���_�|	d�"�������d���G~@2@�HVD�Z/~�'Nmٲ5B�:F�z�c�a�Tq����<��aRʸX\2]dٝv�i�V��n��Ж�27ct�4@f��Cb -��T���ȡ���n���\��j�~u��3?2��Y�x�~M�K � �w��C@�7��l Rbh癙��{�I�cD����n���{�}�{��m7��������_r�%�(����#�lݺu��������ڸq�7�@v�K��e�=�jՓO>��;h���W�X��n1��A4��X�Im���o���:�Yk�H?�9�d�� �`�u����X��*�L�	��TƁQa��16<B`��B��Q�B?@/��8�m�zPGȖFXd�sL��#����k`"zt�: (���5��=��d�<z�æ%��GOu�U��P67��1�����"�@�h���u�����_�z<]J�&�7����F�[J���o(�^�/Qa2J9)�)�)�W3��)���d)�X���Y2��8Q������>�I��AҘ���0��CW�vldpdd�ݩ8p��Z`?E3�ӆl���W�t�	�^.�6v&#��N&�����Oe�pAu ��&�k�'4J����
D�����
���dB#�-T[�����V��\&ɉ�0��t�mVY�J���ᕜo�kj@�1<HQ���[/_�|߾}Ʋ7xi�F�[�W-bn�"*-��n�[>j =�@�8�M�}��Y��r9fZ���W��m:�^
�"��@�e�bh׬_ʑq}A^-қ�LR=�Lu���/���K!��r�{���d�H_����t��0�Me�T6�8/W�L{���M�	��%�f���r#;��W����p��'(��}�IR2�f����K�.��	I�Hq� <�A[?�Jj����42\_ΥS~���oϯ�a$�����������3O?˶l�x:-�K˺��x�_l߾}��j��ȩ`� g�y}�'<9��w�y��ǒ0lAy�U 6RǇ*��~����qf��4�M|?o��fZ��_~�?����{R��.~��t͍�j�|�����'�|���~�&��r��i��˫}���S-e����^>V�0��_��<�$��[�cR�0Lc���ɖ��7���7��f$��bg�����}�+���'���wh咮����󗗗���eh3ݹsϟ��_��i�Y�fM�D��W�'�x�nA�p_%=�i��p����q��z���H9�`�� 8\�7D�wם_��W,�|`ׁf�_q��?��O�����u�3K�z]���͇���j������j�FqhX��=SS
�1=�j[�i�(��[Ma�p��Q"v��(�>�����?}��Ya�WP �b���gUh7�d�ݔV�hF�A�
�d�.l�������K�$�,��#�
�F�c�R�#�i�(����Y��Տ�3�8�%8�5�u�I#&_��27tx�v�p�Ws8��d<p�'37I��_�H��kͯ'ԕ���|��p���/@��j�ET��p!7OLҏ]1uj������Ԁ�T�)�/�c�HD��j֝�"�=Ï�~�.L[z��QZd�Y6����d�������F�y0�,V2쯅J��̨31Sw]�-��r�4TQo߾�$�~���z��&ZH�˥F���v�LtM		�{�Ĉ>��6ei�\_�P�m�I[�2M��D"g�	
5��.A��bf��ӭ��#�lf�C�$�T��f�{!�Hޤ�9�k;.
3 dͶF_6ͽ[g�V[���j�T��⅋��ػ�[*�����Qqa��gG�e�㖖���)����h���O�vǰ�~�iK7�vw�W�nxZӦL}�o1��y1��*^��Jd�I�k8�m�d�%�����|+� Ѥs@1ْ��
�Kl*�g����q`�� l��F�=PEM�}��z�n�V̦$v�H�>k��1�ߗ�XAv箩Y�_���dI����L�,Y�m?(m��{6j����W)�ggM'�
d�v>U��F/${���\�J�8
J����"_=���
�� @B�����r�B�����C��#%��&�&I>,�a#?L8t�����\M�ͽQ�9�k�~}��/���%$���xdV��p*�Z�%J��;�K:��aۏ,˦�	B2���g#�ّ�-6�#Q��<�{��.��4�M(j�\T���E#�$����P�g6���y�\Ch0kM�Ͻ��]r�,Ӷ�����4���=K+�̗��&��B?��&yK���0*��`>a�N�N��N��a��ܱ�9zN:3VT�f�I�B�
%â�1"A?�L1m'pL�@�8/�2��=��U�C^��׃.bR������E�_J�]�|�:)fBe~j%L�|h��m��z�P�3g���F7͑K�<�Wf�7�)H���Lr�,�U�D[i/��Â���_@�f� �PAs��XaWS\���)���z6P0��b}�E��\r���S���_���42t����E�� d�2�����T\�|�h�T��I�iA�1@3�X��ڞQpU��F�.
!��l�z�etZ��R�]1�~��^�ޠ���I��i��q�@ȉ1!V�/���_2����C�)�X��c>x��g��4�{�y�]s͏��TО�o�s�'NգW����;TJA�hʗ���׿�MtGK�0R�����o���ǿ�����r#p/�Eщg8�=�淿�0�W_p>��	@{����+���+>��+^t��������|��k�w���[���0x����o����o��rZ�a:���
E�s�>��.J����oǒx��Y�5m���&}���ʳ[� �\J��'af��'c�[1��TW͈T[�>��ܺ}�m��lb_}�Ȳ�v�-���l7�� ޓ`�O�m�7]v�m�����~���ג.i�fW����V���cא8����h����{���_?���
��\��x������������C��i�U�k����썷�V�V�$3��[�8��ӯ��5����@������K�n�^B6!������_�y	c��M���L,ӂ��H�� "z9
�'�.NF�?j]�V�/�v��q��G��B�J(��`W�:�!q_�4S��. ����R�.Y,t���4nԑ���f���4~�h�RB�'DL�u�)�s H$)� JF�G�y�b���Z�pVL"��p�l��]���3xWj.��:� �2;��v���
����z�wt�hrgff��M\�D��$��{�}|<	R>���^�<G�M�#'�f������G�}��%ɥ���?����[,�6��c�=�,�ӭ�;w��3�D�	���\}D������"����ŋ�ȿ袋Z�����;�����FQ�s��Gr�!{'j?���kMĨ�>�8��Ft~��82���z�iy���{8��LP���r�w����ؖ��H�u0�gS�n��+�k�A�?�Uw�7�_�>Vӳ�:��^�랢��,:�#�(��={��nm�������?߰�;=[���⥧/Y������w_��/_�ҷ��.�s�c��s��-��73C�+�`2bd�c~�U� i��f �m���<94>���]5ݵkyѰo���!�b�Y(�4�v{�ڇ�2Ք�[�ޭ&���^Ac.��k�j�h���FÎޛ8%�W�;�c�9�88p�g*�=nش��_�r�Hn$�+�I��i� �[%�w��ͻHo��R� �{e����Mɐ(}f9MC��B�"Y�g��Kw�@�@j�d��[�r��^�ւD�H��frru���O���]����#�n[Ȋ���@�bV��r/7�(�p&���Zj��K*[S�X��UpQ͘��~�2����ʅ=�L(]�aE��?�~d��<F��BcJ��955��Nz�[�:<���O>q ���rQ�J��A@�[�A��X)�Tvyd�=�^���p-� �'��GKE4,�$!/���J�;4��#3���g�%C_ٴm?��8VV�ZF�IZ�d�-R>�����T7���M�Yo.^���Iܔ<�_DU�ZY4�$O��+�}�ZEԯ�l���4�ǆ���I�)��4�
ސ��7NM���
���x��*��|���������6�T�������Qu���p�v�邎���1R���m��A�t`_gzzzj?)���h܍���(����W�^=�d)Y�R����?�����)g��.:���֧����LۤU?�PV�IK�;��)U��<\�\��U�%n�����C�3�����-�$Kivf��K.��}�߸�7��[}�*mR�-/~�~�_lڴ��c���~
����ln��g>�m{v�W@+h|l<�&�D���ؤYZA��/�
��n����G�����/�ڧ>����/q�I'���什��2-ZE�)=�������O��+h�׮]���̱��X7���y6�����yϸb�L���q·}�y����D����Ͽ��y�#�L�~	|�`<厰�t����4X�j���\�dr�y睤��ޖ���k�=��i[Y�r�����vȲ�l�K������PЕ(��4�����*���8P�\D��O~������D�t-�t��c�9��,5�4}
����������[}�#���*~�R�P�|��;8�I�
V�i
�u�h\�g	3�2�8�@��_K��A|�s�T�ܒ��.RC	�;�<����?�>����a\*�$W�y X:�$H,�Y�yA9�hZ-�1b��T������c����0�l�����\$���8�� �l���I8��h�E'+�-C��>cw+6��,�8$ ��*�M^+��W�o��oA42?By9��\���w�#� �A5!�0K�
�C��A����,ĘL��p��̡= Ml��4��'�8X���ό��r�x�����l�c��Fx7�DK;Q:UoM�:m��j$�	4 !�P#&凞�N���(2��Z.����N-O���g�Z$�����L�x�	g[��c�!e��0��ߦ'wLF���l�igqK�m���J"/���p&����N	ʥb�+qH�:1lY��AU�z� u1HӘ^Q��13C�3�6?������ãŁ���;7n9��CǇG�N��j��e�1�vcrV�h�yi�,�#���153�WǗ������Su�<��R�.Y��m�k���lm�����G2q�9x^�P.y-�fO� ����4o������Jɤ-�^ylr�0��(Bc�AYF7)��i�Z*&����"l1B/T�`vE!p/vH�D�F"`��ݵ{��ꐕ?��f�ā����0y�a�Ж�{�^.����C �3@"^�X��Yի*̃�꼂%e�C���毣��rN޲L�Zl��!��0j%�#z��H�M���M�N�̌�����l�	���
3�W8]�I���ɩP��w/�ʦ+��4���<����� ��P1�x����dȢl,J]��(�Kp�d:l���D�o�u�rA�ǹ4D�9��s�����ƩT�I�<|$j���~�= ޳"�if� 4]�z� ����� 
f󄅂�$�Dq
��� 
���l��\�64�_��Z�u`멖GkzB��ز�n�����)rvbU1�r��%0R�P�V�wg��Rz�6�8[%w0��Mt�Ɩ 5>��C���F._���'��B�8�x.���q��F��+~��U(���o߾���qM���������RE���5�v0d}�N2�KN	4��<��ɞ��K��T&��٩c1��(к	8S��f�m#71كH�$�I��u[����F�l7u�%�k7���6��5dt��`Y�3�u-�Y��=�%S���c�����h֚-g�ZhԢ�`��LG>�C��9�Z��.A�*��� 8�tkj�1��z@��źm��S��H��h�a�K�,���(���Jh&�J� {�QUCſ6�'���O��ش�;������?�;��W���:�O��>e���C�oݹ�5Ǚ��Z�%�΀����3��eː4�N����z�W�(A������{�>�>���l�)�R��ǳ�
������?�跿��w}❍8 �6ٍOo:��5�Q�-�="z��8D�:Z�1"����lJ���)N�Q��s:�Y���k	r�}�ju^�A�ׂ��TW*' e���TǴ�r���/�ڧQ�T����(N�m۷���@bT�{�9W|�S7����_t��:�SS>�л�������_�{�t��Ow��t�G�=>;[_�b<�
����)�7\v�/n��ݷ�q�ůglZ��7t��^y�Y.*~P�iV����B[�f�Z)�uŊZ؅T=��Co����7/?��XM8-�l4��FL�����<��.a�qzƁ 04��| E{��T  ��IDAT����=�2m�u�:��(��l@0���g�%|B���h�o}!U"��*�?��&'KA��D�Ĝ��7�e)J���Y�H��
�2@�iE����]b�Im7mF��p�=+�RI��A���,��bTeDn�%��W�'��%��LS�����^/k���m9�����&6�(���I�\&�Mz�Ej/�Y�Q&�>�����߿ɒ%da�/�{i�N{ɉ�{.�GT�Ǩ/�����[-��?���7n�5�o޼��Fp�,N"�k3�薙��~��ׯ�{�j�9�c����k�?Ъ�y�:4@�=�q�}�����݈"
�7+�j��@>�0��O�c ��"�� `J��A��4u�&�o���`�^����l��~=�d��f�E�s��i�,<dՂ�F@�6�p�F�|�����=�j���N"�ߺq�-[�?�����vl�[����!��x�8��mW_G���^�2dQ�����g�.2-�zի*�ʮO�8���]�e5��MM�������$��\,����LB#0YC΁V��А�#'�Z�p��ʕn��Az�*-�s�=�t�����n1�<�Q��4F),�P���^���^�c��^�~�S�ӽ�����eH
u�dpp�q
/A#O�̷�<z�/������2��3?��sX;$5�<�SF�0��!3�\rK_��Tν;4[�l�yG�5e|XmB7
R�*�"P����X5@�F7���0IQ�I�Y��M0~�����3hm����T���Y�tJ�'�J3S7�������̰DF��,��c���3e��0L�X�L�x�b��[o���GUR�R�9a5���Fn��"�^�;E���rҊ+q���	Ւ�+��q!sl���Sv�2�
ش�=u��h|���F�H�l,Z��u�{�ۣwٽ� ��D.$_���:4G!�w#�E�.� ������� �QH�]��c�SK��;�3O��r�Q���'hU�<82R���$Q��7���*$6��Ţ�0�wH�H�����u���ܻ�F�vL!&Rt��J/��w�ћ��I{�X��7������-�iҸ/��i�e�����){GR�O�����D0~� ٶ�wh���K猍Qsx����ҥt�G֭۴i��(�ќ�J7�˅.�m۶П=���$]�r�ľ�4,3�S�ж`B��f���V������;��� � I��t�7Rt�\q֋\����~����w<l���*I�a���Yg�%��8�����;�"�c��r�ܫ"�����`-	?���q��I�v�ؑCG�ґ�t�kZ���I7<��-K��;�d2�,��O?�R��]�6Q��|�SO=ult���~7�C���Ї>Dw�A���Q���p�g����˭�LT�5�v�~Vvq�����>W�:��(����N0�02Zd�]M�gS8�����~��7�x�+_����Q�{��bq�֭$���� ��@�}��Y�k�����>���J����Te�{�f�����|-Q}O=��޽3����ҙ��)nM��,2�I���R^K'`	+j�H�Y�^[Z����8^�� �I��09ĥ��b����ƥ�X���
*�L�I�@�$F l\�FԄ�$ʛ��'���<�e1�柣����m$���,��������6�+�/]�Q�4S
6�D砟�k��$wª��:�Y�0�]&Ъ=oV(�\$&��v��g�N�zP`�\U��9|�_YJ��F4�q�_)���2�x#�&�2�.5�TM8�%�X���HWSC����H	)h�����D�%)����eA2dF���h�-;w�G����K���l�UO�ʚN�&�b�ځ��ӱd�H R�W@h0�n9~��4��B����]{-[۳g���8�%J��I�f ə���Lm�ݻ��I�T�4rJl�"������jj��^�$�A^�S����|B<`䊻nf����*l�$�	:���4= ���ax�0貿�vș �'`���:a�}p�v�3�ܨ���d��ff�������� Yh�IO�gF�s�Z
$3��ZXi��ll6�AC��G8�5�d)��M{v-]�4���ұ�ə���5{�Q��A�/z�=�dI�w�Uڙn1:B��N���>"q��L�>���4����3��3fj��DaL�1�:����HgZ����`� Yڜ�r<׮V�3��ǝN�l"&���)��?�2�����hd|A0<Bs}Ȫ�P��SS3###d�-#���U����7Ro, �(D)<���*R���5�/�M�28��chJnI���O���v;�{
�/b��@#CV�	T�#}/p���x5b`!%�y$r�S{wa�x�b:��r�!-��Ì�0E!V�ǰ�4��cM��lx��CY�*w���뜩&Þ�	X��oײ`�8@�X�ɚAr�b�8��6�~8:G�4���.F��g�EpP �>=}�%Х�@�08�ph �=m��K�� /C	��m����~؃Ň�F�c�w�Q�9nš�D^�Z��:�����#�ӈ��3
+KF��A�x&j��h����%YR,�e�Ԃ:P��2o�i�Ч�n�g:��TO�Yň����"9S��7<⎂���;ˡiiHhx�2��N�zU�<Ǣ��4[����Ck�69��`9CK���3�.l���m��(�V�G�Pa$��[�L�Uȱ�L��ztl@t�p�Lv�8��+vɤ'����QU�Uc8xl�Wn��I�Z�C��Q��=��V
���x�ZkEq
&�=����Җ�Z^]��Cmٲ�Vk�J@O�mSz"</}D�2�S���iXt��1�	JM׫B��:��n��eUFi�}ϮZ����Xs ]�4+�Ъ�C��"1$ b�C��1�F
U�ȁ�d`�UA~���E'�t.�Ws}��A
@��55ӈ�{�S[I��-=��#'��/�n+*�2?�����!iL򸠱t�A}Ï��7�p�y睇�UZ#��l��Er(��Ƨ�����Е跓'G ,\����袂]t�N�:n��,������W,\�@��[s���o]��� U]Naơ.Qx �$��0���ﭒ���y������3|�y�V�U��E�2�44/�V��y�?�P�q]10o��b����|��g/��(u(Y�ۿ�����._�򗝺��I��Un���<x�9�t��/>�\xj���(�{mݱs��Cm/�6i�vܡi4Lo�8pΩ�?�_��J#��U��`�염�m۶eA�b�pU'��.�B`ŕ,r�;x�4�?�B����m\J�A�8����xZ/�Z�<3����{���#SDz��	a��I:R?�5r��%(O�y�i7ɑ�)FO�����_�W�n�~e��(H���&?,Ôx	[�qe�Rϭ
_��Dq��W��h�bN-��^��`�srL'ŝH_�����r>�����?�q[V��J�~A�3]AA������=,T�1�Z7ʸk��VT��G��n��X3� �0l�l��tG��*#��o�K��Z
�L.FE|�,�Q�Z-�?=��}k׮����v}�K{���g �M4�D˫�'�� ]�^��Z��� W���_�� eӥs��U�-����?0F�j�DV/itF�VȮ*z��1{�����1�� �-�`�󔞙.Nw����8�E���}��f��裏^}��dٜp�I.l'�]��޼��tɒ%˖-K��]w���vN;�ҢQ�{]�{���\��1z��6n�x���7���}Lax%zZ�ے<2Q	�����E̾Tܾ}�c����;����$P�Z]��� �a��lu^�*�X�����o��	�w�r@�ô�J=�G�)gv���M�#έ��v�Ak����W9�t�a�f8�����hp�'ɋ{s�B�kFxSӜ_�/�Z�m�>�UY6��5��{ShR5�H{�l�p��š�Orf��1ʥa���#���F�q㊡��¬�b���	4K�����N�Q#�q*���[6�����q��'	*]��Y��3N�o�ʈ�W���B��p,R��n�%O�P�Q�ߥ\��Y�2�4}�:f�|K�$W���L��իW��}�;��tڕ����䄖9]L6dx�	'����d�:r�z��z��;���J3D@ZI(��R��%נ���3�fg�%�=��n�$M��.�\z�h�Ӷ�M��9$>���a��ܱc�g���4n����iu�QO��4��H�[�8��EO^]~��lԤ��g��"J�����$�0{���ա[��8�dŲ}���Ù��J�B5K,;��S(�8l�����0r�(�\GvO���2�p�	�Zh���C�+B8�M��,�������"���.|9-����ܲ��?24Lb�M�6�~��7�t��]���po�
�Y��kc���L�1Y8^�Q=��C?���
��`Atl�a��-{�����M{D�ʘG�gа蝦��X$W�9yV��F�L�/C�b����H���(����H��JEL��SOw�q:C�hC'��GW���N�
ms���W�}�UW�GǑ�o}[�����]s>W����/�
a[��!]mݺu˗/giGA:gFTjh�k�J �ZV4�YT��+��Ra�/>\���G�|��i 0����I���Q�>�����& P�y9t�w)�ڱ�u�j9�2J�u��91F~���7?�C�J�X�u�
[���w����(�֬Ys���T�����/|߻�G;���I�Z�;�[��}�k�Z�t�?�A��궡F��EUΫ^��ۯ���ģ���~�;�9묳�+�O�uv�f�@[��oo3�;c��(����,F����<GOi\�ͽC=�<�
�R���@�G�I���b��)bMI#?�m�u=�1,���e4?��Q�Ɂ�ɫ����31��]�W�E���a,.��K�2��\`���!?��T�*�,��4��8���
�߀��ٳb�'AY5�y||�$�j��kG����R��)����&�̔�f��A�
(�,P��v����PK8��=!�}/ڜv�3Sq,'�b�v:��)~�FͶF�%a�v��"�ÊeR)��hf{�RGLZ���E��4�d��j�g+���͠�8�i���v+`���Զl�z� ��A�Q6�˚��穕"0,�����-e�:zWh Fӛ䃆�O�$�V$�T%��ӄ|0B��(DD�'��+�--R�^�v���΃�s z2�5_�ɢѡ8;�L�Ƀ�u5^�dpd@��}+��ZT���kz�@sz������@�ţ�nk��A�Z��JJ�rʳi�؎ͺ�Mk�!CհݤUL�g)�*#�U�*�a�v���ڴd$w��lL���]�U¦OoM���Xӵ��ڋ/V�� 
��%v���c3E��b�h4�Di"]4*4�d)�3�?j�h�nsZ۷͉�ɝiJ�T[5[`)J�F7�&g�,**���P:�؟1�
�MoA�m������p���W�J�a��i�_�r�A�n���!u���$lY���O��,@���r��c�W�*l5��p�"Y_b���1������.�N""=�9X����*�ش�8�� ���2Rk��ROa�9���"t��*�\�蹃�U2;�N�Z�����Y�Z�Ъ@���J��u%�L��%�E�� F������ZZ������'wPgk3�<=���32*�e��lhOrt�G�Th��"/L��M{B�h�I�˱؄���Z��{Ƶ��g,������YQofq`%�ޫq!�Z���pMr���N��ȳ�%���2�����,�z�D�f��2M��ǥ�"%�819�b�DJ0�T�3�y�C%�HU�&9�~�ؐc�A�Aˊ��02H�iL��D��9��>5���/KG�ISQ����&O�,:]�s�����F�Y�������f��Pa�d��e��4�ZZ������j݆�s˺��,i�TG���0��s��l���<��ly�6H,1�;�&�O"E!:Ҽ�� U���28jy��R�T��
=T��xb˖m�w쪅m�QŴ��q�A�۩T,r0h2���rM�y2M�DMmKaL�MA�ui�:a��TzX�LR���S�<��_�A�Tó?kj�{��q��c��}����T��Θ��*�����W�C2h x�OЅD�3:ȯ&�2���>��;o�K#���QDۉ����cpZ��AMȅ&ͣ�Q�sc-l�<�
�Y�����_���{��^{u�i$�����K_��[�������!k\@�����X�uG���C�1�r��%/.����'�ɕ�(��!�$5�^���
Z0���U�qH�l8����7^�����t:@æ[|0%������b��M�[��|�o��V��6���l��,ڴg
���Е���O��&I�v��)|�Y�7�x��ǯ~�3���\�F=���B��:]�Pd>C��)$�\2EZ@��4��nе�9K5����{~��k����ʤE'�S.�6M�S�s%1RQA��ı��A�D-F�a��z�"g����ƿ�#1�\ �[Κ'�>���4���C�N".qэ(�l���!1�S�]�o���B�S�q�nru��^$�ߜ#z��|ބ��ϑ�C��P�WfJ�&6��Z���@,K���l��]4�j����9#u��W���=��������#����	�����}�|F�W��\F����4-�kƜ��z��NNRMgd��
�ٸG+���@�LD�D́L�J2b���eKQ	�F�Z�����8�����V�����@d���󪉌�s��w��G��_�qö�F������?���'K���ç�z��N>����_���'���|�����y��l���N1��_x�)��t��4�<�����)�u�g<���k��fiu�Ω,T�eh���y:�F��z]a���܊�M����P�ٰ�uZ샃�Z��&���r�� �-z&h~(�B%��ef2DmC�@��i��Q(а���={�����l��J��s�����hAI����	ʟd�x{�r_+y������IE��B�N��C���:r�nA�Pɪ����Еb?�9;a�qbo*ν5���<���uxY�dJ�^��h��C���QT��>S$�mz�yu���V�0t����d@�H��\u-5Y�u�`=�tw�4�x��Cʅ�$���Ց�M{���?���iU*��=��ch	�F��'7�4���	g)����͙��%
r݅��L��h�"���;@�$_]��&�l0��h\o3^[�Nq��dh'�|�̻d�T��n�(����;:&�}�	�щ]`�g骃����I۴%LA��S��y�	�t���Ig��K����"���������v�������\OT��l
��p�r������ٜ�ř�&SV�RL|��j$FH�q."��#B`�I�`݋�ר��DE$>	#�a��j3AP�ꪫh�ܿ��C=����9{��]�v톍��뮭;���]���2�i/ϓ�=v�("��}t(�F���O�Z�j��՞���7l��;���G�\��L�DI@���Ӈ(�KF��d�a*r�$�#���K�XA/��r��a�������&�&WJUn��'v��uآ�t,�di\|��oy�[�-�i�y��f���t����7�yѥo�Te��G(�hH}h�����:Ѕ�H$bݺu4\kּH�R�Ji�hz/�N닶L�D������O<���.�G,��w?��Ooٲ��{챍'��+��{G�TU�F�[i-��m~�R�,��خ� �9����D�����ٓ���fL�)�-������ڪQ�C=
��44'�p�K����ꬳ�R8�GO��¹������R�s��8�ٶz�d$�Ѽ�e/�������˯��:��K/�T��csNV+-�m۶�X��^/��(�7o�Pҹ�|�D��p��=^�� ��]�{�Y�1�t9f��"l�����v�vu� �f��o����lM�T� �m� ��-��Kx�]���"(�r��KF�+�%
¶ѹ�zz����k��+(J��&��� ��x 	�e��'Y�ҿ��*yt�����q)!y�Y�=�1���3�}k}$/4���N�3U�
�^FYա�?M�j��e*���!{�$)�Ԅ��(8�A���-��u���������[��S�jz��� �Tʡ2h3�[�X��k�ֺ8�}Z0�ٹ�C�������nBUl�%>2+�TݢI�Ds�,����J�K0���P(������?3u��b��v���O�药�'����h%��SN9f�*��?���'6� ����/���h�Ҭ���U�1���(=�x�j�K�����%��e�t����m[��ؽ��CV�$��]o����/����n�.w���I������B�ozu���'}�_��OZ04�h�N�;�&?28r�%��ٶch�R�)5����N�8T�z{pj-L�"j��
�C��O������!d;Z���羂&��/}�c���wm�t�� p�;�G-;>�
(i=JA`�Kcę2�i����A\�e��vq�������>���۷�������Ⱥ�]�Y��,���Y�Z>P�H�hc���.�(v.۽}N�qd)�j1��3�*}޼��?sQ
X��H� I����DW�������0��s��?��B.�f}�䇮�p�BR� �7ͩ�iRz�uӋ�c��A34����l���罂2��W\��7*/l�,j=���sk���dWJ��$���t�T��I�����I�����1T�k�k4]�@�Ao=[k����d\mS�x�wь���\NB �q��ccc��X��!jF^�=1�,��Β�/_B�����\��հ;���
:��Ձ!T�a�7mq�< ��+XY62>t��q��nu�nd
	K�e�X:�0a}�bI�����n���C@�P�0����	#�G<�l���2�lYeh�:BJ�J2E�_�v���^c��0vk�*�&jF?��lV�ڱc�l�I#�4ݬZ)�j+N���J�Z�*���t��2Q����v7�Z�&�L��%d�e�ml޽�I�yri��e2�-��H�Ǚ�� a���������44L&1-ؤ�V��!'}z*53-���
��Pq~x��$]����.�F��e���w;q�j�G̻�H*��5G73�8@35�n�ػk�<ػ�E��
�]ꠔ4�rq$�[vm/z�0�ep��VS�):�ɕry	�3*Wj��-�n��ݮ���0*9�[,iX4�LW�Z.�}���,f�i1�c.f	�Y��_��Wn���է�PC��Д� J�aH�*C�uU�e��n)��@�w��m�]7Ap��Q��>s]e:m�����lZ�o~�e7�p�?����_���1%'4A������� ��,�D+��t���9)1H���P	�k�-,����b�5��k����5xwm�ڻI�ZH�H��q4���:�s���U�U�gf4��wW�zDs�N����������{���v����?vб����|�l֛�<�z@�����'�g
��΅��;�k�D;�~R#M.����vC�G*����*&�`br��2f-�l[)1�t9�V�������>��.WZSU�	�:�dA��M
6���V�=2
�`,�m!t7���:��/=����7�wwz~=�ۢGq-��9cfn�᝿�;������~��w}�W`ḵyS�tM���=6�[o}߷����C��/��sC�+NL�<��3��v���b��t٬��9�̌'��s[��z���B�͉�BdBǊF����3*J����� �zxL樟��F��)�Y/�Lq�r�}v7��@<�hs��2'�k^�:~-�+"��OUuM�%��*9g*���)�^N�$K	�S�İ��r0�Ed. �|�����3��6?s}�����H��D�l������(O
V$1�Bb��lԠ�r��k```߱c�a��k�,Y�D߹s����˦HP����, �C�v���3rۆ�c-"��V�|<F�����r���Pu"A5�`���(�L�BH�f%���N���I�0�w���ܴ� ��3,1�+�t��~�����񎎎N���^�l�1������8d���3��	}e�J�@�`�p73��sO�>=93���s�-�LMM����w�H�����zxx<}��c�����b��[o�u`pў={�y�x�+�z�ҥKG���w����s�W���[3EdY�uĪ�K{&��>�j���X(�����_�岵k�n{Ǖ��e2p5�6|;92r��!�^��;2hm�JSxsߋ�$i�l�$��[�F��X e�q|����qd��CCCFF���ݼq��͵���l߹��'��d��WT��q���_��J��f�>�*Q��I���#�RB/Ɋ����!< +�7 %�����T�N����F2�G��P��$v|�o�.˓�3|�<�S?3�m�a��6�T�I%m�C��h S�	e��ZL9��+�Np���
3j�<?��e/;��� '܌��KM˼��"��ڰaÅ��aAE�5�jxeoo�n̍ԑE�XM��>r�0u����Sӎ6���؉z'�;�BV͙�R�Ң����gf�[\���k:���eׇy^+�j��aN�B���E�ߕ2-ޡd�P�dh�&�[itt�&#�e��ዢ+�d�<��T	�3f�V*0
�K�'1nY�h�H���RE�̝���s�|���9U�59��e:M2���c֙LC�Ӽ�i��rޱaaU@#h'&������3_�@Ke�^G��b���	��p���8��'{���FD?`o+�WT� -�>fgYr�O��P��3T	�-j&�~���� ���t KС�ؔ[%��u���'��Yu��=(�Ȣ��4h�<�乢�Q�0��{������)Z#q5N;�Pjyݭ��4�~p�:����G���>���-^��;� b0Oө���44�a�U�)Im(� [�F� �*�+^b�`@�]�o���U�V���)���/�j9N^����ޟ�����?���?�q�w�V���zMP~|Q��~��6y�(�v_֙4[�0L��0C���F��?<��߹����llg2L�D!e��ܓ�~+�:v,a�E.�3-�K��E-8X�)U�)�@�'>��5_���}-�D�U(:����x���M~�C�	/�����xw ϕ|�M7}�3��ԧ>s��on�ع`Z��h���k_��5�\s���ނ�l^q�p�;�9�A��Y�J;V�y;��ZopD"���gi��e�k�5���7�fK�fCe0,7rr ��v�F�H��"��d�Px������@8�ǹs�,q�p�X��&1a������ע2X9(�A�a2���&�P�(7@��Lc*E|�H�ߠ���*���*zV������.l��65�I�؆�qp�m(Fo�����8�¤�da"o^��(�n��Y)�ߥl� Yڢ���}UD���o�.���m�W����ك��;�PZ����t��K�ޫg��X -&��~	��:�Hn,N�'���)� ~�**Ig	e Ri�0�5ݐDH�d�o�r� �ZmC��rM���Q��x���x�{�g�:�i�Q(X�4�6��;{�-���Y��N�:�F~����w��`�V�%�P������qٶ�*7�U)�)�,��]-���c��A:��լ�U_�4�sLC��Zyr�Ǉ���kMF���#+V���m���8٪�x��S�����뮾�Ui�����É�m�.�6��=��cO�r��WBI|饗 7��F��3_��3y܇@��mK�3�L�Ũ��˵j������.]r�%�V��3���hΗ���h�ν��
�I�:�����K~�<MnJAIj�;"+�� +Z�**1�t��� �={���>�y��I	��Z�f͚� ��U��;��{�U�>9[aQ��@�$d"�Oi�JA���"�kdjIg����8?U���D2�-��Arh��Rm�-5 B��Gq5>k�#�S̊��DI��AcP�1Uu�  E�Eg<e��@�;�bQJ��l������+3@���93�E{SF�&gh[M]3S<xr�!�\�X��2�UkcIƅLd����Ȼ���64m����@��x�'~�h�G������V0�p|ɡX�|�b@������4�����1�a�C�7ڋ�,�00Jh��_~i�._���lz�o��o.�t����|�
�%!��A����T��.�T!��4�R��QPg
53��5�r��rM�`���N�N+(bN��jW�s�+hʚ��DУ���l�ese�
��TWYS���0�M�Ѩ���b�Zh �yC3W�X�c�GJ��e�V'���HF�0'q�#�obB����t�~6Y�ĕ)�A���e���7k5��_�R�J��d9��+��Ŕ�$�UC�I�u@3/�Y[��3�J �e�R�@CP��JC�Q'�10�Q⏀sQ(��R>�M
E��r�A^�	��DηZ�5��A�ԉ�Ӭ�lٲ�Z�w�/����!ISr�E�\fvt�Jq��"�M��<D������.t��i�j E��,k��Ȉ
l,2�E�(���P8���5W�$Sc /}+Y�����u����>������?����"Zom޼���H\[\���n٭Z.���ΐ�`J$�������,�*k =����ߺ��ڶ��������XϕE�>�ɿ��oR�o���tuw�Ԣ^c۶���G`9�s�=�}���x��7\��-�\$Nlġ�k���ATؖ(&D�L�Ό�ڢ��$V�	-ڣ[�$�;�g�F6��"@z@H�p,�&C#�41���"��, 7��
�.��4l=�+��l�p����q]'c�F*��
�[�����_A������_bk���B� ��9�����;�m���ϯ޸q��M ߣV���R�1_}O�շ�m�-7����?Z��G�t�G��u����KH�Ҝ����4�4��_��y�����ύc#��ᱲ�ؿ��_�y���"˶��چdxn���U�V�__�K�G9|%B�U�4̀H�9���2SZ�����E��7�L��,�v���u&
\"������~���N[���n���'�x��g/���'N�⋾���}�9�v&U��~��_���~U�*��5k�[��Mu�G)�C��-�|�s�u��$����� $Z�hRi����18	::|f3-|Uw=зͤ����pF�>��d!K�5��RO'S	m���A!�J�he)j�0P���aXV˪��ȑ��s�']0�FD4��{p�� �aL����G@&a�0�=�Y���8p�jy'N���������>�I�"���!ηf�<1zmZ"�y837�h
��]�h���h�Œ��ӳ���ǩ�_~�e��+�����_�{��^x�*�à�� ����[�n���1�l�JVtdHWP2
or�h�0d�6lh������R��ܪ��C��~���c���ӝ!j<=�f�K��jXb'_#�;M�0���x�'Y2�L�μv��&�>���+[��^�;vؾ s�ެ��&��xUԝjn(�@�d����1�{�jU��jPR�!隬qgԖRht�	-!�O��8Yȋ���`�!�(���m5??��t�,���-�~�g�� '굚JՍ�s"&+Q��D.ۂ�c��j�v�'msz&L�7��L>O5���N5���L�0{���0��2�㉛��,�I�:JR+v?�e�v�$kd��99��Ϟ<~�V�ᙙ�ix��$�eR��t3:�(E>�٪��*~ٷ�P�0ϣj�#��g�A��YGi߉D��C�`-,ްa�Ν ���X�,h��e�Hڑ'/4�)��Go�S�iߒT@�E	=QV��,�!ngEQ�y822g�,�'v��+���:(۪fqv�_�3�Z`�`Y� ;>�{	Ȗ��K�l�SZ[���k�R]�f���W_ug0ld����Z�����{ Z�\	1�þ���0��^zi���X���i;��&�S�4�E��ls�<t���U���} 	i�?�nAK8�sb�g�@�%�c���0��\� gi+vh����q��*�Ha�0Y�d��^'�V
�lY0\�� 
]�+��ʱ#0���}}}�V�����0�vn+7���СC�a���Cb�������G����x��T<'y=I!	*c�;���g~򶭿 {�&\�0sD�	
�����>K@�g��7PN0���!es�W'B�c��7d˫���G���k��@��!He"(�O����~;��,���<��e��w�~�4��ޣ��o��o��q����#�&�{�f��6��)������Y�����ɒ��@a¹�Z�Ҩ�3����o�r��,�V�x�dh����PB��	]��g�Հ�z���O�o��6\�4
Ū�����HD��:����+��=������Jq��RXtȊ�'�{�_�?��+_��$D=�O���?����_-l��8������-���,�ީ`!!�AQ=\��gOM�nh����e��n �T6``��T56��"�7~��ӣ���W�T�^|Y�����RФ�n��)�Lz�k,l/pq��g��\�4�7�8"9C�q	SiT��!G�0F"�K���%�m���w�����l��
XlGj�M߳ُ�P�z�!lC��W2e)�r�m��1��C�'�X���:�<4�Gl��b�M�- 9|�D�#�͖�^ +hX%sGV"����~�*�q�5�rED)j^-�S�u���'l���}Q�z���25��
P4��1EdYBٍ碍�힬��*�a��"I�L�J�{�El�,����ve�����2a�3�㶰܎.,^ރ���@73�>
���07Fֲz �F��W�)�5��c�N-���@ϵ�\���i���Y�r��Wv�G&~t�rT�g������Vk��ݾ�{��<0�(x��m������~N7 ���䆼"رϲK=���V����k�^��HaoO�>qh~^?���< *��Q���.X�x}�@�v���Y� m�K7��e8v�'O=b䱤���A@#��@�S�,հ�Lq��"t���Ό�vS���G�7o��拶m�H�Z����A6��b�h��s����3�V�1�>i�*5���O����,Z���<�Z@�8	g�L{fc��E�a'�Nb�i�CWF6���S�.�]����o7��_�6,@w�oi��%�CC� L@\�`��T7#��@&��OF��n*���!�QL8$x�'l/�n.C��p�V�"췁k�N��\����]]ȿ���z�	[����\��Hr�n�ڞ��n	�
�p@p9�e�yQ�-\�冪�SU=�������HP��ñ8�_��l�Ƌ	A3��׆��Aښ�57 UC�uv��713�i��}1t�Cg�B���^�)��� ��j]��`ݠ�Ì�0
0�,_�:H�d��ɱ�'�yj��0����Q�����[:Ѓ�����{�]�vu��
��|ds^U�,�l� ��躈<�]T��-j��ȱ��HUK|% oa_�kͲN��Ӥb��/d ����C'���F��(bZ���ϻpረ�_r��� ��''�V��=�s�c�=�������%�ܬ�7vy��O��K�m�W=#g��*�H�[P������5[��W������qW�㣿�{���@QD�sՊo���׾cݪ5���E-;�v��=���d���oM̕�O^=����z'����>8s�;��ر㥗^\�dŪ��N׭]}��o|˲-��%MUP>5�;�gs趂�l�0U�����).��"U�\�ᕂ	Qf�����T)��u>35	7,�ȫ�D�F�Y�Z���h�I�T�NBB�� ���'��Q��	�&*�Ԕ��dq��ܜ���&�rzq������<~�剉��O=���:::^�}P��#'�q��.����-SS;v������`Vh.�C;��3��dͪ	*rc(�&�
٤]&���I�¾����i�J:���<�0���o����_�v�6,�$��e���������	ؾ�$��#/x-]�Z��,)}�F:����^d�۰�j)[l5a5����[���������o�p�"Y~x˭���}�#v
H�	J��-YY�����}�1�F��~��g�}V7В.`a:�*kȹG�IN�+b?y�
�v�9�jr��z�"&E��='Q�,�/Mg�ߪh�#/bBJ�w�(�e)
<�_�Ї��"�T�y��#�iAo�$z�/&t��;<�r��,���:p�Y�dө�<�U�V�"�\2��k�����^O�\ e��_��_��Ǆ8k�4�˷�C��YUPS���M�P�C8��.��Z�c�<��Ѵk��o��·��Dc%cR�:b'�V����=�o��������t�R�".���5���~��?����3^�-��	^ur�U������9�M�@�8�~����}b:����/|�M7]�w�w��ԧ:��]_0�瀝�v�С������lF�1��G�D1G�R���S<AJ�(=�ۄ$c*5��	��@���{���u�J-ă�����~��Ɂ���|whhQ���s��2�$KH~�>E�r��L�ק��D���b����Y*���"W�b�P(`\�G���Θ�����6�B�.�7�J��$Qq����M�6MMMu�.��7n|���ڻ}�v��(/w�F��+@G뽙9N��'�ƹ8n��I<-�m��iX-k�ef�K&f0	�%���U Ƅ۲v��YѴ�/�.��?|t2��.]z�;�}���?����o��&C� b9:s��dd�����5*�?�w��F���H�:�wäP
#8Fc
��q�]���ƅ�W�6f�CJ������"��>� �Ԇ��-hJZ��U�+�	�/S��<P�Z�2�����(lݺu��^|�ŀ���ޝ{v�X�r*����Q�<��Οٌ���H���	O򔠟m�|���T�C8	��X����CCK�j�r3[�^ '�i�#6�e�Cqȓ�p�a)���]s���~W��*i��۸:S�H ��F���"2w!w��#�I�CWv�b��\��(��Z���v���$�b͌�����E@�* �%K��Kr�+;a֭[�
��u���\���t&�`횑2��`���*�w����+a�@/&��b����]��83�Ɛ̱`6�҆���(��&|ulb
-,=]�o�-�`N�F�[�{&�b�X8����zux���8�@�/p���qn 7����=�˲9��\9@/�o��%=�Z>g/���Ur9����O

��A;a�=z����4�y�{�O.��8
o�p=�v0o���?88x��Qh�{��^���prz
�7l��Pyh-�:�Ѫ���/9��A/���$ɑ�U�z���u��|@Yya �jewV$��b�of�-��H��d����#'�#����|���|SGkH!�c7#��ڕ���@=q�ĩf��n���F[O�b^�hϞ=��Ls�ʕ0�����"��������D|�2?���{FN�����%��Ϭ׶k¼6P�;�M��a=+��⩒��^@bPU}������/A���a8��G֗�^V&_��W���S��9����s��z�MF������hN�=�ut�����Q[v4�lR/M;X�)�v5/h��ܮ��_�����3��X���o���b�3��㟴es�D�xC�1!4%q��kq�������O�x��1�t�(��~�U(&5����-����ᐣ�'UI�����0�����.[���~�������;"]��Q�$Ay�W.�|L�����ǟ$wHĮ��/�_g9��[r��K�Pq��l�:���ݢ6�r���=����:���HJW( -X$J�6��>��G7myۇ��<��}�����~�V��B��xұ��0�J�T��n@�f=�J�굲���+�	�v9E5s"���@�#������b*>�%�>VO���\�+��C�z&�ɣUk��]q%�\p����_��
��ıc0SJ�<ݣતs�:fL�qA�k	f��!�Q�}+!�t"y�u��<hW�2P!������0�%'V*#�yd�X�dp���@e�]3��� �-d��z���u
��<�j:�l��J��fxq�V�u�~����^0r�֬�t�Fؿ�*�7�]ݰ���5z|�h��*ߵZM�vh*�PX��,�r��$|+{qM̺UsU;���ط�00�Q��Z3�L(e�� �|1�9)p��A�'��rY�h/z�/����}G�y�Ak�����k�9u��}�gh�e[곘u6�D�O��An���R��=�e�r�P��>Ա��e˖�==��5����6��3=2	�uf���X7�G
Q���]=Lδ`-Y��#��&`&\.�d���R��129=�d��ݍJu�� D?}Ǯ�8�e�Bg*�&|�d*͒b��<E�,I�ω�_�b��2G���vS+�!���&I�GU���bE<����@JP����z���{�ea� ,$���d-@ǧ"c
!ջʀ��!YG�~/�	M%�ŪIx֮��F�g���}�*�&�ck�U���F�1q˵|��� k{xp���|2{���Cr�4�R�2k�Qd~������a�J3���C%��I� z�Ztj���5X�����n��ۨWay��U��m�2��Ƈ�{��[*�2�֎��,�U0���lM7�9AAl6��[c3�]CN���A���f��6Y[+�gh��	Bcv:#	݊�~p�$i��B�e؞Y�)��*c�}]�6Y+B��,i*��g����I�T��Q�l����g�0�+�ֺu�׭�ܳgǫ��]��S�U�ȯ����^>8,a�$�4і�u<��ֱbxwO̅'�|
k��r�Lᆇ�����K����<�X}��bj_�a�H�|�7A�#�"�l���|��͚۶m��F������*��|�V�-(�l9�od5,P���*����l����r(8(��,Ȧ��-@
5�G��iۢ��^1_m!�g&7[��\���ϭ]ڳ��=�/?p#Ϋ�Ƭ;wb�D%�2K�g����C/`���-�����G�m�]���勋��n�0����H[��r��������^T�R�->��w��8�#22@�������4�m�Q��0�6���"~b$@e	��cs���Q�5۲t��#�0��e�(<��D"�����-$sO$p	��c�����i�~R%55���� 5y�<:Q�[���|�ä�1S���-��g�\LF�]͒�N3L�On�t_ē ^1�j�;����	����g��՞[��	D>����^C���x �l�[X�4�*�k+B�jV�Y��������g>󙫮�
���~����z+lb���ޟ�ٟ�����wx�g��q��|��uAB�)$�O��Z����贈6�>J��S����iSS� ɤ�Id��~��z���}h�֭=X����u��n`K9}�(��Vm�L_��PQ��vmC7|���	?'��dԤ&|���m�[|1�n1� E[�"6<<�l�FPO�<��Rs�޽�O��,������k/"��|__�A:���x��I��R%��D�V�
E	ôb�,�*� �B���s��5�p:J��˗�����/�|v�S�GO�:���{��@cPL�k���l��X ����go<���ի��=��6lX��wvv6�&�J��/��R�����a��}���e�_ɪc}�
yk���U޴cY�+C&L%�m�nR��TE�*:D���^f) ���i��kϞ=��߾}���@{.���\s�S�w?��#�'����������?��SE��{�,�7�+��젟�y��"4� @rp�$x_i�"@�.������#�@�}N�'�x�~���ݻ'�B&#���6m�f����F|-(�2���;J]lk�&vv��8<;��0�m�
���<9��p0��)�I$��a�@à2�F�"�|.M��bk�����NA��3�Jc#�c��ȩ��X�`U��n 0�ӓ8v��-�+�šV�~�T� ���Vu�$.�ćK�:,@��:|&�0����H� $�T�T��l_�i;�e9a�X�ނ���E�ېu#L��A{C�E�T�@��)'A�JYD�-p2�by+S�M���=Z�������=��%<z�yS��Dp�Uo&{��E��ۛ����r;~p?V��@�"9@��|h���Kث�1pHd#ù�<��E	�[��-����<Z���TqQ��<��)}H�����}R�����Aj`JF-���\�w��:q��Z&iʰ����8w��� �,��S����l��R�V�6m�t�w,�6�4�yU��;�����\�$��#G�� �>� ���[�p͚5�+�]�;x������eI�r��\����s�l��b����]�z�ҥ���@aҞ9	נ�]%ךUJ+������=��_~��r�5ybx�Q��3�~WT�US\��������3�����Gs95���-����>��*Оٕ�����O��r�j83;62��jB��G������m�z�M7�=O�~�S��~˚QMqSΪ�u&�����g�8�?�*�T�ZH��xT��1Z/�����wv�<��0H���K�D��l:��F��&Ɏ�4c��q�xT=9��Y�U��4T��e��M(KJ{�uT������x͋�w^LH���"�no��]Si��j�˰@�t6�\0i�,��9k7o���U�3+���t������e)Q fu�ׯ�{���~�#����������#�^��"Y�ߒQ����>2�#q2e�X ��<�V�>��J�ѼI3d�ڝL�
������v/��&-��b�i��7⪤I��è^	���&��?��?�eK��xC����_����޷o�֭˙He9�'�g˳�B�헾���ݒ��x����_�r�E���'�=o���4�&^l��b���+_F_�K&�T��T�_���0���%r�v�tu�8p`�à1ttw�NN@'�TZ��/�k���.�R:�23��n��Fm���8|���+�����a���L-�����-�V7�~�3�,s���uv�y-g�J�=�:̓��y��j�Gӣ���zs���J˞̠F\n�y���VcW\	�-�*���|g�b��ӣGv���:5��&��;��������@zn�vl�.kjv�T��x�>�>�1��Q�2e.i��aUa%�w�Wb�h�k�j�
)B@� ]n���'�F^Ġ�x�$(XÆj�3W����̞:�dɒ�W�c��ʋG�?~���+V�X�|	�DR ��G�v�� rs�.@<}��呟�"�~�hZ��� *�����������W�̲��v���+���bP��ڈ�e�� ~*���kG���ҩb�LH�ǲ�*�*��Σ�A1��n�m��bL���g���K��^��.��9I�*�X��c*3$���^j�U���
��ODEub�Fgm�Fm�x�gېm[�"3�ae���DJ�衠�q��C$F�D`�l�v��v\Pd�����q��r�ۤ�3�.���x�|�Ǳ]�#�'�#RS%�]*
IHa�Cb�XIH��Q�3
e��Ō�+�Β��N��B!&�(�%�����a��ˡ@� ``Q����b}X5 Gg���@����oW*s�.��Y�Z�0�X%����%QhA� ����jO	k�M�e��-Z<5:ޛ�;�)�*	�c�-_���low��cπU�x2Q�z֝Y���R��+�#X�s�}�����FKB����u!�n���:f$��/iJ$K>f��;0��������:b�_/�;��$�Ih[�݄n�������[<�lٲ��VԬ搮�\�*�����̪"rE�agc�ـ~�J�qjhz>0��e�oQqQO_�ިL��"$���ج�b�R�bu)�׺�Q�#ZZ�cW�p��M
9�i>����=�Z{mzFv��ĄY�8l��5Ȋ�r�\.OLNl��y�Zoa�13}FE��� ��Ĉ�r�
9A��^mFs�^�s��Aa�/��Z�����m?���8���B�;�]���CpF�-eSWBW�۳V�ݷ��+��c�O�:r�hA�d]FDQ�u02"Wx�w��SK�����>�&"-K9�,_U����W�ࣄ~�l̰��Y�9���D�!��3�A�kzp�H��>��G�jd\C���5	9�P�F{J��"�C1��c[_�a$�U��axqqz%��BCl+�ގ+��Σ�,VrR�0��O���#�.I���=�S�'��+��L:x�/ň�wdlUΠKD9d~`�ң!��J�����I��+p�1�C�5��\mמ�޶�?g�[X�^6�A@	õ���w��}�u�uww�M��;���o��|p��aAc��(�>�˄��rLKz7� �(8.5-��I��L�y��gI
d�f��6H^��s8]~� CD{;���1�����޽{?��B'�����'���?��?y��?�bPX�i��������QL�\`�~���|d�Ï=����������.S�g���y����j�������$&n
�
#��O�:��/��[Bul�Ӗ.��X�x���  ��2(���ի13D�́�/���Z�bC��}YM�sFE!��L���H��/�)���˗�{[;�a�D��n�����/c>�,B(�WFGGA}?v�X��'��ة#Kx�`^+"$�(�Ks���'�xb���,Y2���{��}��A]#���!=�/�v}S�2ܠg�좣U�5�(�Չ��,OW��b� R�>�hA�xә�7�&@&#� ��� C�cǎus�pf�x�)���?>|����`OG7��R2SS���r�:���E=�8�C�� (�p7;�I�N�<Y۳�`��829�c2�
Oo���#+��RIB�8QȠ��_��ܱ\�p�BT�tҒ�gf�ɭ�K����-�;1�t׮]��v9��d��\�jյ�^�ᢋ.�䒺��������G�~�i�*���M����y�`'Ή����2)9��%!�d{*�bkEEnʄ�d0�����S-�f�R�@w���	t�jG�3TCF���%�`"����C�uN�T5td���!�Vcͯm٦����Дa�_����h�-�arT$NrQ��p"X�\M�+/q��$ƙ�lA�$� k��,�Uy饗�~Í���v�	2�4Ux��E}($�X�E���?�c?fmy�֓O>	0��!���y:%dJ:�&�O�.�? 9��\#����L���7222���;Td��=����Zv;��#�Z�v-#��k@JL�O�z��y�ZRb/����Xă�>[���	�NHq�I)$�����<�"t���pf|f����5Ǟ��n��s�e�m��K ?׮];vpl�ƍ�Q=������4ouw�`�>|8 gZ@���0����fgg�{�-�֯��
<8�� ���4�y��I&���O�4N�YDȡ���e<fᡍ�􌦈��m��Ek.�|�p}�2}R��P�W� |*�:4��#�l�Iu8Vx�2L+Lg���S��uW]�iӦ��Z��֬y�K��C�A���l��������瞛���F������3�F�	�h��ܺu����n̲k5`tK'��i~c$Dgm��9ks<ߑ��� �@Í�H�tÀեa�`�|�x���Weŵ�U+��
�Â"�E�I<��JE����i�1�� ��(1�i
~��]�-<��.�H=R����C�E&H��W�<j�?&F����Ay�0=�+c��v�xV\C\HC��ř��'�3s��F�4z�����z�C�T���mf!�]ڵc��\��;��r�][�t��@�7������ٙs�HUA�1$k�8�!7��m~�םE,v��[Y�S�r�Ns_gAr>:9x�H?�%�1�Ϊ��)`�Z="Z�>���D�{��_���	���K���A�fhɶ/���O�4r]f �&k�m���?���|���1������o�sߗ���[�������#��ތ��,t�D�!�/u�G`<$�WlB��H�`>i���(z��#��l���Շ`z��g���3W���tqrr\��v�����d��h�|7�.�]�.kfLCk5�Bd��.G�Ӝ�ԬkY���6mO !�2�ΎlwO��W��T���;:��0=:{�@�${��Ij�	�ޘc�0�#K��W�/c(5���R!�,R�/�Fvzw&{�q���L�xvÞ�鐤B1�kFx��Y��#����Q]�Ƽ�� �ԋ� &��"km�=dY��! �O脶�)�����S�?��	�HF8����PЕ�Ĭ�I��ý�|qX�"��������K�l���돎�n߾=�n��4r�z�!ij�#�(?�O���s*����"}�(yn',.�nFFf%yb����C�H}�n�`E:Vːb�2n���uKә�ƪ	M��U�4���I�!m�&Ϊ̐:1��*r�CLNO���:~�/��?!Q8�q�&��\]]�R�^g[n�#�.��M,�L��mڶIFa��ђ
�a1w�+���`M7S����A󯲋�� �̌y1��Ԗ�P.&!�� ���0TI�ҝ*(*��<b���v�6#(7��h��H	5|�d��{� ��J__�Y��u5))P.Q�����Va�]悗��W�ZI5Wj	�B("#���U����wr�o�E��� �$�N����a����-�}S���h�`|�lj��l5q� ��P�`���b������m;4���l���>U��*d�kh������xu:g����Y7f���a-�5C�P��r=�)��VM�|�Y�+(䳎ݪ�ȟ��Q�O�S��[Ȑ�-��P}�b,�@C/uP�����j#�5��9L��k�W�@�z�ś7e4u��U��đ�m�8U�����7��B�[�c��Ra����X݋�� G���3�����
P����{g�'A�^�hX���2e5C�l�Z�'�H�N$GYDڪ��Q" ��ëL]�hpI25�RЕE�EUp~��[�������e0�-�8p�:q�^+X�{�{,@�-+a¨�*�'��߰��8;u�b_���Brbk~l���X��;l	��(��a���ih��^2Ϯ��bid�"+Ӌ-ו쳏?^��[�n���}7������Pm,�����UW����ۃ�!�@i��*��ɳL3���?�Ӷ�(R&^�IR*氃" ���7�x?�W q@$�r��DI�p�,��R�%�q��� ��� �	�%E#&'C�a�9�Q����g���OEDD�|�)��}�F�s�)�2ZH*
���EX�RRkX����N����(�	W8���C�m�n����	���6��F}�s�X{���z�=q%CN֊��b�g�֥��o��xf;c���M����oa�78��(�9�wEC���g?�����n��;X��}�{�_}㯞x≛o��H�.?p���c��9�¹1ǯu�m��aM�Bb�NՑ�<X]P�l9��W �@�MVl݉�Z�I;�;�1Ca t9���#��P~׻��F�ah��Z�'�_�����/D$�������G�&e�b{���7^�x��'Au��}�ˌތ��_�8˵%��!m�+\�1J�I��[j�����iv��c#��Ț:??�b��ꫯ�/Ww�ڵa���{�=zvqEG�����~щ���/Bn�dΰ�3&$Í�;DKv$b�.���c�	y���33�&B���ߺ�
�#��^;�����:�9��Z~6���1<H'�=n"��4#��!we ��
�<���p�נ�����!R}!J+��Z�R�<xIvn�s`	�C�m!p�c�7]�օ�`�.��+�� HH!k�!k-*We�D WO=����K{�~������٨f��G�¬���e#��Hf��B�ЄѠ�<&�)X9/;~���!'[^ì���Wv���(IX��7f�W���s�0�QT�"LE�N���'�J�M�D��� .?~���\e���6����ss��K���B�u)�����j7]	�Y�������p�g�!EV�:z�(t8G�a6d�Q��:��ٴ�% �8����B�:I��gB!��s�I���Á����DmSsU<oè�}ӷ��9���T�@�5�M  �ɅL�&��5��I��O�X����&�Ar ��u��
���
-���Y\� �1ϧ�@B�r��q0����QpB����!Z���0����|*t�B�����΍C�
u�D��؁��Jc���]�T� ����G�b蒟K�H∛Spr��E�ߒ��6w�"����O{�O,Ce�ʶ��I1�.e%)RR��Z;����ɓФ�N���T_G'b�Z���ܶmL�x @�R�<�u��C�/�~�t�Rh���߿|��[n����p�"<~�I�bB����:����86�Ī����"�:�����!'���	��r�J�(#$�s�<	=��߽aÆ�����-[��/�вC�e�����'�Gt�g�\����nݺM�V�(<�ēpO��MVga?��wTs�pg������'N�B��o�566���Aʹ���_\�d`�ٹw�>N���/�^�9�[?�U+�$Q�{�ׄ�/��2e�\��ǔ.�"�{hD!��'�b�kUR�=���.�# 2�ĕ��d9�+�����4�������C�ގ?$,V
�K<,�!Q��P�v�����*B��_�u>U-Jr�����K���G��%L��>}���Rv.�l��U����h�჊7�������5;�e��΍��ܟ��-��G$P
S���|��ib�[Ƣ�!�ʙ��z�!��}����o�7��f����LgJ � ��2<+����z�3�x�Ii��Oܪ�
+�-�׼��䕶_/�����>bN%JXhqO�D������ON΋jD��T<(�dA՟z�q�qs�x!�*ն����p���g���R���̰8T8�b��3�p[�@�qbO��۪j!&�H�&��wGA
���FH$�2n��n�V�. ��d�՚5k0��i��״�=����:���T���֫Tf���1I֑�WC?��5L]%�
Y��s�&�bӔK���c�]��LV��ܔUo�:l*��%{v P�ؑ����7���U��� l��� vD���EM�hwm�8�\�6�0P%�K�u]�*b�Zcg��6<�@��	W����Cu?�$�y�+F�m/B�'IhSTx�
q|&lE�`�Pd�k�"S�i��V�I#����j��GU@B���H�yN���s�V�7X���O�:z��1"-w�GO�>0�qO��X�f.lYNK5tM4��q�a<&T(
�蘒A�+��G�B+�C�F ���}����2hb�����,4e�WPA�`]�h�TH��mzI�rQ�eS>� ��M�V��Q��Z���������z����c�=�����ׯ���L��=��u�桟�D�ͱO�d�4C ��/�U�&F2�Ql�I���9��!��w6�¯��|�%&2I��$u�l�"�G�B�F��a���1=6��P�:�;AV'''�Ogϣ�����ǔQ@���tN����0UtX"|�1��tk�e[�Ԙ�U�"��B��p>-D#�1l��M����Ͳݲ�����4 ��Ƽ�K?s�Em45�Y���0�U����S���V�9M_�j�O��9��.�a�x>ȇ��+EDY�+�57S�W�������h=ܭ̹����T�+P,��k�靵"� =�U]��VV����6��S�U���_�d����呶<���1�b�:�CRe4��
l�A�h&<]���s���y��������01j�q��-�;4v�x�n4�{��4�e�	��%Y���8��׎���XVPIϔG'�s��c������*(�v�՗^�z�]h3�a�aj\�0�+ջ�`L�%�NR �C+��D�G�i�ڕ}��(t*�������A2�Ŏ��v�\�f���Vm�����������O`
F�-D��9Z���m�j����/z����w�	D���8�p�p?�S�e���a����5lk���P��M����G��6.>���ӧ'�>�|�D�661���w��/0��i��+
y�j��?��m�Q\��\ﯽo���4Z��`�3!Q	��s�)R��A����6�D��A��/7G)� Z`h`�G��P��Dɏ���Ab�.����
1@3#�X�L���D�1R,ĵUXYiנҗM�ij���%��\�P	f�f� �\P��1	����*^\�>�(ڈ�R�����J1O�PCK:�t%�2E�y���!u(R����|�HL��C�|�^?TpUd�����-"F�x���!U�`$�3�xR�a.�ɸg���d{���W���A8?�}�oa�780�RA3���>h�>HW�6E�������9����nZ�F��S7���-�B����5��8�Jj��j7Ո	sj,a�i�h9Պ�����w���ML��SV֍p�=��'�XїBa�[����}�0��N��u�"��F�����=��O��{�]�<�ԎB�/�`jY����B#7�� $��<�v<�Є���-�R�PK#���̟��WJKg�AR6�#	��6E�z�*����A\h�aV`�+>Pz�3�<p�}��<!�ؤ���I3�"r�U-���R�~ Ss�LSUTIP^���l�R�H3#��F��W��EgT��p�9n	n����A!wsDUb�0�%��`�`�ΐd3h���K�m}�9� ���:M��e���g���&���u̐fFƔ��j����En ��e!���8�G����L����MB����p���,���[�J�{��C��P�i����������D�8D�693��Su��m��~3J}f��R/��q1�HT�ۇ����a�kXI	��g�O���	�xt��#��#����|�������6�Ϙ�	������g{�,z��ꀘ0��0Ȋ��H���P(�£+Et�a>A��l���"u��I�	zd�|�/��6h��}�3rs]�]X)��Tn�̩G�$�1LE�R��wg��&k��� ����ԡ�)j>z\A�A;�i:��������Y�v-<}���7a�g�Y޿?�����t~I \H�"IUñ61S�&"�;g�@�+3�:|���s�g�T�����)Җ�3諆�5�����g�9��X6������1)?χtudt40z�7b�
3�odѬ�,h��'N�p��ֻD����
�3�bN"&m�ւK}����d�8��hF�!8}�t��,Ӯ���T�0a�B����]@���p;v�S-��;�b�1u�V�c�;���xZֵ�+W������2q�Au�X��	�U>���~d/����T6r�tb�@�#�Z��ŋ�f�ؓ�Z��?9>>�>�E��5�� �C�\/c=�VǺ���
^�?�.��4�þ)����� u��pD�E���k*XF��^u=��<�!|K3��R]H0	��_�1���E�5�R����bY�t,o6�F0FfrX�>�)\ �"�7��Cl?q~�d;�dx/jK5O1��B,?SuΧ��.��@�|NAZ����<����b�''�I+$&{��,��\5� ��$�,��(ۮ���Q�$$����XkCHV1;!�9-�	�PX�0���Ƞ��qX��ǧ�.M��)��>�����F/q=$җP�l�H\��9��GV�oa�78tل�b7�B���{�Z���l�P��֤f๲h���o��?��Ï���H�¼����b	Z�S��"F7��h&զ�|�k�/^���/E!	�M(9#K8S�OoҎ�8Ɔ�gj�/���K����j���.�,�+Ǖ�9t���޾-ۑ�d�`KLХ5�ӿ������C߹�#���\�=�|��;������LLO�y�/>��w~�w�Y���R��V;�ћ�O�B�]�*�m�:�d�%�Ȼ%�(y�д���+�Z�qQ�!���}��ݲ�"�t��,���	���.����F-(���ȜU�;J@93�+�7�bd{�c�N��0<ԓɘ�M�������
h�,�e��9�ma�Q(X�cS�}�s�3]}��W�Vյ��xT��%�� ��K2h�nro_�X�a�We�&%����}1"�WB1�@O��e$=��a��0v�ZT�7V�)��m������Ճ�LF���m#�P��8z�( �@uاJǺ��H�� �R|tMX�X��>�}��<��3Wm���ĉC�S#����k4�|�Hc���>z>ećhm�#x��rK"B���AP'�Z6c�p$��,;��K�9>b$M��2�GjG=�|Q&��C#��Y�7m�qd�C����Ŏ�C1_�8�Z�R�����̌�?��#��_ ��P��0Ʃ`�0M�s��5�l@�wg�_�a%b��C�0���@��R`)���6e��Q��ĄG*ä�tR0�#�<b��H ��G���2f0��a��B�z�ZP�e8V�L4@�9F�ͦ4��� �A�;>����$��9�UB���t���MbU����t�V��ų]g�sp�|.�Ѥ0
�V��������� �b��9�b�;44K`�@���h��	{����H簺-�]v�]w�t�Kܻ�UЕ��>;	5� f�Z!��M��tARr���^菃{7d�;>�|�A�XV��_����S��]�2%3�jѓ#c���'�ۺ��X���<�V�8ͧ��Fg�NC;�
�S~] `�[:V��W/�^�-��y�j5ʵ���ǎu�"F�$��%Ј~X��� $8רȨ�F�j-��g{;{0[u��/;O��XEWҔl1�k&�
��rd� �ڑU5A�|b_}W�����P���T���Eq�y�#Qv=�;��ZI��y����Gd�0Z�*�I#�J1X7n�<A�>�Ι
����,�i�j���S;��&����e\�f-{����S/]}�,�l�����̖�1>�Ѓ�<<E�3�:��o�@��GF���;qj���1}ֶ��S���L5�Y|�%�Tld:Q�ʬ"Uݲhhݘ�&[�	���ݹb�8N��	s�w!�Q�ˡ�)\ER@�� ��P�(N�l�uN��k����%®���;�t��p� 
F�(�Q��5�c*�/ːU E>H����T-A.�\��nY�_0��=\wN�5�uU�v`XU����C�CHG�ff�I��؊*�o^Cw��Q�����m�(�y�����5ڭ��g�e2�����["RkczC�Zi2t��������6�8a�;��X����yHv)H�W��K���T�O&�2G�`ͲP���U��7���z�쑇�9jM��Y�����2!Beh� 1�>��U]^j��`
&GFJD��q��LdHZ��$��5�o���[X���Y^y��ӧ�_��aI;��D�8��p�֭���_���~�.4P	It_�E<V&h�i �`Y���dӧ�m��@�/f�Hj;���ilLzq*�&��u9���m��MA������vE�M�������T�w�q��P��I�l��6���o��G���k����o~�|衇8:.ia���_��Xp �D%<��{(K��N�_�^��9LO��	�f�P!YȒQ !2�>�cLв$���1p���laY`d�D0�9gi�49t�t~�r��PU�f���>������������wC��9�_SGfV.��tH/�{fߌXd�>�S�d̑Ïx��H�3g8L�rߋi�yA�]t���2��iZ9��1S�O�¶c����.R���_���j�����7��(8> R7'_T.�W���&у4k�Y�d���]���$�n���:���Gi=!5�9�t���b}zz�_ ����$�	f���,`-��D/>�`� iy1.�"R�L.7 ���X��31�F&�B�/D�"(�(��̶O���ĞK��	)x�)O,��yV \���s9��X�Rk4���Yb��ܵ	�������&l��!x�t��#J��4�t�\�F:�i�jo� �h���?��X�z��H 2*-�E��)���w�of�*N=әK�˓��=N��H��T�����`جᐣHm\)-6�(2�b[�����5]
���KJ��O+�J0�H���m"2�����l`���u4)�����E��bf	q���m��L�_
(�0&q������a��Ν;%�v���{���� q]ۆu��1����|�V�ҥ�k�/`W��xr��9Q^�b
I���r��j2Z6��0%�l1D�V�HN������8`�P�7�'b6�	D�{�i���3���n�o}��i��m"�V쟞׋�P��� k.�Kq��!���iL�& ^����^�ʰ4��q�^��u����	TĎHI�J�a�H<��N�mi|��.66v����]\�8�s�>@�����eZ^�Dt̒X�V�r�%SJ�c^��B�G�J�,�8������i�)�[lo���p?�r�ir��FR̖7��R�^f��a,������.2��j�7����8j6/���I\�Q�����yȽȥ�`^���k8�*��;GMqʓ����ҹ��E��:����)�0a�	�fD%�������ď󓹔VS�8U֦�a6�N|��^\W����8�P�^>��Դ�X�aYq���r����������ތo��e��T�&��\�S�$�S��P�5����Tl
��ǔl����٪�)#���L�<�TYK���j7ԏtfΐD�M�rD+��2u'�-�;Fɉ����ryNs��wBH�ꀗ���xk��qUU &�����\E=��o�ba���"dUk�����?�Х���7���/�P�:���XWM�4]*���lǅKVZ>j�t�=�F/����qH����~�;*q��U��YErZ�P1H���J�w�$"V�Da'�������a�\t�;e� �"�������r�]w�}�����7Ȇ��_�µ7��X�[�������*Q޹�K��(�ߓM�Ҕ�;�ÛP�� q�P�{�)�͉��PP��@1�ɬ�n��˔� Yj�b�T�n�ի�rav,i�˙ydG��[�H�E�0���� ��HAӵ%����V������z����v�1_�A��=����c��N�9���.˥�@� ��Xh��j�14����~�Ĭ��t�n�v�-��]v����'�]��S,�/�%MrY�����L�"�%�T��"]�}{�9T����A�b<�,[ua�ը���
0���=�����G��#mp`t�I֯_h
��2�R�##���T'�b@ t�^?�s�=1etu-1�e��q�ݾ}�4�w�E�9����<i�������j���J���.�8��F�2I�K�Ǧ�i,P/�r'�6&���-��V�FS��}��'�XS�[o��!a��)�;22Қ=�w�މ�{�Utm_wב#K�VsGq�S�����������{�|���ѥ===��{��.�Sc܂iZ�'�i�h�j:sFI4alNa
��d��؞
�!�G�9E3q���d&�gtAi]��&�����Pu��.��a��`��jV�:�&�q�DiاX(�\>��h�U;0Yo���z����-O���\t�G1�����]���Nа[t3haa(���*�#7�{���\�D�X8-�}�/��&u-���j�ha�J��X�焧��"gj����6�$�j��z�ŦM�6o�|ڱ�!�[@���;ΰ��!4-�����?\�58'H��fsǮ��;��u��n<��5�e�[�>,�뮻�E��w�;,P�)G���Ro��c�ٶov����|�9���be�j�n��!��.�>k+���xa~~�Y��ZbU�@*]��^���9��7!�1�b��䅊�,�Ȫ�����V���ݻ�nv1�X,�:+"OC#r�����Òg���^ ��	�Hľ�r�'�5��]d�M�UD��rYI�q����l&c@�-1�hFL�B�Hf(��fĺ\$�CZN���}���՜ S���J��s����ҩ�曍�	1�(�V$��Zsltlrb��v�~��n,Xyc�p/LVs��m�4�U�=�����J����{�s텅��tx��
G5ë́� {3s����}��������XU&v��_�Ua�����V�Q3C���������͠|3������ԟ�w}� 3~��řz8�O�鈱���FYs�`-�)Y��
v9Z���D����n�����(����N7��¸��b`�X���:5Xw|4ⵜ�l֍��� ��5�M�+EF"S, V�,�U@0J��b>�*�����_89��G>�rEI��Q�|fQڰ�0C��+�"F�q��6K�(����d���k �;S3|��H�}���)Jjh��!!4�a`�	�7�p�G>�(���"���?=��s�P������#W~��ii�؂�܅�Իf�+�.��jG˖������Z�H���o�-r���Ko��f��e�Z-��sυR���uie9 0�i��:
����ݸ��;�Ӳ
"��	�7�=K"��=9^�Z�r�f��*��}�=˖��x�	!�y`�۵ћ�/ap�E}��_��W�r�Ygi:�NS3���硰��[}�<Y�	���$Րq|�Qȣ�9���DRt�3_rV���S�[�qW�6��Ҽۨ�(<�-�ȵ�i���	Y����y����(����+��6����Ѳ�я~��?�	�,X�l������z9���MS1�}W,#X(��l�����$�Љ7]f\��_��×1�B�E�Rh��a�	Wu-K��H�%
���1{�@�S�R��;������,V�}�ځV�vd���*MDB���[c׵ S�Y��p��!�����2����X�Xd���f������!��av�,-^�>�&;�6p�Д���+9�����AVZ0,�Ck��
}�2�"�A�g������Prv��I������i����#�pG1��\F�t0w��դ�bG;U`�2"׆���r&6͏<�H�Px��/���;9٧Jp���c�ziTI����C�rIA�������mttt��e�:���0lv�P4���!8YM��:���G�sf:�8�_�<DY *;�kI#eL	[x����:�4�����i)�un4>�ND�`��)V���&�E�4��B<GA�%)Jn~��P[
����\Z��'�	m�h���m7�b�ȧ��b扨�k3��#.���O�o���֬YW�ܷ�&��������g�ZOo	l��B�??����\mz�` ��#(�mW97	�À�s0�D�!qfr�F�7(:��f`���*!رI{��h#:6�R�pSLE#ؿ��,W�Ф�$̜tl�h�d�xQ)�^R�o�;,���=�+`�$:JpzFK�c�1ym�ҥ�{{g隨�,��
=����v��l��#cZZ���a!I;:��FT�/21P�?�?��.`�x~~0>�Q-ʇ(Lt4� ���*b��ex|�����Sc��t1��aÇ
id������B^`��jd���L"q����q6�!Qq���O��OD7AI����b�/�Rz���l��^A]����?EV���o�l��*G@�?�яλ����7�x���q!���q�bsu�=��l�X��mgݺu�������5l.ר����w��� M^E�·���7|n�玠qԬՎ:z-����J(ԇ�
�*C�g�-[J��K�:�D>I���X�J���ó˛k(�&Ei��,�H,���\����ItX�<M��DY9�d;�B�
]�$cNx�}��s�9h��!>��8
~�%����{�nl�Me|�R�Pk�����4� d���ÏXU�r|cQ��A<����뮹��+%"s��/��x��}�sW]�)|j�ך��<�c�T�
@���~�i���M�ź�����͘�c�W9��S	��B��m��M3Cr���X�zh�C��E~;R���{��j3���|��W8ĺS�ϑyA\����f�U��ea�p��gVG+H�0m���ً���2jb�qe�,�������D?@wr+:lrq�cidL¼e%�Y��oQ���X���ذB���0"�_�5�
�ny����(y2&���3F"n�$?�C�x���O*��{tu��\l�N�d2W�`x�{PJ(�<R��*rH�������F�c������\� ڮ��[fv�j���Ғ�^�P���T���g�g\�#kD���-��P�ON�]9v�1�Fd\�Ҕ�
0�B0H�a�_OwŲ̜Y�|�٧�T�����J%s�Fˀ��i� K�G�*��"���U��F�p(�|Bu��k��|�`�)�`@�a�P�#eTJ�:��.G���|�6
���Lʹ*-'<��K���v���UI����d���z���u�]�����T�1�䢋.����au�Q�p�`r��
�f��a���V����&�6�~�ʣ��rmb�jʑ"��P�}��p��U���m"ǀ�-�VS����ّ^�Ŵuѿȳ��<4�;6�v����v���\WTԲ�]���Nz-?�yG�7O�{~zB���3��e��Eٳg�9<�e�ք{��!���k�۹Bq��� � �֫5-)�\�$u,c|A��ب����GQMr�Ă~-RuZci3Y"����,�,kQ��SKA�Z�Q~�ϩ�l��i�x
��BR3a���z�mT)j��tyb�*�FCr���i))��&cڔ9ͤ�S�0�a��P�s!�ˡ��.b!RzJ��X�~�6�ou>�]�m���O�/��)T�!X�`^&�`|��Ff�e�]6T������ݿ? �][[(�m��`އ�>��s�s�م���������u��c���~TX����|Ė�m��/��_q䪰:[c��(Z�M�0�g��Ȏ=�k�����/]h�ž̓�\8/�ֱJ٭��ފpm�!��R������"���� �a4t�@�h�t�[�*_�'6��x�wLOL��?��cv�b���0�QSa��֐�W�QVE5��	�*u���/�0�c�:�!י��J,<0�Qdc�9���Z֨n������9{�0
�,�۶�,$u\�-�ba�z�`�-t��;*�8*�K��BS$;t[vN�ܭ�u�(̙���^M�.mzf��&�!���,�'�n�Rp�D(̜n�ZKj����@+hz^s]ZX�R�10�u��P�`}ԍCm!��R	n؏� lé��?�A�}��_�\[A$�eh��z-�}�hq����I𧻓�bX��"{ei�=����7�[�BG�_C�I�D�|�;���s�N�*zx���)aB|����# �˖��r�-'�|:�XP�1��LUՉ�I��"�k���~�
$�T��Z�Lًo��O�V�_�§?��.�Iʺ��p���#3�� �j6�v��ӈ��\V
��]��V��R�4�0�V���,��ʕSV9-���;�b���:9�R�4ݜ��� � hi�$��(�~��O�u�Y�.��n4�o�����7�aÆ���8���>u� tU����E�|;I{b݌�O����o}���x�O~֎�.Y�b��r�z�>'�����f�v�[���zU7x�|�W�����o���x�>��Ο�韂����~᪫�2M��v�����g?��?��k���sE���U���Z�9XssFXD�9�"��S�m	?8� G�Ai�lX��D8I�_].��(�W���Ë\A�)��g�Ɯ\�y�5�i��NX�yD5bۅ��E�DZ��e'A0s����;�ĮDI2�.d�e��
�ȡ�DL�K��M�t���l���"�H��܆*qyK�kq��"~1�;���K���G���N��$�$!\�,6�\']WG�^ ����Gm-ctq�ҥ�V�򜧄���2d�>��j4�8Π�Э.cej/]�]�S$ӄC���X�D��l�g�L��� vg�/x�>�6�X���9���@���``��s��L,"��ߤ����FT����(����xf��j�1Mv�����|�	#Y��E�E՛���U=˅K|��*@߼Z��/+Ǐ/'<WI�<�0����?�h4�#\� ��?�4�m�<����K7����;m��k�j;D��Bޱc`-t��-�~���
{��3�� p�V�NJ��<33�m�6���h�]���m����#�af�R��*��(-F���vP��|����������[�����j*��pg����d�*TW@�EZe���5���?"����f�F��9�(t�2��m��g�1����B޿XW���i���!A�_C����ͅ*��c�^09��X83�#aR`!QZl:T��t2ݴiS��~(�v���`G2���#[�N�H�������F�k=�ǖ�R�6���/��f_!٘���<�c\>r:J�i�����2
�2�D���T��ň�%R8�W�T�k��@*�|>�}�K===�9���kE
�֖r�`��d�,�+K��S�D�&q 9��)�D���$\@Q/��u��D9���gj�A��1d)�(i�9�y,��"Sp/s
`ը@!�Օ��m���4J�9Ce��R%]J�*��`�R�pV-����,x��<�aB�Uj"�)�Ls)�J"<���(�0%���+q���H"����D&+R����֐��YB>���g�yn������7�HC�v��u�	'���<�����\T1�@���?��w��#�ra�O|�������7�y�qo@Y�%�!�M�����?~��W�\����◈�������׾��/~qŲ�w��]LN8>>N>B*�����ۿ��}���?~gp�k	}��4L�oSo�$G��A�AqVY�\����y����볰U�b��:BJ9Ka��u�j�!��g(Գ.F�O%ODyO���JIDAy�%��i��暋/��b���z2K�,��]����Ǳ�+��$��~S7�+�/��W����mw�}w�VŬ�4e�] I�
��O�&����Go���_��ᣍ7^z�/���@?�� ŷz��O}�S�} z��O���O�|�� 	��{%)���~��`���u��*���Q�K
!��$�gL���0D�j"T�?_ �i@��g��a
�B2�;[��3�O��|���͏�5+:�������>~U�)����������b	L�}FҪ�3B	I��U0_���ikHHe$)�%�����h�F��$�=���;���'��H��P$��)�B_��Ɗ����{>�#_�tJR��+�A�d|xJ:��㊘0���h �qJh�e7��L��Q��kŪU�b��:�v�{[N�����+����0�B7X6��E��h 55�trژ׊�6Q<P�?4��P'���ؠ���S{tKu]'��^ %���}�� ��ǖ(��n6lߓ����ЕI�`�U�B�t !�h;Ǳq�c�T�Z&إ{�l��'R;�f�=��0j�眅&�+'z{�#�>��(�B��1dGM�Ew����2Z`JG���ģ0s��ʕ��TuժU���޽;��)�t����L�XE�@�Z���V/���0�-W�`��;k;R��ڮ�R<���+��b�ϯ6�-��j6��MU��k9�����&��'����-��0_����}�Y B���"<'����
���Ő�3ZHƶ�{�zm�L�>�Į]�򴃖��`�d��WS�P]1VV��&''�v���W)u�z�o��`�휛�駟{v�3ϼP(��ט�� ����C-��u3�5�D=7�tUf����8h�)I"	�� �Ѱ,��;�˯�̠�]����Q�2�8e�J�g45��Q�-��z^�f�k�`�ZV�I�� .�JBw��_�>Ț�S\t�r-5�%�{
�T� K[���06n� b	��` `DHFQ";�-cߋ?҉�]�p�b)�����I��eP������C�I�\Q�5���ry��m{��f~���R���_��� �S���)��V`m�M����v��'��p�a�o|�9�gk���,W�0�;3m�A�v�ݲF���G�����ӏ&����;w�Kk��p�5�k��|�*�uC�rU�a-kϞ=n�<g�:�2d�t�B��X�����96q�&���R
ژۦg�T\�r�ZA�m4�'�!�z�����r�����=,�%�h1��zOF���'�d(˞�H��Fjƍ#6N�I̴/� �bpǖbݲ���׫�
j1�+AU�^�ױp�k��m�;]Aʨ�m���wq� s���Æ��׮�j���!�v@�eDξ����Nmin4���u��7�q-����@E̥)�f�(+F�Kn�D��r�;MϷ��1s*���%#�����V��*;ꓦ{��U�t��0�T?D�� vS���D�c��B�%
U"LX	$$�EN���bJQ��'f�q��H�r��DG�"-
��/�T�o}�>������f�*�|hdv���z���M���p�q��)_�|� {It�d�_��ݱw�M��Yu���N�0��䖢�Y��uI�E���y�ah�
�{H"�)�0B���/�\y �]��>��S�C� Ö�Y���ܩ��^��ǟt�o��wl}��!wK��Ӂ�� KQ~q�\J�RE��ճ]љ(R�M��]�$7�i��_�^� �1�&�]����z2X-`ebP��Ϯ�~~b�s���Yo{��������+~��]����V�9*���C�]SʻuXEe/��МQ��sܑ�?��}q�)�*X3���+y�Z���[��9��/��e��E
݊]��fNoٍ�KK����{�]������d�{�{r3"���Ș�Y*׭[w����fC�I�l����p�+� �A;d��ױ֫R�ڱ;���R�z�b����:C��/�&��"�RG���������^��4&:w��a-�T%��O�2�8X@t�����A�Ógd��E��y?�(�6s=�{����D�g��`��͉��,�[b
8������2�;v�v�m7n<��Sg�g�
��?�����!�)u���M�l��/�ݱ}`��I�B��v��3��<��×�|���y�իW��́M����{��wYLrXX�s��jzz�d�dn��]�q�J~�$�����y.����.���*�d(�Nd���B�+�0���Ѣ0�š~��s���H�b�}�w;��ݟ��' �1��� ��	x`�#k������}sib�Z�܃�0} ��\�M��?�
�\����hضE���%���y����}Y��3��jCO�9-�,�c��`pK���čB'H,���5�Fn߾}���c5d�oٲea��b�޽��N;m͚5��-Vo�z�P(=��w>�8�ߵ�H��ѣ��o>D�t�\>���GF�����_���oD_)QqE�"
���T�	Y�K0������ ��ƺ8�0!ˋ=�<���NPj�����1�!�N/T�$ػ��-DDƼ�����j�p�a�*D�OS�M��z��������&n="6���QZ��I�q�V3�'ƬbR��X�a�#���\��#"l!SB�L��q0=8<B=���Y/����S��׳��2s��x�?x���剉0Ac�G�����;��aj��-[��9؞9
�z�mذ��<t�]w��M�U�8x.��Y�=��3���}�M�� 1��>�mj�nx�a�Q}�d�b� +֛��oZ��.Q,Υ��-ղ5cM9�#�[�nw�g��=��2���;B�ɽ�n��Z�5��`�K��6V6Vl;��L�db�/����XK��(u�H�E�TU���ڤ,�+��R��8CߏDˡ�o��|9�y���kƤ^|X2�n��@������ڽ{����{-���`d���(�J],�`ǲ�6B'���Mϡ�!������Bce*��A066��GЁ����z��n7�.�lv�֎���6��3C�ɹx�������r��ތ�O"�K�,_w�up{���g����>�"�-&�X��}�c�N��\��]s�hQ%����[�+��6V�N|����k���UW}�Ot�	�ș k��`�>���_��+���o}�Wa���}��^!Wx������׾Fx5�H��)�_�;�_��l&u�x�i%6�-��T>��� ��gd�������<�<��p� l�TI� �1�}�o~�ǐ�,Lv"/u?�c�	SJ$��	<�� 5"�ա��Y_[VBJ�\��p�'�|rww�SO=�m8N�0c�X(s�8:����;묳`IS���x����:�\���ױ֫	x8h#i�})����2c*��o-�R�(JD�����Π�H�V����o{tn?�	�`��~�j
'��>I�_�Bq�HiqV$�����l8�����I�U�l�������*��4��!�8�l3ޕI*$`4�0���FZ�Pu�������o�������B7���P�Eު��e\0V7���|�V�����M���m�����v��:O=�l��U�r'�x�\kF7��������ׁ�9d�Η�Q�ޜ�oy�\ox�+B5�O�l�,fCN��O����Q.��
&@�l՗�)v�ڒ�.*� �{aI�=a�
��Q�-����Q��ЏR�	-�@��e�*E?0���Z�U�J��l���m�WtTJE5�/�D��d���\�b1�/����%0i��L$W���D^Z8�p�l��`dc[4dA��Q��s��F�i��Wpp쀸�$�~�@-M�3
y�EdP��iY�j�Y�v`�@��)��.̈́q�Vmv6��3Z�@�P��px�>mI�hŶR�LŊ��4Y�꩔�J�ő's�d	+7�4'f�D�?��{f
���X�400 V�ҥKO9�@0��7od�Am�Î��	����T�s�Bx:L-�,8	�L��U�kD�C0��BO'B�̳#��i��Mn�'}2Dԃ%�)FD�i �92'1�.f艐�Do��&�Q�bJH&�%b)4�ѥQJ��GfK�>�!+6nz��}� Ɇ�˙=����܃����r�D�3�����(D3�	�,[!Z��Ц���"z9�w������;�K�c�	�*���k���ҕ=� E�z0�����ON�ر��;n����V�s�p�^�2;;����o fs���L���s�������+]J�ɊI,EȅE�62�R,c����D��F�c��V�4{�#��	Q��\�G��b�4j��]�5;�U�g�1�q`V�\��i�^��j���!w�nad���ZG���h%pR���1���u5�0;RcȚ�; 2e,��Q}`�v��Һ�� �F}�b
 z�>z����R�)�!���d�*�J]	�p~��f)�u� �ǧ�&z���}����}�.�x2�i� �X�zhdhzvndt���C=T�ٺ�W�Yհ�]�>x�Z����d�n��-��9�m�aۡZ �q��[�,� �
�R�s��z�,bU�XQA�"�+�	��R|�_��-�M� ��T[��_<�/�''�/�q5W����ͷ�����7%UC��ț��O9������30%tCSU�4u�����x8��m���M;�sց�Zd�B���{ʛ�>+ [DՄ�t���������ۻ���͏9���~C� � ��_������NXO�dS$U��kq��_��>����i�u�s崱
'��b-z�/�#���� ��Ǿ�����'7���t�h�$��CXϊ��B�&�yU��b�8�� ���H��p]+W��>������o�h��0�*�!�xj�ŀ�]ۺ�	U��._b�Q��+%썆�:l��-�����qǱ�R���N�!�V����gϮ/��(:*Q�5I�$q}h�� q�3�ױ֫I���0/��3�4��@<>��	1xG�'ۮ���M��y�3�$^qQFԏ�*BEKjfԎF{�i���頠V�c���^�W
����<���G蔶Q��'��o|����� 	���Hw�}7�5�W]|��3�GuT�>gsm,��� �s��n¢;�,X�%c�4Oh�P�={��.����mpY�a��ny��F+4��-�����g�ynbb�6(\#QLww7Jiߟ��D�g��a�V��ը�$�ɓ�4p?�� zt�6/*��K2.W)���ի�y�)�)(���P�z�L�l&b���9c��z+�4g��;66'y�'6^�n�9vO>�䑕C˗//U�p2LP*0�x�1Vˀ�����6m*�27����F�}���[�@0#۶m;�#���7�38҂�(�$�]vي5k�<-?�������>����'٪�Y�&o��� ��v?��ꫯ�n{]�>8���������o`���c�>�G�nc��g���-7�8�!�Հ�se$=���w���7�r:"����n��W����C�������`Ä��<.R4�eٱ� ����a��g�$�l�!>�J�p�a��� 3����OvA�иȉ�1�`������N�s�d�&�W�>���f`0:�J��x.����P�\L��0`�%7g��8�&���u���+�llӆK{G�d26&��r��*>�*af�C�vp'L�(Q	;�Er���v/d��C@���6�$)�a���&x�o߾�}�{�z۶p�\olE�T��b�z��~�n����=�\�p��N5���sOD]V�\y�1�L��+G�֨
�
�{ (���8')��۞��v��ӊ򤈙�q��$����M��
75�$21#�*���X�Ѭ��ԏ���������t�ҢP�r�*'�JT���m����S�3�u��k'��<ؗG�>N�/i=P�At�����z�n��P!�>�'�i�r��H3݄�XNzd�T�G�a����b7^H �F������<ʢK/��N8 ��t�a�	.�,�������l�QaF8�)9�h�?�裓���<��UG��پe.'��U�*��v<\���_���h���Q�#�M66i��^�P�Z�^6��$��nQ_g��C��o~ȋ�����d5��緱����֢ y,�
���=�\�ƞ8�D�A���}쮻�:��`;����b0 �22�0t�,A�K��%|��0z0,�"9~X�� 3�1������A���_�L5�1�J?�s^�t�%��o~b�q�-�.��EI��R���0��@2�pM�� v=���_���蛆��$ղ�>�����p��8��W"^�=���ᬥR��(h~��T2��`��#�<Z��t��@����}�j��������z�'D��,i��{�?����� �iT����{�6��X�U�t�f�����;Q�BR����3y�	!S��3��s�#�M /D����.�j�_B�bZ�(����$A��Wi+=���M|?"��,�T�����Ҳ���Y1�_�f^�q�0"��H�"�ΩB�+�O�7/\�0I��׽o;�U> �d5��Rt��n�w���푫VK"�O���5;;���=���۶���Ī�v<�H�Y�)�|�q#�ԗ�O���󁇋��3�8c��嫏Z
���m{���{ם���8>995=m�}�X}�/��0�l�2$�0��7�:4�dfA�-�B�X�t�-X���ҍ���k��*�g�ǳ4��eVD����}��XD���B��Y��}���[X�_o,4����<|�J�W�*C�вѨy��z=��a;��Y1R���(���k��V��	����z�n{���-$ߊ�n�~ 3���F��]kh��](��w�oU1I
jxp�X,���l���,=_X�f5�v�dbc(fMWA+#M7�B�BP_D�zU/�F�����'v�N��c��mj��K�,�q`<E�QU��T-��57�ʠ���ڧ�/�+�ݳ��h03�����[`0��GL�	�G�n	�Y��"|"P�`��0�X��T.<���`�H)����v�,T۠L��{@�66���D\"3��s�è3k�����)���i�2��(�?Im�W�l�`xoa��@�Ӫ�3�aE�:.���ZZI�dF,�`���l�	�t��+���LM���:b�sUaal��lAD�X����a:F����)���G�1L�j��k�����'����`�
d���i�Rt��o�0_Z�m}�y���b������,���"�����}D3=>5#3�d>ݫ<TR��&%�X����
;$��I5��}-��ꂲ�b)�E�ۍf��a'r�lV���\�=00�^�ț%vb�E�@$;����T0_]6<�՛���]�5��j{^!g�Z��Q���(.�M��u=�(�P�v�00p�D�a�`�܎(��2���8m�h�*R�ceV��[*9�as�F���v���*�S���9(�/���?�M�L� XdL>5#����j��c_����_)���/A�_� Y�E'&&Jf7X��n�w�}��Mo�9��%E���2Ct7hc�v���s[��r��G-���l�6o��o��զ��xvf~ll��g�v�/o����r
�<���+.�,E����k�z��Y6��ZI01�Z��n�!���a��`�e�䘀�F�%'%�/i?Hl���R<DD�X´]�(�,~�g��*�������k���+����56�%�y��+ZN��+����h9-nJ��\��e笏��H�a�t�SL�4����lݻl�ZU�7�����(�tLiVЪ�o+�|ҩo���[a����a����?v�-��q����}�4�$O������z�e��ʏ�i�eGF�ƽ��t��`�с��sE�"):܅f�:V�SN?��_�jzn�(+��ANHX�J��8	�H�G*����rjNk���i|%V`�Œ|�I'�y��0"r �*aNF�I�q�rތL���׀]Ѷ=��AD=ăw���M�ܛ�[۰acWd��b%�8��������/����tJ�MYZ�ȍ���6����c����%$��4�,��EP[�N��Hخ���&�o��/�ӗ,u����A���'�Z)3�{�#d�)^���8�����.ޠ�o���#~#��� �dN�͉�d$-6�b�-0y�}��d9v�����f��������1��ntMۥQ�\#�:��y0��؟��ch�����XAD~ba��������]꣏>j���,T�Ɏ�{�}�AӶ�@f�sH9dr��M\����q 2@��9�;��7m�422�����Z�vնm���p�o�`�/[���IH>WǶ�fi���rh��&Ze7a�j�S��6����t�Mp���N�����w��X���`��A3;V�X��}�T
Oq�6���刃��XJ�X��U;����ov�&F#S��cǎ����Î:�Cx�E������[�������O\��+.	�}���)�J�+V`�G@����'��ٖ�wq{4���@�J�p��/�x
�pԱ#Q�{�����g���N8�5G�>��v��{��W���)O������5� 0a$W�Zۗ#9x ���F��sfV�a�ا�Y^�����.�Ѽ�S�H%�_�ԏ�Q:����1�TT&�U�.�Ѧ��+r�Ac�6��I8����U̸�8͏}眽Ü�܆@<�v`�D)G-J1���` �PƷD�ɬ�\�	g�� �2,8�����f�i��T?��s�t&�?=9-ww���t)�C�lCԧ~��_��4n�v�����uC���3�8C55�}�����?�K)Ӻ�C17���L��#�b?��R7���gRңa�<�Qߧ��� �|�Ow�<ꨣ�V�b�6w�°!�=�۷���={p��=;w���02T��#�1CE���s�E��p����=�o��'ӊhD�i��	�HE�6s?2�[@ͧS�C����� �`�G�*
[qr�"�rh�+2�p`vS(ֹ��&�?��B��}�477��C=��#'����.�U195����;@&H���y��k��?9O��S�EG�)����l1���{졇_��3�>���q,\��2���>��[_��w��m�ؕ�B\����#�Uy�a���},q0�10Z�]���T�'�-����/�*��":��m�w�v�D$�|։����ʀM�sh-S絊#���u�t<��n��[�W�(9�H�rͦ<]X� �R����b�¼�P����X��f��0��>H���������,S$Mڥ��xec�%�\~� Wĵ�T՜.��"�N�&��or|!q�*a�+V��'��x��`�]/Y��>���.����������n�61B��^ݿ^�����d�K�p=��\��p-�����W�?�<l�~�V�����E���w���{A����J�]�vć>�g_���}��_�b�{�S�̖�4q,>d��k�xk�Fs?H1U0s���{~�9�����<	eQTÓ�y4��1���?�Î3t��L�}�CS�0�ej��悒���8O�!'	cu����eI 3�R|�4���E�,^T^뾊NIG��e�4�`'�{H3�����^���	ȃ�U����k+.h�v�V4}�Vw(���B����53 ��c樦��B*r�%!L�����E�D��3[:a��V�m�m���1]�M�}ɒ��-�8$��h`�&64�R�==`'��F����r��2��7^�n}MѶ<��.��9�t���s�r �*�����tݩF�V�%f����k�9P@�� ��=��C���}������3�6� ���#�J�#/���d��.��.���n� ��0i�2���*��&�c�Y�Yϩf�������և�D���Xܒ��� ]����=��bvVq��a�`��ص�fc�ad��]�;��_��A&u�$ka��q^�"�n�O�֯Y��K";��}� l?�i�����X_́�h�o�A�\"���>I�Q޶V�����N+ey�Ms�ڣ�zꩭ/�:03��R�r�R�8�`������Ё�^��jTQ������� t ٺ�M-��v�[�1��Ku���!�R��@AN�e4������(�(`���$+��ɺ��r~,�� �� L��4�d֪D�ܡ���I�,�me�Daڄ0�t��8VWF13@�����3̉�	���UkW35����2�:Ǹ������N����Y�x0����ڳ#�/��ǿ.��}� � ����wnG�6ې��a>���`Iz�l�3�>M.��JE1����'@��ڵk�޽��?��/_:������9�Lٵ̼��*�p.��D�1�%��VM�,"䌖�"� �+u��,YQ��}宠�jA�1��ؽ���2&R.��p��]?���)+z3G/]	;ezrzf/��Z��97�m���=Rt��Z�pK�|����K��"��ak��#~����4=�[��n@�K��O	�!��i$��$G�М� �@�"0�2XYz�:k{
�~�
6�b�y����haA��X񒚓"ō��Gx��S[߼cx媍7�=�DX�-avn��>04�>�gr��y*�sӐsfW˷���¬�HBC7E��lfO��^ط{����r�e���v����N+z��q�/��ѡ�%Ł�cc��i�y]ɧ}�ecb�1B-)���^��}aS)IE� h�D>��X��o���)�h�EZήR�c����e�`�<�鹣�=�$<��%�~�{��>�:>o�=qꩧ �M�kϩ����w��O�~��p�ΰq�K"�TY��X��t�����lJ��۾e�ް!@;�������eU��u�ɇ��ˡya���{���7ޔ3Ko<�,��"�2����:5))s��"��ό��O�"RJ+Hi UL1���!%	�pK�|Ix�ׂ�i"�E�\���`����V�����
���OV5س�@�e�v�uX�`�Z��f+4���3]��'P�*�n�hF�l{�_�R���0VU+�·]��w�~�m?�y�Ֆ9 yM��1��P���{���W�_)��Q�֭W}�}�������mo{��v�y�&�h�-�(�`ƈK�d�/���?�xk�ʑy����κ,qP�����~G�9�t��G'F�_1����Q-:���pvRF4zً��\��#N1�x5��B$f���^�;�k��\���}���ؕ��ㄅ�~��P@�`�
��r��ϫX&`�fB���c�2�1{�����1��N曶,�݁�Z��T����f�����hmn`�+S�vUALe�y�ndR�C�w�l1���AI����&�i�������?��?�p�聇����FFF�:�.M�f\��L���53�����w9����y��e !�\g�qF����m�����$r�)S#$-A4�-i�1ziӣ�28 K�wua���f� ���w����ۍ%.8N�+|4�̶����;�ԽqBӇ��8���F�:�>U�I-+W���F��ޞ#�<�9�ؼy���$�.��;���(+��k`5��K�η��8p��37����� l2& Ｎd��x��Ć�����ᇫV�ڶ�&�G�>��\���+�r\��A>��,�Β��O=>
>��҆Hg�KI�+g��Tr�T���GHU<�e&ՠv�RR�E���2�
;8ږ��ӄ���\��>���X�
�T�2�0�6���f�)F��OnX��(�o�=ĐBI2-9��|�'�k;v�عsg�YC@H�}:N�X�#;U�pab�n��=�⦛4C��;�/_���@N�a�
�)O)�O�T!f0�Y'܉ʋ�\�.Y%�U�V�qh��900�kzv"<�1�gX!{��Р�S#Ῥ����,���]��lE���bxx��Wn�^OqĊ�
�(+���J8A��$�a�	W��:	/X���������,jx���#R��h��+aU�����z�d�7�f�����1�)]E|�ꫯ�3�[wT�R��g�հu�����%%s�s#��I�� C���O#!R>��W������V��F�"ׇ����O����������mGh�W�E�m�bE�'UT��c�N��[�9Fh��\���/�q��j�N�Y8֬Y��;�<��Ӱ�CN����!II���)�A���������t%��q�{�oY�˾]Y�R�ߡL�v���W�����ׯ_3����4V�����>�+���B���'h�Z�v�����-1�����<�/e�@{9�
Gv��}��a-1sl6��ˤ�0 wJK��8	:�%�\�W_��_�o���xyz$bAɩ`�2��(�〮l4���[N�lT|'���P�zm�1�� xq
���������W��s�=��c7���b���{Ϟ���L8�IڪP>��O�ߺ��^p�
&a#`����P|b9�;���?^�Z�rȂ7(��1��J
� D�Ɔ.��|B
ZJ��B��fS�9��B��'�R��[�`�E�b��!�K�^"�X��;h�,��k"��^Ĥ����Qd�T���"�|{�c^�6d�P/r�ai��a_HjR�Eq+ΛG�Jz-LU-�I�Ȃ����A�����I�N�{�v;�Vi��� ��3v�8�!��<ʡ:lɴr<�m��qԨ!�+i���w䀹{�%#�5Vk!c�ft�0����YTT��C��nQ@��uS��Qġ�;��R��U�W0���PU�v[ ���d����Z�Vl#�[d�R.o�9�o����A��
Z^�u@�k���P���Ҟ�����AM]@�]1�'�]�v��Iv�A���%��L�5�F�&i�+`�Q} G��ʳ��md��� ��̑k�ڨ.4@j?�g�
eE��h i��nń�� 	�����DNKS��Iwnfz|||�尀�b��Ʊ��4�Z+��<�Z��k��=LMO���bO�����j�L(ϛ��.[��(D���ؖ���%����O]5:�grrjn��I�ԓe�Z����s�oݲ��@���{��`���uj���y���D-��z�Y�(��*�q����޿e�#�<��o~�97@��2�\���B�vZ	�;�yd�/���Fw��^�U�>������0N�׫��#����"u0̸c��(�I�ݡ��6CVZ�'L��c�8#� l��
:!�ef�v��G���N�Ґ�k����h����l��=pU�����l\6Ñ+�ʮ������߿�������8l[j�R�c��0��MĨ���|F_b���F��>d�@Y��sOEG�z��x�1pŁ�Q8[��N�*��	�:�|�e�^4������o�
���{�0b���w~�-U��>�1� 1Fo���aT���X2�韱:l]�zlo)��.�!
:S7Ɩ��6{m�H<3t�+�Ǝ8�TX������I]5w�ܫְτ+�/�a�n�t1��YXl%	aO���o<Z�Y===��Zm�
�ʋ|�^�W�{����nV5�d&L���R�i9�Gi!�,��{35]�Ia�"k� �-��Vo4%Jy����ڱ���r��@$`����^d"�g�����0NH3	S�x��2s:�w������U����z}�����уV,�t��1b/o�9�ˤ-�
� ������h7��\���j[r�J�0j����у�F�oە�f~U.�@��Af��V�����}ꤩ�)��!�r��셪eY�*2�������}6�i'c#�D�%�i/U���n�"��Ҧ�Ⱥ�@�������K����o�fŪ��������iXtJ�%ƍb���O`�*�X��P�-l7b���I���*�gC=��B	;�Q�ػ�}�_�է�����y��GoP1�P�UЧ��������D�*^�+u��D�p�=�5[��������!3��GC)�X���$b���q��4#�|��]ax(�r��6�I�a�w���5K8"wj��Ϙx ��	��p��*���c���_�9��s��}�����>xDq{�t�u����>��*+؆AS�(���`�N�^�@3�(�)E��`�B��k_m��`ĚY���;��7���7�}�[���`wŋ�O}�S����p?����*ݽA��C^Ϳ|��_��뮅��ʶ}J�6y���0�"Y_q�e^�xMdK���^�$�pG=-�VV�
Nr3]d���TESM���Y%�&��6`��(��˪�y�b`6�}��x��b?�����N� 7���S)�vB�쐒��}�%�t�fJn�R���zq�����!�F��ر[\�y���|�=��v���f:I`J���B	l���׿~�����������e���0<aeT$���M�@�W����x�92�J�.�QH��������lZ۰v��ÏY����{M꽃�Y``�R�Ḁ>`0W��٣�NVA�M|c˦���ĳN6%�)��z�|e`岷	u_)`a�ɪ�Z����iQ�9�S�#�M���ls�1'�x⪑��V5؎���$�a��U���4oc��ӧzy�M)2��m7��S�8r�u*��Ι+� � y�e�*�o�Jd��ԈI��5�[�&��@�5�m��?���Ҙ�T��*�4"Wo5)��z�y�'$�/� �3��s�=wź#�����bŊ���F�ǋ����f\7=7[*���S0	~��5uy���t��$
�pٲeM�>��ұ�;�`���1G�ݻwU���B�x��g�����<��&����4�8�����,�s3I<uww���>Kt�:w�r#�	���c� �1[�r~V�I�E�������1��Hr"M�μ� J�N���s�2���l�q���\�����S�� .���/ު�{��v��q���-��&���x� Wf�e���Wy]����+����e�����D��\���G3&��^���?\����s�i��E��o�=�Oc���A�Ȉ���LLM�%BY ���衇�%���,n�~q�/e�ɛ��!�1٭Ɵb����&Ж�չ��fw���TCAQ ���t�hƀ���Db��8��y5%������&j�6��D�b�A�AK��h
��NS�?gw�_��oνw����{�x#d��d�9k��������ɭ�i*�)�]q���~�����V�F�,�� />�+���&�V`�"^H�I�;a�����ʕ+�-�^p5�EOq �%k"|Y��\JV7-Q���I�<���y�Ix�&��N��G�ett�V7���ݎ�;<<<8<DgN�L�}Q�EN<~��g_B
���r9/��r)�4gՖqWn��i�ilM��m��M��Ϧ9�gۤ��m����~��U�g"A疄�$��ñqYE��KN���3^���$1(+��v���f��?q��N:�����O�i�Lu~b��Ɗ���)TF��F�0M1���khV��ǰ�5�靠�rmw��;63EӖ0w2~�^f1������o~�I����i6�H!��N;m��T�%Z��ы䰱m��(I=W+����v�g-�IČ0��x�����?�տ��o|㟱ڹ�������/:���ZWY���sH�G}��Ib�.ҋ.%.Dd��5w��i'�bR2��%�(ٞ�Z����a��O��S�lL�i�E�\D-���YZ��'Z�?��m��T�e/��m���/{�$���f�<c�.}��}�{�oR�e�l�!B�엥l�kh�j�8����9�K�{�_�ӟn;����b�&���,���>v�WB:�Rc�o����w��-ג�O�ai�.��]�v������ֳ���$�,�H�"s#cn��_t��}����͛O����m3�<�F颮R���oXyp
��p�x�o���1�v��)=ղ�G�W��L��僜PtKre��qԥz6[/�Eb�d��ޞ�&�!�f�e�<>���娎�dm���;}졇$�s˭?<���J��2;�SW�k&a86q𵯻J�h�D(?�K+:�4{�;a;<���s��&�v4򱯯w蒾�"7���qfhëV]��7�����أ�{^�w����&�I���S���X�u/βj�n-,�D7�,32�e���QY���B�EW�����&�	�H͒_�u�P�`;V��m��V\�2�l��h�Q���)��_I�%�GR��{%��g��y��`����Q��͙������ӷ�M�Yh�i�\r�e_��W���7�s�9� K��ܩF�D��Wl�ou���y����k����L�Ɩ	��tf�� s�֗����.�}٭N�Z9�fvi!��5���5��7iӰ�BCK`5�R1-9ˎ=���Jz�jٞ6�&�g�Y�鞅҈:/����2H�:)���� �c�4&'d76�z�	{)H��yxG�/%��e�-�׮]���>�xp��ݳ05i�s@�ͤQ�*u�j�t��	���7��Ҫ�0a@�n�d�L�^l��*�qd�����"��X�{�� ��=|:�k��4-�-'n^�b�k�'�x�y�_@�C�>q�m�m`��A�EY��Duqaan�������Q�X�R��=p~����7�+�~�F����G#�e尬�k�o���;5�]��_�$��L�<�sP�r��KHt!X���M���f��R�8M.n����bY�ͱ����G���N��אX���2�\�,����&�!�ѹ"<��d�q��ТM�8�q?��A|�4�Q�^뫴�W��/|��������I���_��w�^B҄���ŏ�u�g���졾4ʭ���ىɥF��=�q���~�}�Y/h��|�"�x<�ڈ����t��5E�>��41�,�s��;n�d9c	D�eZ}e�'l�<x�`34,W�_m��Ǧ'��$bO�kߡ1H��u����!ں{�&Ч.P���Je���b�ު�&:D�e@�$K���j�$�~�"$(�ڶW}�矰�d�p���h�]'�x��_�G3رc���C{�U֭�����S��׿�ܾ�ʊ�7��Wќ���~��;��(9�]xѫ^�*����ħ?C/���#lZ�=��F�f�xe�^�i��L�0�0ր�L�4uI��7rN��+}C�zW�"	f�e�8��Z�t������^�Մ�-#)�\��T�X���<�R'�k��|��6�V�������ͥ��P��+.��3�8餓��v'�Q;T�^��7���?�Ѓ$�o����N;�͛�n�J�����z��d
Uk��z��7?��n[ `ٺ����s�T�/�������wв8�0�)8�I��WP�u��m��z�%�?�}�@� �JH�[�Pi=��C���?�G� q�E�U�#C#���Y�VS�i�k&i��2d�q$��[��z�w.��U7��7�o�Ҽ� *��P>��?z�տI�+�@*IVv�\�I��~�$H�F�Ė�/{:�</�`-����=��i�� ��b�HH��2?��L{�Gp�ѻU!E7PN��HЬ�V�J�	�	��Jǳ�k��BC�V���a����P�����<��]?z�e��Ц�=3��#�ȟ��%�"d6�l�/��/�Ȳ�'hP�鎙)�n�q�d-�dI0��[�����s^tv�%���Ч>�)w(��7~���=$R,�>�����r	�x�����9��`�:�밸>�syHP=W��m�g;8.dt��࿡M��#�LNNҿ?����~������>�<�z=�7
C������oذ�d�oH*<�~i����n+�1�z2N���� ���{H[q��u��˟�������,\tY׻Dp�xG���h�Z���gH��5����?��?��ʕ�A+�(��� �%�����k���D^ȟ�PGO�4�f���=�sA�`�48�4�,72����$\r-�]�ܳ�:�Gw��Y�BHw�������C��fgg�ng4����-�ۀp��pu�����^�s�{IP�o� ��0�;-�W9�fH��^
�¬����TШ�;g'3��@�
��~p�Ey"1������g���.%=t2�n���)=ݸꪫ�x�[nQ�2g��8�ѱY{�Z��G.4���љ;w�\�b��_N���A��ƶr%ri4He��}��1��c�)��<��	4#�'�ws��j�Z���d� }(E#i�p���\_w;x���>�l���m���SvQI�rKc�N&;�V����f'��F�b�8.;??ϝazR�ɸ��f�]g	�O�֢Wo����b�-�	�u�����P��q�&�y�M5�~��f��P�TQK#o?G�[�4\�z��G�U��y�Ӂ����4���EzH�KʐX�p��q-m�/��e�c��n��Gt��-�I*#*m�F(�O���ډ�J�m�\Ј	[`Vtz%���$��(Vo<=ϔ��$�u����C�W�I;�6B"L}�]�x�ŝ�'5Z~|�}���|_��>aRZG� ����%�9������Z�el6��h��q��4ڵ�Ee�n�L��633F	�X�j��$_�fFzXͷ[��IK���Ǚ����k�Ak�N�s�@��\mX�E{��<K�r�9�̞-[�WJ�����=���$	A��yM�\,<zL,�R'��:5�9����z�^֒�4Y��X�8��s�J�[��V��_!=/]��VH6X��y�m��%��.Is��_��ι�կ9�3&&'��Y�~�y�G�4g��w�M0)Z�I([V�Dcr�c��"�䉡v�9<�d�c��5��Ø6���J���6�x�$NESMC�e�35�������I�����PtB(�O��z�t�Z���E�+���ٳ�~C�%}���D�@"����O�̡��c߾}�z7m�T����)���*^I�ދ�����C������=�-Z*�J�;myi�eQ�����e۶m�]zrؼ&������?�1�R� �h�iWΡ�� 8I������5x,�UOtnrP����ϳ������}�oI$�A�����}���K^}�u87��%n/U�ٝ$	?Բ�-��<���)Y�4c�G&�[�K��zf��Z��e�0��Y*F��d��o��e'Q�Rd���6�#�B®"S�[����,���a�'�c�9����ˮU%ű�\s͛���=��s�k�8�{���)-0�����E#)7����?��g�ݐ�/��
<��S���o�Z��k�_iZ$K�IS�5�e��X�����v<ok=ˑ�Zj��G�w�}���|˛�p��?>86�v�0��I��������V�}��?���G}3{�����������M���?���شL�.��o��nA��0z�_�Q��@ͺ���:��F$�de�����+p�_,+�*:<BG�<V����Ar�������^����ݛo��[o���v}�p�OZ��m�!Q�,��~�������ǧ�Cd���A?\�)7�:	��_>�6N~��~ָ��)�1c>&��M��pҦ'�49?K�ɭ�W�,4�߹����G֌�p҉��v�ر�8Ir� ��̜���U*����E�z�3���Y�*G�{�I]d��bŃH3�5B�Qcnv.��p6��v�s+W��Z�G+�՘�1a��`�Jb�I����>��v!�S#Y�Gs��U���/>�ԓ7�F'�CV�٧lY�W˂�Ё�諕se�P߰zm9)hO5���k�^kpt�Oe)r�J�uKq�Kw�� Y /իa��M�u�]���lc=t�g�r�Yʺ��S�Z���3H��Fj���]ͱ��F���=�H�Q3}�F�\ͮд�~�-�X�f�n�I�^7*O㰽�dJ����D'$�b�y�7���%���{������Z��uV;bJ�����@_Yo#O�>_G�SV����f0}p��	jF��}[��Y^x�BzU��#�&����Q�_p��/�|Y_n��઱It>��?��*X%��Ι�%�]���ȆV$�֜�ʥ�e��z}q���i�0�p"9�(�M��$�1��̍��gh˓�W�Hcf��HM3D�@���{Tj���<�Z����4�d;��g�,�c[E7y�I܅�ƄtC������������4���bS�����(�RVx\'#a�J�ʖ�#4$��A���+%�{k�H��ŞGOD&�����L�����622�q�Z�����7��Dv���j���s���"TG�w
O\�`d�5��jSK�<I��-m�L2�mǵ��s��C�NO��5ݼ���>8%�zыb����vFBɞ'�W������~2rj�O���W]~��G������;E��?��Ƀd����o�޽���/�+e$��ư�ʀ\u�Z�0O�O��ji�iEYẾ�Wi%��'����?Z�y����Co|����q'm�K_���F�������Z��֞����s�:��g?97W?�����}�|�U4�̱�à��ln���A<�k�hl6\"f�|	bh첤'���fK�XXX2̔�6 wI���P�Q;��r�+����$b�iA�Zd�-�"��Gͬ\F���e��Y􂂨M�n��`��]T�"�!#X�Y�Q�4ڍO=�qӆ��V*%����}��k?�o/zc��缐���V�����^t��M�y���ʡ�#�yŏ���3�r���-�(��e�l��k�� �eN`�䘳<L&
{.�肔{�$��=?�B���\��$�RpFj�鷮y�[�MJFL_ncm:	��0{������g\��U�j�Ks���V+�ħ>�ן�+�`�f�[�)�tM� �4��?��؁�D��F�6�.؉��,����u���CuͰ^uV�ԪW�-K�H��RZ6���.7L���'C�n�o��3�)�2za$��85���Qf~�8�]ׂ��ʭ�0)z�LKv� o�QEL*��tHPA�2ok�!��d�rY%<�d/Y���l������� �˶���*5��]؎�j���0��r�{ݡ��hxF��~�>Q(yW>#f�e�����Z�r�BGU2��������7o�LR�����~��׿�5�^N�,\�#�F}����^��r��7����N߶m�^�Άi�FI���������TF��-ыn��$�;�L񇉓U����{��b}9�uė��Ng�g��N)B��m������׿���]v����_��_^{�a����D	�J��I���~��?���oܸQ�/�U��&�m�$���s��eQ/ǑJ/�u�й�3��ҭ#4���@Ӳw�^�)�$53=~��AUĄ�I�q���}�&�����s�VmYZ��%�(d�Y����=�'�y?\�	�ܤ��,�Հ�;���W\q��|��G�A8�89B?(Os�A�K�7�^4>贻�둇w>;��������K�/�Z�\sM�r���־q��ʹPRRe��H,n�vi,5P1RB ʳ���}�v���S;��]{��!C�U6l	�/�t��v&��|���S�
:k�;�":A��U�~ެ%��<��T��@�r��=į�&-�AdD��Wh��Mc��*2��F���Bq��E�_ZB������ХY�@��2ka -5'p�
کq숳M��Yd�5uE��7s�'�6����X�쬥���W��K.Y��sϞo�1HЉ(
�P$�B�Q�GF�{ݨPRlZ;ҍ��ȡY5�S�-^�^����ñ�e��ݱ|Sh�˭�އ���?{Y7`�ST��LL,��aۮ��1K�)����$R�H��׏ݭ�]t�s
.�-�<7�GZ�����d�NO���/I���$�@���0M�_�k�B��G�,Q�b��M��+/z�x���ϥ�~���Pʑ�iN���{��q:g�q�-�~֙���)
�[+��jVP�Jດ�;;3%�o� �9�ny�b]��(͐�o�<t��СC���o9������d�G��R+����۶�x�/���[�~�3�@]Q*��
Ґ3�뱢[��#0�PA�@���������N�.�o�#����Ϋ��$_�ȓ<Cg�����R�J�-��#�%l�ib%��D]�D}qvv����I��1]!�޴���O?�*;����$%LO�v���8~=NW�ӑ�躴=Q�$$�]�B�Cر�%��.{F��+N1�����N����|GX���SSS��Ⱦ��F����<�[Ew1Ъ!Yl5��0A�˷��''ѳk'�T�Ɖ� 'M׵c�#OH��r	��骳�c��E��g6!���2<�hcU#c��`H��ӈB�qi�����]ξ�\�'�2�!
%��,1Σ��4.���R��4���K,�v.��̾A0�$����l
̡�o\�1�îh)Q��*���
��'rC��zQ/i��k���P�GCK ��C�G^�HiY�rB' �*I�S�a���P	H�%���ê˵H��g�MMf'R\
�a��̕��T%h�Ũ3����z���&3
 	�k���hH�j�ٕ�E�p�8%�l�@���$Kx���β#
k{R�(���j��m�g=$l�F
w[FZ�{7�2qp��󞗽�2�q>���^��+&+��ܷ��eR�"��ҢlW;ﬓn���$k�v�8��ǽo/�I6���{��=&+I~�BQN���#K�(���*�k�)��:ܸ���{��+Ź�8	$� Y���Xf���|�帿��W�㷾��m�^���,-;Z���ꫯ~��/y������Xq��4
e��f"C����O:���G��xÖ�`�dB=`�1�V��d������r�R�:�j%h�H��Q�5;�0n;��[��^9�Y�UJ}h2�P��j�Q�.��� ��';4Q	�N�!4N.TZ��-鯔#��~}	�V��AF��� ��p�U��ڰi��iⲍ��2��q�'�O�z3
��"��4�J�`���ٱ��C�f���O>9YZZ������\���_4��9�)���q��)����]����X�
��;a�V���0@*K��Z����<�u�t����hI�qJ ��;pIu�NZ�z�y�;if'Y%6�4?�P�Rr,�6CB���9�b�8��.Q;j���k�a�m��ܡ��P�Xo���Dv�`�w҉'(f�k���1d�n*a��"d 6����Z8�G ڞn62׈m3Vy�a�Y��ЊZ������0�X+�d{���}2����b�O�G!�`T�a��}�}�׎��&���m�!K� ==H�a+񡂊����8��	�A]�9Q��jsM
����3��Ʉ�=�D������E!���ҩ�kt�4�� Ҫn�n�i���hT�=Y�D.��V E1@㗬WŸ�d�����[�C{��YEM�8�N\�t�гyJ�A���qp�D(W.�HQ�w�,��ubI�
�8XO3OV1��+V�~���-���B�;e�0]�p3t�2]ϯѨ�v�:a5�i֦��V�\$����(y���\[�]؟$l�.�	@
��4T�w��XNm�J��e��,�pm��ȍ $���7��ѵi��E;h�[}����Էy]Z+5�Ǜδ�C^�U������@+�N=��b�:q]�vb�;��-�=iK!�)�3�gAsC��Lu�t2S�SB�N�4Q��rutt4R{(��m\U韟�]�r��6l�J̴�uk�\�5��Z��L7��Y	m�lȯ���f��>�!��|u����G�1M�F��wiwUf�g�4-��Y��u�9�>00�W��1�;��1ڪ�f��5=n{i�R�A�NXJ�Z��咮7U��� �L&`0Jh��j�t�8/"�E�6�P���-���u�vs����nM�?0X�^yfi��sL(Y�.��j-�V`+ݧ5ފ�v��U�L��A%�f�ٞmٵ<��I���|#���[��/���e:�	�7����u"ؒF�d��-�$A��"YA�;�����R��:��%,#�6S�Д����l�p��R�w��\��Uh�ܿ���^�n�Dh'�C���\[fuㆫ۰.\�/��(�ɗF|/��k
ɍ��(Չg	��޺��'��8�š#?��HX��) F�����VK,�^�t�iq�H���U�=�k#�(�҉T�1ِEH��I�皕Ю�M���Y4���s�	m���.���V�ƞm$��P^�Q����M�g+HqoX�E䷝�M��#�W��G��`T��1i![p�0չ�DL"��h�l�uMh����΍��vL6nsi��uY!��lb���m�g?H��E`j&l�(�����|�;	���o���?����s�K�C)&��d#���0D�Rއ<��W\122"�`��x���={]|��\�)���S�k��F#�=��4	L���$]>4.���L���\�k�u,���޵�������Waj�}�{���o~�ӟ��sw���躿��w�����?�$���T1IF����r硞�[��_�:�w	���N�
X������op�'���>��Q��>��/�<TF�\�L ����������d�l߾�`��|���tw�E�M<P��"�^�+�z꩕aD-8}�%��&k�ځ�w���߿dx|�n��K/]�����M�,.6�U�����e��YQ��q��w�kp����Et����������_���ɬ���.��'���Fia6�9;3�x��Z�b�#��Sq<;?�ȭm�����^�nݓ�����kG�:���/��
  ��IDAT~񋧟v��͛׮];�b���t>�7���\�Ț��|��{�1���>�f��۷��j�$e�v�&��٨���>���'�_���Dz|�*�!Q�g�45�s�Y�}��Y�r�2{��mWjg=Ƨr�L/z��������_X��:Y��;:�����n�Ե�����E"(�ɭ��jW%;�,�|���O��в����	�%�8�ʢ L d[s<_x�yiq�M�o�ߔ�� A�3ɾ�e�W�C��4����іɮ�_YF���>����%	6�j�C�D~�&q���%�aq%p1�.�Zz����!�MyԮ�Cf	�ZH
`l����e��J)/�]toSJ�ZR�EA�H���~)�G,?�1Z��U�������,}�����n�ڵy�1^���*`Sc$��\m!Y������kz�7O!����Y{̌6n���������nX��'��pKĵPm(�!]�,�`r���@�$ܘ�^ںu�aWh=���E]t¥���^���*U��g���;���ԗ���F����g��w�=|?��333�0p�at�W��~��U˨��2����.p+�>����+^�
Z�"�h�����C5�g�Zm�J�򢹕����8.�h���AL;Mo��2.��5k�"V%�1�u��̃�+��D/H��(�h����9�f;&�N+��]kt�jɦ��M�ݼ�D����I�F+��O�6Ѓ���g_������MV�����i}l�b_��!���R��Z��4df&���+P�E�COݫ��HVpQ��4���S�e,���\��<���3)�!�;���x�S8�>cB�{{snXbrx�%Ç�\�'
��������e<�_ -a���i�>H9��#����!	iA��}4�O)�2l��E�#LCשi���Q����̔&Y	�pE����#O��y���^��$�v�L��(�%
E�6V�h�x�{eW��A#��%yIE��] ���^$��S
9���4���9Lg!��CtZ�\�\m�>Z�R\0i)�?˄���	Q̫H�e���`TRw�xQ��x�m:
O����m捬y��vI"���z��^q���h��)�_*e���.k��,+m9ZP�W9�����H�ɇ�FJ�U��L��ட_���j�F2M���+��O�s�]��50<�2Q�W �`��� m��=�����`9'�%#���z��(�KUʺM{(��!�vgz��^5m�:rM��v[t���[pC�
Ӗŷrf�JR��l3u m����Ņ����_e��<N߸�ܳκ箻��V�$��˟�����?��F7�H�h����jy��Eg��m	�<tBz'+���J��|�}ĺӏq�����11yH��1�/Px,&�����9��n`�E�o%��z�ۻ;�5�yI�Ԋ���~�n�p��_����[\q�,�P)��2}`��+U��=H�G���f�;�
���K2�h���S�����#+�}�F��'Qݳ��fk*C��v�l&åƂ[�ɜ�����`~n��=OP����0ң���
^Z�U���rm2����C<5崚j�P��+��̠U߻[C�I��<S/��JKhVuHy��wH-�*%��g�9x�-x�W�*v��ٽ����k6�X�j��d�m�&����@_�l�-B��/BFM�m�ɓ}��n�ZaT��T��Gm���N��2�yF�%YiE;l�E�<Lv���;>��v�s��i�@*�[M �Z?!ΚY�?6>�� ��|�rf#/��(���c�<&���y�R�f{׍�,
�or�d5�۴Hf������_��^�l�Օ�KU �C�����Y`�V��sK�L|<W�@+�\�!�A�r{��2,��H��Ȋ���;<�5�<#]А̡�y�.� ]�uQ(��;?Z��s�d�*?J�;:��iGt��Q!c �Od�Et��(#���F"�Eqn�YQ�kv���t���-�^h��d���`,��f�&ʠ���x ��KL/O��n����7^0Q��(��N���nN�2X/���|"���@	��n�Y.^�A�`�������(Skao�k1K���$ӑ'f�?�N�Ɏ{��}G�����TO�f����^��a7yhiN2"LR���$����W�-�P�T�8�tUeji!ʒz8��QlXMKkE��7���U4Z��o��n��:o1}�b��"�X��1���I"R��3�M��i7�,Y�r���}��ﴦ�H˚�t~rbzbrzfҢ=�e�:k�[!H�f��o�iF(0+N]W��u�V9�>=>N?<48�?�nMr�HA/��ܔ�H2�)�����'�~R���vk�F�/�I���y�-�ț�&�HZ^n�G׭F��*̼����G���@�6��(J�����k�ӦY�'s~�����"T���!m������@��kE��d(^���*���6b=[U��I�p a��_�;���uϵOظ>B�2�5;S��iB��!����W����40�14����̕"�e�:́��nL���ic}rm}V�[8|���T3q�i;����C��b������R �)GC��-$Z�V�`�*���܀�y}C6��Y��.M)��΋�@>`�M�l�0�HXv�"��$�Պ,dҖ�b�Kڪkf�<���G�&d�d	$���^f#�Y�P��D{�̂��|��H�+LrN�m(�K�b=i�w;8[�Bn���(E�G�r2�{���3 ����cp�X`�u�,�)F�BBa��s��[	M��E���E�q%Xn�ʘ�Ȃi�f𡗄��5�X���c3�5��ԺR�c�[K�8���b�у�V"��R���C\Y\0�ye'N"Z����kg�����̝��+�9p<ok=ˡs�>H[�Kew�qG�Ѹ����M�s�9gժU���'~���+��e� H\�w�����/���w|����o�IOxV���t&����ł���{Rl�^'��1������v'�w� �^"��d���y�;�;��|�w��]۲^����~S�ij��i���_���?�q��}�����w����]w���xhh<�v�8 #d�T�����kJS�0�O:zo�W�x�)�FR@"�X���'�T>*O,6�(�Z�v��5k֭�����\�� j4��W�n�b��5I�R��2 i\�(Th�$";��3O�3=�"��jkh��&���J�B:�p��͛����ݻ������o[�jU��d�f�����p^��4�G)7�I�t������w.,��g)k������T��P���������4Nd��L.�ۤ�Ɍ��ONN͓��N^M���/~���pÊ���^������gfA�[�>�M��Z'H˔��֭sZ�lԤ�h�����E!�L��B24�S���j{���?��۾�������/x��_=�ft�޽������^�N޲z�j)�pB�)֪U��A�D������"-[FKk�<�hGGG��ruT�Ԣ���ZC�g���L�ϼ�Y��^�S��p��0��O�\��j�&=}��366F�il����e{GyD٧hr�JR	tG�K�W;������y��=�eLǒ�+�b�^�5d�����t>�h������!��s�Щ�:z��^. �GҖ�a�_���yI�A&>��O�)���ԩK'.�����ʗ%''��'�1���q� �Ի�}+��w=�O-���`��h`b4�Ǿ���s����A>X�h7%)�i���}G �]�^.]m׃�i���-�*A?�`;\ ̉�HߥKѪ�8���3q�oܸq�T$�����M��?��-[�<�o?}kx�0�B��}��l��#j]���\���;.�h�)��r��?���S�>���㼠s�v�Ñ��T¸�Ew���y���^u�U�e�ڵ�[n�Mq��O�q��9�j���\���tG:�n:�3.��R�~��۷o��׾F�T�I/��C���-�?8�w|��*c�+�ͮ2i������'?�I��@���]����Y'���Z�,��C��f�D[�n�trs۶m��B�Km�:,��":��y���1��\��z��j�֏o�v1<<�qsA�&Y��;w?%d��59r��O2��s�%�x��7�|��'����+��B��}���,���O8�������
n�@��@䖻k���qTԋ���mN���ή�i_C�����m���m�����(t��Y��6�!Z�P��U*/�%��v�(*�t)[�;E�!�D!Y���'��'�� ��7(��MU�4#�0�"Iy������:���M���%�Uti○��R z�k����tf.va���Ľ��-QJ؇63�'If��arAbf�#!C+ۭ����¤J��79e3��,ö�g2硙�޸ ��Tm0����E��/�<�eˠ[,�!2 �d6�髴�:�����y[�Y&�+t�F�u�����W�_z�ŗ���+��_��������׼�J$�h2�$�B��D�o����������$$&Pq������q�G/�W�`qO�_�����:�Ļ�rYN'$�+D���eS���:���$-ǹ��{�i�ӎff��� ��]7�@���7����m-]�ė��?��d�c���u�ｓ�&I��kO�ǯ$��s69C��E�Z���եh��N%�U4�ik��c��r�m6� N�ԫ�V:4�W-�3st�����SsӤ5V�T�m��@ka�Yj��-�4۳̌klH���d-0k���%o��j�r6Hg8�cH�C�~��&8T�+���lkַ+��C���$�T[�L@�O43H�$KZ�J�E�vɦQ�VJ�
��q��ܰ��`�C#h��VI�N�Il6�T�njp��f�Y5gkJD9t�����X��΅.p��ٿg�ڵ��C�v+h�o�LMg�4fU���y'�UФ�]J"tg}�2��Z�%g>�\�VrLk��Hcz/M��ۤt˚;�j�>�]��Cal��6��8��[�C���Vh�焆682̹��C'Y-��,���D�F:;LH	t;ex%[7�������m.���8`�d�Xdf�蹝TSr��22�fC�ӭZ���Y�bU�\%艴L�'$��B�|�@������ʻ�z0�Gb
%7�[��q9�0W����*�e�9s/�ÝL����;K[�G�3`d`�!D^.�I�p$2�;-�<粩��9>1�B�Q$}�Y��G�#��1i�G�Z�p�44�h�t�-:2����Ҽ%�(�,2��1�K�k����+dÜy����r�P�K�X��&����@��	��Fo'�v�$�CW�,�HR�p�F<�.�l
��V��kd�k�8�O3��Ig.zF���J��KYV�۩c��YQ�
���[�o�FZd���Y���i0����f⾲�e�H峍���A��s�?B O�wR(�����m��
$V��%EIO|<�W߻{��`�1��}���M.�ځ��ǋE���,j�P2�i��z
�L8��v��0p��+G��4��O��m+��}O>Y�,�'�|@/r(9Mc�C���,q57g�g��D�H�h��K��G��`�m���H�����*�I1q��EJm�Y�pfy��V�͉$jY�GiB u�D�D�I�7KI-��~��ڃ5T��A�Y_��
.I���qJ��9�P�<t�R���X&h��3S�e����FK͚�M����jzt]��sS�f�����ܴ�N���tF�[וf�cr�P7&������_��Y�B-볧ؓ�{^�ī�(�bd�hE;�-�p���pM�UM�x�p��_9R���=b��E��u��GNJ6�E斦�1��<K�+a@��֌��୪�R�H�hL������iZv8�Q�w�5��v�Y�R��ݓ!�r�SwՑU��R�%?�'x��*���c�W��0�9@f����BH���+�O��Y�d�ByP��`:��	���/��)�� �e��w #"���}��T���?,[n�!jZ�	y}���R%K���>G�T�ݙ�SnO���ɨ�(T����y[�Y�(F�L�ˎ;&''��W皧�d�Z��ǯ|�kEw��⟾�Oo���ɟ��G?�QC7�>�E#-g��pP������%��Ql��X���[��3�9$?XB�/���P��%=A?�n��P�x@UX����Aٳg�Țu��6P�i����{��_����}��~K�P�q��$l�Z'��q��;���k='������x�#�Rx��C�}�=���A?Hjjj*�3� d�T*���������f�B���T�:400�ҋ/%�2<<<>>.�yq��mj�P�G��mh�O'��j�E�^�c�=��D�@�w�bNNz��^���ѥFFF$J044�b�����S�Һ�]5Id��C���J� w��9��,��՘i3G!#� Y�&l��2+�MR��}d0�����-Ч�z�R?�af����ݻ&F�L�UY�����D�
����G�vL(���u��0PEӨ�"ќ���=�� �2�q0�T�]������a�� �攣]���;ԥ�y�m�������䌭�J=��DIE�P�Ȑ�77�����򭎾^�eh�r�`�܎3�S���Em��V�B|�P�N��,UQ?33K��t$X:��'�|r��x�y�t�I�zի�?���yzŖeJ�f	���4�䍉|B4��z �D	��x`-��x�qd�9�dۭ&��8����n�'��2h!�WC�V&bE��٩��1���k��F�����#xu��u�5�4{\[F�q�m>_q�� 6z{�th^�!f�\A����Vr�(!:���8�����iCm���7����y}��}��j��A@�Ivͻ�-�����4����3��g`
9@�nu�����O��怏J�.���Ŏ������d9�L]ڳ4N�
���'w�9k7n"i`V�d��V�YrIv� ��ԏ�G�jfffv|��{�&�g�n�喕�W�*���/�53��H��/��m�n�Dp�gB�<�{�G.I�@���`m�Ν�~���L]�%N~�w�/�dW���M��}ϩ0���Єӷ�<���������ӟ�t�	�����%�]���}�.�L
���3�s�)�g�
�A�w�LH,�A��@sH�s��ԉEIH�T��DG�>������r�m�QJ��6[�D�B��b�h��|�����(Y�$�:q�"4rp��իW�ZE�8}`�flÆ?��8�}ՄW���`�A4W�<�ݡ�{�	ܶm]��5�iJMf����fn[=_��=�M�MM/����ÿ�6�:h���FTS�A��O��A|=`ӥ+�>EPN&L��_�7�� Vt.p?��8��"�i" �
֬����M"%h�fr�R2Z,�;��:�"��^������_�,?y��-At��A�'�ZV0r��{���z���յ6IKF�@̔H�U(=td�&�(A͒z��8���e\b-F���3Ƕѿ.��X�q�	�J<6����蚩�1���B��K`$��`uK���ۺȸY�^��e��z�>���V���Z�r�����L��[߽)7m4.5�6!F]+j5�����#;b˖-���Q`��G>����g��_~�;��a�GWI�%qz��2\p�XY~s�3C�i�r���Dr�|���y�&�NT�����ű��WFs��B���ݿ��_v����$��h���s�=o��;��ƭ���o��7�=��?xs�.1#��w\�kW}�_|��^m�b�8�g���t�x��+2P�Ѫ �L]r]ķ������e�'I�\�������k�,����B=�<���a���r�o��o��]�V��zl߾���BO���V���6�q"�{��m���Q#��(%��WL�̒iRɥ��b�@�n-��eq6?=Ә	���"��x�X쫏��n�3�(C�Wǭ���F�%S�2L��34qIu�8�u���X�Zg��9���!��J�T՘�:ig�3���p 6��,�M��|���d�_\h�[Q�,v��J@�$_t��0cL�N�0�o��z�.�p�A���hirj��ͧo:�4�ƾ�'���d���c�c�-�tvi6`���ɻ�>A��cq��|�艪ij��3�l~i�ԯu�׿3e�Hx�6m��+W��16?�raDY����մc���������O��\	�n�5T*W�ܼ�����=�r����Fʕ����v�}ֆ�+-C�e�O.�#�̹������^���?�3�����b�q�a�8	���=�^��.^ZXZ�ٹ��F�����Nӧ�z*L���!��kח�X�r�&mM�0ky͚U�:�Jhyת��� d94���}$gj}%(��U�W86�C��R���@�$���9ʤ�}�A�G�k)��(���lk����w�M�#�91~��/r!T�`��@&��j�9��aڑP^uӋ��eXp���I���]�k���M������hцX��$���GǍM�	p�t�M������C`n�B�p�9�^ܶ��Qk�ۛ� ���Qu�*����
J���⨚*���?lXI���͛i��v�]x8�B������<8lf��?�Vw*�����=P��`�>��5bC�e�/y�54��՞�x����������k�l"/:l�������^r޹O^�jO��o:8<���S���ɼ�\� �/v�0���el���("*^ڍ��pe��~L2���|4[����Z�j�O2:M v�:T)�$h�|x��N���
��W����ĸ����w�Ga�Z"�n�=o�nMg�:��i�i.a�.�Cc߾}kW�����}��i�={���"3a�6�f�~�:���dZ]g��8j��?Nȴ�Q�6�N�M�Y�[)՜S7o*4}�;k��7�p=V��^sE���/ظz���Dṯ���{b�YOP��Z?�k��A���_�:X2"B�v�'[�R� �o��.����e����L��3s��&8{zYR 7�U�i&�i��	]E��̙!}����"ڎ�������6�0�K�JBR���_J��/�Z�hB}h�N��p|�!Ҍh���T��r�(,#���qu0b�B3e��H��"��F��y*
JD�)&?���{�e�_�'@��o:
�	y���
oSτ[�����É6�vP.�-t۳��E�j�mK�i;+Ft�m������e*0�&�25<�V�əJ:*oB~)))�7�|��%A (g�"�L�E������V�^���Ef����Y
��\� j�!CBT�R�9����D�+���6�3���܅�G��Z�r�o��Y��o}�~3>>>44�K�$'��տ�緿���׏|�#�̇?��O}�S_���{�[ޒ�"���3�(qx�è�{���+5��Rm�#�Ġu�$��ב]�u��5�FOl���3&������׃+���DR�,@���#Xw�)��
��O~�cǎ���R	�k�U���9��Dg�SQ�)��p�
MӞ�hy\�W)�����=.�M���K�p�mڴ�@��訙��������b&m����c �''�$nyrD���VbDtv��ܝ���!�bsM40$-�@}\�XIWPo�Y	xF�SB�?%�hYf)w��2=z��o��(��i<�gkH���(R�<���O�] ,!�F� d�\t�Et;od��2P6��w���o�>�``��d�v�2��>�-̌�O���̉���)�@�Z����#k�4h�W�^�%����"�ni�Ӳ`�Z�Hw��a�uA�ka�n���kN>g+-�z�ݻwϾ�H���dG�y晰�ܖ4���O�'��-,;�}L���H��t#"">�$��?m�Y~��矟��֮��i��}���cc��~ZQ���(r������<���@�h��,�p���P;dܝO��F1e�5�� iPY˳��u/��&�<!Z^oX����q�8&�"S$Ce�.ի�1�����O�� J�5$���6\�7�n ����n�D�J㜚���XIڴm�W�h�x�<4j߷��[o5"�|�6�Ou�N۸q��`V��y��33E[5	�Ђl�Z�V�%xxxݺu�/�D�BIԑ�;� ˙�mq�E�Xu�ҹ�8�@3ǽ�C�*}kaa��\���@�[����¨v����6��ؘy��~nҳ�	 b�Hѣ������Ag�xTHc��P��!����r�����^��,W�E�d]
`;���f�W�v��
n��ݜ��,5eEu:��L�b���wc0zn����8��~��ȫ�@�m^��٣�ĥ�DJ�C�I�z� کVi~觮Or�g��
+W�f*�7{��0�f;����mן�Z����"M�!���W/�f�@B�֕��ԯX�<�D̠|9��[��Ocn�*�ؙ�z�':�]r���ȝ����W�kr;8��;���x�{@��N`4-��@I��Ϗ���6�') ��4O;Ta&V���0*W*JCwh:�2-2���M���:�#������|�uZtɂ;J h���_*9�����J=����Tu��'��c#��<���x�[���J�B��tn\��k�i �Bd6Y��n��yh�(�,x��%���3�}����F���ia�ٝ��b�=��^W:a�<rA	�!(ߧ�O��� ��$�z�_���s�x��z�C�����/��[���>V �e�K/�u��|�s������7������|�������˫�V0�0J=�٤��i�`@v܂���S�z�\�K�=G�t�;�u��$C�k]&�(`���X�'�Tmi/�a��@:",ƿ��'��W^�:���|K$�dA�7^s��?�����s�y�k�Л��-3E�oJ�����77zTZ�{�_��K~���ѐ�[��z���/��5���M���I�	}�ڦ��1���^��%�=;7�{��}�oP׬J�?��4��s��$΂�����XS.�n��\�wyd�~���I8��׬tm�o�>���r[���$Lt���LqD�l3u��dիT�V W�����y�j��$����5�XAB�mp��V)�^p��纤�4��8O��q"�<�m�E���d�9)�$���@B�kL��FG�^l
G9���z�K/���?�F�m�,.�^xڙ7~�_jzژ�y�'�6�4561^���5��v���W_�F�V!�ʳl��*A��ߞv !*N���J�@L-H�0��E�.hsè���֭YK��;�k׳ׯ]y�U�:���<��SO�߿�ҟ��t�yL�����#���?����ccS	s�2�*���g�E����]N�`,�m(ɱ>�`q��Z��kx����m�~�[�?�s�Y��{lz�_��B��RAd��m��%�"pAp6�y��$�`Y6��蔏"���l�-,��SfϹ۩I����Zϊ:�ZJ�@F���f'�iu8��e#K�u�D�L�9�O "�޳;�=��U�6���[Xu	�!u	���݂�itRA��}�3��Se�P]�� �M���a�P,�a��`5=餓�z�+�7��3$�V�]V�н��Պ�}�{���X�8޹s�Rs�����հ��>=�HU�-U8���6�N��r�%��ӕ;���U-WL�1�^�ʃ}�充(��������$
m�����M�ޜ�?���}A^�A��+ˣՐf��S�|~va��݈�8�v;4�\7�3�>��Y��"��8Md%Ȓ�8u�;�h��	!y�F��LP[r�ڹ�58BB��22����Q�Uha��V�{�g63�E��˫�5�V�eX��0�&���mt1]3In&�m�\�k�xwꌀA3�i5�
���x��XE�v�
]C!�X{���[kS� 'm���,l7��fp�%�[xj�����ڵ{-'9ir!��!�O�i��_����M� ��f�j�ŅF�DpðM/N�;w>����̑+l���k�-����ӓ��<&���1=�W���Ҫm�r���(S�-�b��=�E�^���<��?7����u4�ő��GZ�+65u��	 �	��w<�f�4�\V���BYiNJ3��04J�%��}%u��<2L]�6�����F�^a��
�,�2ɭB�	�K)�7����M 
�0M��s���EWȸΎ{k����rܯ+���$ ���rfyY�vA7G�X7�%�M	m�[\�(=���yX��(��2,o0d�7���`W�f0����:���J�[��s�(ǀM�j$ɀَ�F���qWa�YⲔN��cM�8��n�l�ķtR���9��MAk�,�A��D�?�4�PH�MW�
��݅�:�t��s����Z�~w>��O����_��h����xpoy�[>�w�p�w��ʗ����9��w���}<$��~V�Z�=��#�n]�`�����C(h$���^��S1������J1��Zh��]��V�(��Aqp���!�[v��q�ʇ>�fPasB���������g� �G�A����5�K/��E�jơk��euI��������{8���\t�rʜ�3ҨK���,7�c;�1C CH���B��%�	/��{܄�l0�w�ظW����h4�̜��~�[k��#������,Fg���_V_�����1�ʄ��Ca�0���z�n�M+MG~�*BE�ARkԬ���G�#�暄2������[��MLLH��`�.i�Sxm���^�f0hI����|D�L]� S��đ�!]޿���xـʑ)CU���0x��[ӂ0kK�,���JX�s�Mő�Q��#h2����p#���y�V�U�G�jD�_A'[��`�	�[�7�73O�>1~����/G����]dbb���6:t����-�;a�ڞ#ǯ9��s�\�rFK�|�2m���KW֫�G�����߱{~~aH��5\��m��	jAC2��O�QE��Z���-[f�ƃ>x`fN��>==�lv����ȋ+�`���j�Н�om�\��4�	𬦎w�����!k��� ����w7�_���1\��r��&��C[�n�;1�n�:z��˗'&�M�'�V�/'Y��Jl����H��~IP8�j㻶e���@V��|���)~5���B�z�$ �O*M��FY7�.h���ɒ���_����J�d薴j�ä]-XG���7�1�W���$b�К�fQS�6W�=��-���N���HZ^�\Q,)�H��A������ذz���l�Nkx��=CCC$�֚F����Z���ʁ�0<餓�M���j~^�z�M7��P8m%��p�Y09�MTo�˝X�H 2���\�k�T.�S��	�
@JJ~<xp�}wc�., K��'�	=���	�D�@k�c |�6�,6�52.���Z:;�Z� �f�;C7��Y�k��Szrn�5S��H4�|	�ʒ�!t(g�Ŋt\G�*�����<��1�a~QĒxO��$fvDa����%+tq�ȲG���#	�V˯��c��L�_����ڄYB�pVe�¸ӨY�]I��a굺_��)Zp�i���B�tٲe�:4/�����a��M�q�� �59�j��	y�XG�x��^F������-~%ϴ�j��te���K]y啗���yl�'U����x�8��y7U�_���䏃 `�T�F���ob���+Y��ڵ��n���Jo)��N�R����w��'?�	��h����7��GW%�,���pr\f���w��}�cV�S6�z�7�s�KVǩ-A͡������KwĖ��ٔ������3�ǌ�1c۝xa��I�Y�EOr}l�;�.0�b_q����?L#����UW]���/�%_��I��E�|ཿO�m�(��y�`1���3N���Y|�-�(l���S��7����\�3��!	���߹�J�����E<!���;֪Uk>���z׻ޞ��^�k�p�k7��s�w�]{��ǟ�.�8R5�[x�;/�����_���,q��OH4��rOO�ւ;B�L�ZJBVI��[	Ye�ґ��s^(��"C�i�3��A���\'7��R(�������ƈDF�Y"���=�>@�\���ҹM��Y�b����QAA|��v��<J�YU��T�H�tG&�bܬ�6!T��ز���B��HS:�,�a@�SA�I�!�iR:���ΉLK745�}�5�V�$�e�~XK��Yԭi#��z�)��	�?6HS�~�*#;7�Q�
ں
Y�&Q���u�j�&���84Sq����(kQ��+�)L�ZÝ��|��v�G�T�����<l��'�#MG�mjt'�.#�@6X�"����f��"���P'c�Ђk����2ô%K���Qy��T�kpE]��Eײgj�g��cm�Ugf��J����KnE�uS�j��a��Ú�|l�.��7^�f�4HS"?�&�f����4�4�-,�d��h��_��u�<c���7�pC�o���ބGd��͌�q�V�BolP����8X���S-�����Nܸq��ի���0qx����ٹ��_�(X*�ɠqm�%��5�b^�LmfF�p�^�V#��b1�I�l�"lQ.����魐�F�?99���ҥK#hP��yd�7�����A�} ��Bd�k �\?V��:,^��e�+��L��K2 ����ն2Ɔ#���j� }p��q�DJ�B]�ú���d >b��X�ᆬ
�d{5l*x�/w���{d��̒�l�F�¤� �:������J���A�8���	�X�9::��Ӵ��T�.h*P:j�wHm���s�r#��\˔
�7|B	(�㉉��n��[_ف(�B�<�0��^60\VPŋ[��Ԕ�C���k5gfW�\*� Y?N�x�g$�}���t�}�Lb��Z�d6	ߣGaL�>ɎR�0����l��ͦ�V�V+�K[����h�=���<����<|�Ϯ���w��۴���gP�M`�۳�Ȱ�pji�d�Uq8���߿h��v	h!{�z�(d2�1�
��z�]Y�yP�4�M���1�Dv��_������aqz05�0�\a����Z�0�P���h%�5��n5��i��N֤Ab� ��\U^;�7�'�N�V�EC��-��6C��$���,��)g#c ���٬5f�Oj,�*�J���)U��>d�c �ű��'�l�����E۶�}���h���7>���I�VK9�6���luv���e���������y�v.b9������Fl��0�A���`�h�7'͸� �I�*�d{����p�#��gb8R�%�>�RE�Ѿ
��#�<r���잆�'i:��K/�'#QV��]p��+zS��#1_Z�H7j)��!��O;m3b���E[u-�A��
�����>�mF�
�2�뮻�����}���3��mi!�ԭ?��?�����fKy���I��ؾopp e-���Fn [S0���G@}�N�5��:?�iy$H�y	�KD �n��q;��TXn���+��2f���A�����������4K5tS��Z����}���?ںuk�p�L��S*,4ZJ
�դ%m�Q����?���S6E�f ��t��a�w�η�������-�����]��\�i>t� X�'ҲCO�������:��F�kշ&k�%.��A��yc����~�e
���3�0�b�푍�>�/���(�ќ_�/Wz�����	���Q4�
v��O���f-L/����M�{�:����c�+7ب\�CW��ep�*?���r ��E~�#!�g�$�h����>v�by�>��ڱ��n.�"vfD���-��h��+�F�|�:\�M�-=V�iH��F5-���H+��3��'�W�q� 骀�	��w�Ak<���D�����LC��G��-�"%��|"�5q����p�.��
?!�8���~���V��e�dR�F?D���S{&�0 �mץ�W�N!2@v��O>́=�JeQOIJ���Ĝ0��S'�p�k_�Z:_ �ˬ�ja�	Ɖ)�]+lӰ����t�摑��哱KCz�E��#?��t?Z���  6�s��T�������K7�� ��'�.�`݆�-�{�M#�K�/9餓=[m�Ķm�H�eL�E^����-�K%<����@X|Q� +��`B8�.^��i�2^�f�9眣.^�����;v,�q�}�������(��,Y���ܜfg`pޑm�
�_e�"|��H����@�/Kf�lw˲�2���c��<n���¶T��Mbsd-���H"D�BQ -�C j���莓�_�	�P��N:������ݞ�1ɮ�_�7W�xb?I��"�Z�E�(00�D�RD$�sMn���;tQK�Eْ�ЋTz�iT�o�N38�S���!�u�	/'?m���~ �����Π.�ꩩiڨt��0٥�����t����|-��>W���^�Y�n�$��+�Lh#e��:$�H���)R�n��R(�l���N�Yv�-[Fˌ���͢�7����J:K�|_o��B4�k/P�<������DKr~���	PM�g�,j6��qĝ՘�X������vS�_�Q׎,N��<�B�DS;̨c�9�g|V��������^�*-�.�<3�%��W�y�b�E�K��W��h�4�$�ha��,��kg�l��޽{�8|��'�ǧaB��@UJ��Ml�§]K0��O��Xo��UѭH�{^�1r�>�游+��i���&����r5E=���<d%����Q��C�s�o�-^������!����?����^x�w4[�]��V���;���]�uڶ��ԧ>�_�ꗾ������ɐ�@�'�=��������я~0!y���ǿ�}�s�[�z�����(A���;�������ƋI�kL��K�|�5�|�k_��?�;����&(5[m��ʿ�3pTԩ�xA��\�c��.�V���?���K}��^�������U���=��r�L�N3r�=�{�W�,Ұ���Օ����*�ܙ�8j|����ʗ���o]� �� �8�K���;i���ox����j��a���G?����߿��/~�T�e��'�ڄ����!�����nWt��,_�P�/�Z�s���r��Ɓ�Ը��㾺��U�T=O��mh��H��#o=�l��j�&)����E5Հb�!�!��xa�i2O*�)�g<?�<�]�V��JS�~	���0�8)K�t�*�6�Kɡ)��W�$�:r[�[�3��iJ�k��a<��#���5f��X��<�*�q��Rv2H�`G�5X��R"�N)T�H�[�*��[�\���&PVu�v�X�@�ӳS���X6(ԟ���3��4�5|�H�5�( �$U��F���ѥc333���M��yU�"6Q�04ڷj͊�e�a�hף ����5,=�r���|R0��h�{��A����%��oHGq�SUB�A��*�}�3����]ƮΎ5C�1�����j��Ӈz92���S7²�>=��Ql��5�ٚ5��82�m[����>�� S������7�p�6��"x�r`[�����������_y�Y�����Eq��o8����8Z�9��[)��>U��3~�ջzy��l�p��}KGF�=��̡��<��Rlm�`x��X�|����g�ZԴKŒU(��,�Rf�帻�`��)ӳ�L2n�'�5i�g6sUg=���f�u`|�^]@���CCD�kŊ��)�m.߱o߿����.��Ͳd���עo�}t�xI8NA��{GiSl2�iڶ��K\�|�Zٛ���� Վ*[�Jg˪�T.� 8��?�]H���b�d���
y)������5�#a�	P*�2=�RI���.�|Pke�M�zj�.9�Y��1ѓ�xˉ�� � �k�G��4��������?���B�=�k��HѦd����r>���䙩iz�U+�=�LbI�y5�f�[n�ς��i����\=E�R~83�v,��n�0Q����`��yC��{Ɠ0iցp�Ƒ�ܤݪ%�:{���c���2��|�e�nBb+jE$���-_��ė�.ME��O�RM�^@�w!X��GBr+<���Ќ��-�����={-�Q����k3��?%RK�.���=�B`o<�ى��0L ]�Hd߬	:�ر�%��䣩���s�3g0�b{Ekz>�8J$i�v�m�
�(^Б� %���+���␆�i��t�b���� rl�&�	�Z20P�7�����Tz���H��P$''B�w���@2�4MOM�L�QX��X�-%H�V�7n�I�b��
��������}H�h��������v^1(B�wGQ7A�Ƭ����hk�L&���H��:qʑN$���udm�,b�{�^r)M�W����}�{}��#�0�0Z2����ě�q�M7����[Oߴ)j�P��m���7t*pq[����S��o����ّ�azJ�*���Ic:��>{�{�c���7�|�g*(I��EM[��/��>�'��~����k/|C�N��ۿ1m���_TnI�Y����Җ-����k��O��X�t�v� �Gm
��X��;,�����ft�W�W��@O )G�f��\�x�������=��ϴ�����������d�a�.�`����[o����>k�Y~{�2��X-�ҵ��|�3���\���#��K�kD�ZC���?����M�7�t4�t{^�����O��u�Y���:��eKW�N����G��9羊�4.�Ur�ڧ��$�~�J���x��z�C�4��k�v�t��7� ߎN֘ldT2��
#_�*�[`a�����E`�����g���0�0�g�e~���Qq��Uf�����P"H�R��z����g>�3�{���J�*/�#O�p* �'��c.Cs)G�?%~�����$��߹s��.�����>ڢ���O<��=�呑���������2���d߬\�h�s����)ߏ����Τ��ۅMĖj�<��A��WpmD[׮]{�y�/���{w�?@��[&�.|A��dG��a�YV/�����{P���i�f+��t2\�l82�U�g�N ��z��0��Y�ìZ��|���St��ԳGGG����"���8�������I!b_��W�lْx�իW�5�]���M���S��Lc��}����?�t��5k�����;��O=��lm���_���e=F�k:y2��C��9������|�<�Ʌ9 ���eF��7o޼q�*�riP�O<|�O<�ҁ���n!�Ũ�)����\�L�+V,���u��&�ZssU}x�>���}���zY�/;u��Ν�h�C�V���[���Oܽ{���C��Ht�Ҋ�/`]��&�dº[ kg£�|#��x^]�ti�{zJl�2�b"Q��f S���LW e:��!�N�C�0:��VfsNe���#uh�:��`ɿ��,JrK�鮔r�)�<M��ُ���"��f�F-��-�IeH�L�a�'�8K��^A�>4����b��"O���3������~��?���X\������؆7{�W,յ,b�B�z�jz}�>�ٴbW�-#Y1]��J#�<[�L�j��!75���@�$mp4��|�����5z���1z������BٹB���x���Q������̊�+�	o���x����"]�� ��5�
�:)R=8},^��L�Nъ���Y�Hj��Jݩ $qf)�v�X�'��-�$
�����ct�-pFq�Z�/g�6Բe >!3��9�_�gİ:P��.�e�X22�'�{����$�Wc�j�s��U(�
WI�t]�Y;8�_خw��q� ��<�ԟ��bvT`.a��LNNV��%/��k`Z�e��F�b,��d�SiQI7`ё�����wk�\ +�΅$	���99��U�R��~g�ĔQ����7��MZl�؟��]�Bw��[�Ve���#�ȡC�N:餖��
�ɽ�̍a(�睴�-��¯�Zz&|�q�/������?��/�q���\��ς �EJ�_����?}�k_��c�֪$$�?�|�85�x������(��w�}��y&q��/�t���nҳ�|̷�S�#N;�%*�����׿�uR�����/��n19O���v���/���Ɇ�4�ex6���?B&�D�@ ����r�a�"�m۠�B;���n޶}�_|�F~�@;ǌE�����������ɕW^��}
Ƚ����׮��ٳ��\��_�R���-�_�6cv��k=�A�*�ZVD�"m ���v1��m$�� ��r�,�|��ܗ$vM#}�8�ǽ1/o����u
71KE�=�,+�ې�gs۞n[���N���V@�3���/�iI��/��J�6D�A�>M�γ�n��)�����/K�%��͜�|���ƚ����	.��\� K)pt�	<P�qw5^L�*/�4Niz)���5H�J.Y����\`���I(���߶c����� �|P�/Z200�Dn�Xܳgvn�!��㈮����*f��`f��i���EKI&>��c���۷�T��E�j��ZE�8'z��,�V�f�v��IP�}C/jE��c�6�yC-�q%f�!�{hjz������`uz���f�p�I��t���Y%�.�dE.�9�0moG 4��wnظ�+^}>}��k����M���u��w�띤)������y����V�u�z��?���u���hf���v�hGF\)�Q�\��
Ţ(�����/go��m{������k6�|��'+@�3'���)�
�#fG� �����姯W�+w���{���6�%����l�X�������v�Z��48��-�[qhr�@N�i��ȊrU�KI���	��,A����j�~R��v/�iFQ�ј~s�s�����s3�מ��<xp`�ȍ7�H�&�;-���Wh:2��9��2�h-�zV����*S7�%wp�wvf�),ѯ%��#$aJ�޶!���a�t/"��2��9�;�4�G8�:��N��(k_��GJT���fSI��14<,ƺx24��&b���"��&Q��vs?�V#?��G���!R���B���JW%O�Ic4e����0��E���&\�
�$Å8�lJ�#��N�	��l��^>�]��!7��~�;ߩ��#��,�mO��V.ӟC���		@�D�K���W�\�M읝��S���%���V���a���%�\-l�l�f�YvJcËIo���2��٩F�z�
��?v�um���͕/{�B�f�k�k��z{h�5�x`�XA7����ý�E���f�M�`�j��c^$g�����-Z_4:�Q���^k��V��z��Yn}My���&�)�!��"�c�U�@�`������w�Z5n��dA6��B��lp1��4Q<i�Ђ��Lr|�0�U����)���hAG�f`�Gu����g�xf�p�hϐ'D;�����۶S!j[	:i}�"��_�l�����:�5V�Yiۨ'��@�Ga��V�|@v�ѯ��z��̍eK�^H�f���MP+Z�]����
Hݱ���>�}av�V5�V���Ӳ����*P%���M6*.��x��������Xe��3�#�ԑ��k����n��ˬZ5Jʚ=�a��i1J)���wҍ�򖷴Ѫ`�e9)L���j؅�9g����iۑ6ST)
eш �
Eժ����k�j%�[��LvK�T�f�q�����q�k^M�΂�FS���4�X��������C�k����l�ɛ6MLN��W�-8��d����߶
���h�ӄ����7~����-��>���bY2Iű�Mr4j׮=�W��B���f�,�-Km���'�s_�yw��Χk ,N"�\xM	���>�`�͙>��㤬�R�@���!m���_��W)���H1IJ��I�^A�%}=��\pn��<���b��|��קqVx,a>z� �0�_ĕ�/�Z�s��L̶�ć��y�3�@���3t�B�腈d'R��Yr�D�)1�#9�rq�B&Ҟ�p���ɄSbɿ�!_��A�����&>������f.H0�K���p�N�J餬R�;`#W��Tu1g�</��#�UUX��k���<?#�b
�_��S�y���"�+'� ��T*MLTgg��c�d���f套^J�ۖ-[�t���=�w���d`������t��bǎSSS�g=W�*��R�Q糝�f���ի׮]K���8��O��^�ZMB�Mu�N+����پs'��3��v�A"� Rs"�&O�8��'���-������D7���1%+��zu�!��'���1汑�T�7�� ��ޥwx�ޝ<�3/^<66F*pѢE��V�kN�;D����s��'����uxύ�����ϙ^T���"��x�I��vU�l��CO��_��W��(��n�:�)�i6F�W���|����S�v�}�v���o���q[�ܶq�F�����EzBu��|���cQ��F�,q��3G$?��`R���3&��5B��g \t+�s�b�e�7o��G�.�VG���G���[~y�}�F>w�����;��¯�2��"�p����cd�^܈�JB�����~:U�5����F�J3N0�+Y$Z���E}>ۤ;�$��y�w�4������${�OaZ�vu�}}J���G��1q��Q�.,�n����R�<�"�;�JW�ė �I��C��I6m�d�!LS�
�LKn%��k�fT*�����z�qk�
�w��^x�뇆��.%��
�����p�4��T4��$�<�d�� zk2�iUhX�8au���|�~'����Ø����h�.7���{�K�.m�[�tb�S�����DZ]�3sbpKq��I!=[�%k�܅�G�2|NSw�p�����O�S�꬞���1<�ɝ��6�d(�R�)� �-���m����ep��6g��]zH���q�f,y�<ۦ2�i=�ܸFW�;|*"��N!?-rV�VKO���Q��G~���$=�E]dZ�$�ڵ���|���o%��X�]��ZN�?0<Bk��G��~��,�0C�d��e��Ng*Von$yBfp���r�6&���鷣}�4ڴ�$ϖ�d��3�r�i�|���G���ҽjl�됑xMDv
EY���&�k�Ȏz���oq��Y�]�t--����AUX�lf�Jת�4�-F��f�bΊ�4�a|����G?z�E��f�ߩ��ʧ�z��^�lY΅%S����KA��.N�tff��?��_����l�^��k�.��Ƿ>522�167�A�����^С>gY�y�\�I#>J�}�q�1�i�䠆<���p�$�SC�OB�4U��s��r��hf�5���|�����&�8|,5�dX���4�4Jt#���,���W�$mh��Be��2ޢ���&Rzpr���^d��ӏ�|��9t����E��5]4NMI�a��Zt˦M�F`҂��@H��bZr5��� 9��]u�H���(�����%�A8[�b<��϶���:{�R'�5B@!����)�.���^TA�wmI-g�2VN\��Q�1���u<�񛹻�@!HI�E�я����Vc�޲y�%�T�c��+A^PC���Z�3[���I���:�[��=��#Ac�U�z�mi�6o�72�GGH�{\�`JU���i�|�^'w^7K@�ݧF��F�I��l���������BO�NX-�Y��P'M��
�Z�#4k����ԡ��ٹ��m���]#��-�\��V���bޅ�jGA �(.���U��]��4�9��"UӐ��9+Mso5; v�]�J��\�����b��h�X\r��84up�����A%��-�ܰ���q+��O<qpێ��X32��p-�;܃�J��i��bg��p5Ӭў��m{�.y����`��6�ڨ= �_@��W��ۇ�����c�Ѯ�O��v���ǆf`�F��k9Q��iXzB�k����mM?�Ȯs
�nVJp�L�)��ʨ(A�c��\�'���~���@>H�Ǟx��� �O5�߫V����o=���_�ѧ���05�S=Ԋ�r��"�ض2l�cۧw1Ɂ!�#<��W�ZAw�� �������|��c�'�V��A@��Z'�Ŷ���*G%�"�l����W�#� �WZQȱ���rS��)��
7�Dh^k{z��Y�pc��-)1�� Z9�{�nI�[���-�M�cO�����}Ѷ�;=90_��)�)پ�A`�PU�� ��#/�}}d@�w�y��^��S,T��[/�X�5k�鹭[�(��XW|X����E�=�Rmf�t����1.N�Ad�*0`�����=��`��~x��o4rK"������;����#ɒE��s�ol!�y\�I֮�*���X��jT�5��z��$�gKa3� rH¶�T
��FdB��e�@�X� M:a�8䁓f$o�����h:=G����x�9��f�zF ���x2C P�etC�J$��,ũ��2����h$5�C'���6����C�"$��*du�� �������I�cO�8���>��c}�29 ox�4����9���w�2xY�J�lw� ���rO�Qcly�h���KTEF�@���5&�vld��ͧ��T�m�V����䇽��W,_�j�n�5�<���?������h^�C�n��̴+�2E^9*G �v���^L���Y�-��h��畇J����5Z���N��Bfq��pۓO-[��D���N����{��� `0�͆m��o����oZ�"�s����|��� @M�EN2���O��a*@���odq�
�Z�ڣ�m[�r�StZA�C�0:.��B������u�]S��i���}�?p�)g�|����ҽ I�e���Ǯ���A���8]8N�Ljc�t�]Y�*3Y�����1�*o>r�4�r<��K9HJ�{�Ol�x���,�ɥ���?�������X�,������1X�Vz�e��C��
$��fm^~��HIE�Ù�8LJe�ެ=����[MK�*�^t�M��B %@&�J�<c�5�\|�T�ضl��1!2�SY��,���>3#ы�x��z�#�b��-�%���AP� ;K&���WM�U��u��}�ф�n��v����M$㰣�KBʚ���� �����/�:��I(��q�ܱX+ewQ:�Hz��HS�;�!~���8��NRS.�K�L��J�_�����`{+����,�r��Z)�ja��Y)R�;u>�sS��;E���C��.��������Uˇ��_w��+
L����c�
��+����~�އv��l���w):Il� �\��	M'��_�l���Ъ%�7�|2|?D(����];����r�/�o߾m�N��5��'��д��&S�i�8�C����Q���֛��~&?��s�!@rYrA%�:�.�4t�T����w��쩩���=BW�q�t�%���^�z�����W~��ǥ��졔y���g����l�4?r����L����;^��p���@��Vl��v��郾0j�8���g�q�qǝt�I�����^'V���TI��^�dIߚ�֝|��j��0��~���X����!ƙDQ�i�&�Þ3�'�m�r'��`�����d��Uz�Q0G�ѱu�ֵ��������6=��S�lْ����rEj�5ۭ�d؁&~��@o
h���*�z�j��}[|�go2Q�� ���i�@�Z=����y<O��3bզq���Y+}�+i�k�������$Q���r ����l[���t2�N�Y~~�Vs��fQ�Љd݊s%ߥ�'S[�0��	��B[���������8q��o}㛨YB?�����b�Ӏ���x��ʐA��lӍ��QD��p=BT�ض$D���J���4����R���C�2�1���MN�,�,�2��t`���I>�|�سZ�V5��Z��Kޛ޺܃*A��lp+w���V|��S��� Q�h~u�G�Z��X.:E#n,����]d2yB��Z�8��y��t�ИQ �%u�<Y��`�&2z�$�G/3;=;599�k@��NK��7���㏧�z���J^�eش#�l�`���/?q=����+�����1'��	vf3g	\o"�c��)�<�v���y�q���+W�.ᾥ��^��޾�;v<�{�}��?B����E�٪2���*�Q�����Ze�-9�ea�q����Y��;���p�}b�EN�N��[ � yb��pP.�I&Fّ�#���K"�N���" N�p�/��P׭bQ:2�EI�xܴiӮ]�:X)����%��}�4)$'ioҸ�D�#�������@[ŗ^z�?�������e�Y������ZG^�K!cݥ��J�B���:	,�u}�#Mt��7�N`$d��R%mE�)�S�.	T6�&+U�ۅ'�樂v��-�=l�F�2�|�Iތ�]�^�)�%�5Vl��d?�G=�xe�g����'�P29��^���,v����^x�_���ÈR���]��x.������Xk�J�s��L�c�`ƀm֌(F�'e�V5Ԣ 	�&�S��?hK����`G��k� 6SǠ��P�E�����n�A;�o!Wu�[��5b2 {M){�l��)�ٛI�6�%�b��i��C'���� ;�XmT`k�)G#2Bc�h��1.�Wb55Xl�+}_�^�["����ܔ�l�-|�h)	{KK5=��)����P�0c�Έ��d���J�T�,P���[ 5P�.a�>��3_o�e|�:��UO��w<��6��rattTM��~ם������4q��2Y�,�L1�PwWOP�C�3�(�״ZmGѡ����o��6n���lw��������[I��� �����fh������|c�o���!�,6� uלo���M6� �dj��PDd
������x���2LECB�f�pRs4"RđKɁ�`b�ũ�n�s���EQ۞����d�� �}���=��Я?;��~C��DMu���O5d�׋�#��(�eU�%+��7B/�����K6�F梍�Jafa֬���*�-_��`om~�I��τ��zH����MJ|�k�5'l:qӒ��qkO���G�
ۭ�T�|��͛7���(Ss���tO�Q�֌��U�@�avY�����.Qy\I��b[$�h�\�g��}�OM�b;��4�M�;����ٙBO��?���((�Э��u�B!;�vaq�FO��`h��=d�&��G���'Ȉ�ЃHQ��HE9�E��P��aָ�^W����G��^���qrTETz�:y1)��M�`d�ɐ�h�DV��X�i��B���c8vA:�l���(�o��!�S�:}�u�A���W����}l��mp^c�Y����h�|T4)y#�Q�0l1�VC�ȖUAT(0)B8;;G���ӆ��k����4N���s�]w���0M{�^�Z�k+�Y�ގ���<O$h=������1[,W�d��P(%\��.�+��/����;�ܲ��Q�^���+�kUt��u�Q�Zu����e��:4�,4H����\t��A֐�>v��*qQ�@̭��'dr٤0�0H��bٷJ����kv��>�z��&�$��"V5�� ��xQg���cf�A '�-�r���#Lu�2ձB]K�T7���H���j��`�,��J	�.�m�$�c�sӱ�(��L�ϴ�qIJ����nx�l�#�~��Y�٨5�ŞJ�e0_3a8��gϾ8h�O53}hll��W�C�r~����O��?8D���O=��c�v�^��FL���RB?�V@�$�Q,6��o�m��h[1N>��U�7x�=Һ��]�+�<o��Ï?�c~�E������lU���*�Ä��Kb���x�VOK����^��.�
�Y��'L��Q"�h�gKϠK��o��հ%�0�=J����f��������v�y�姾��g7m׸�w��;��M5V�o��W��FRPCSq�b���+������T k���6:'S���'VܶVPK=��Yn�ڶ}�O�~��SA�z�˦JJ�|�];����{�-[FJ��LRzg�ֹC��ȵBғ\����7}��?�lj���9$�*�M���t�%�CرĢ�M����^҈s��oy���fIܑ���$Z-�3��+y���� �|`��Y��;��tE��G��n[���C[�N�������{.Kك�{�y�'���4��k����o��K���o�y��|��if��b���X	
~i�c�q�կ�=��駟���.�Eq�f�4���O=��E.�O[�u�6]�`�a5�L
" ���Z2��@.�:���8^�� ˍ��E���t��j�C��*W�#�
H�$�[ͦ[*Қ���|��X�rgiE�e�S�&�%�6�^�C��y0R� �5#���S�֕ �d����\An��I�N����q'%�X6�0|�����^��(���a����X`����KadBv�
(��F���2l>�+�_$���l��eM:G�R:|Q��D���Ø����"�pvON���H��K��i�Y����Ąת�����YC^k�Νd����r,L���童SӨp����?e1��6�㢌bD��Ç�ڵ6P�I7��!�4�*7'�w�R���F�v�.�#8WGT����pI(],i�6_*e$O�Ќ�3¨�s݈�{�9�*+��Jf������EZ��:h�.��OO%�p�6dqis�xYT�Kj)�'])���l����ъ�7O�d�{*wW2��=��
@s�
x������Uˁ�l͊��t01ù�v�s�<��!��X0��L�H!㞇�����5�A���J��z*��\C��5��C+�^��{4;u)�v�u��8c��c7�E�<��%�
�%��&B6:��<��s�G�[m���$��v������w��A.�*�9CO_�E2��'CϠqT^R�H�a���l�hjs�H�%�UḬ�[��:�9�<�%�M�����}���Q����4C���ǝ4�` ;<f"���{~~~|||ώ�4�i�����h%#sU.�k�Ҙ4�5��2�
��n�����S��sGSX*p���4�$�\�̣p�����8��Ö�4;�L`�y��.�� �y)0t)�8C�#d�1��S[��+�#�$��L�O�4`'Ǖa�Aฦ,�2����|Y���-r�m�Ss�5��B�E�De$��n4%���6��?�G�BIF����|����Ζqr]�.p)$�w��M���9�RX�'�®]��m�F��
DY�E���fF�xLD<xP�'�|��)�T�[T�Y[�t)�EV���ľ}�h�Pe���4Z`G�B�̆��,��З�����3UԬn�#�3��ΈB��a��]���覛nZ����3�oOmÎ���hqny��l��"tp������[8��0~�7����^{���_�i��(�"A��4��݇��?�A���޲@F Ӊ%HjWfg`��tj�iz�p�f~� $O��r`��D>H���)�>Fu�`���m���)[�"oeI�x�Ua${
n��m�ƍ��M��/?���X�X�2�B�*�$�AjO< �� W�/��B@ ���<�4��]G��~��DXi\�s@1L�{��Yg�Žv4�$��&�~u�+�a�]Qb�E~��k=ϑ���ť#rYR�P1b��ԖO�����1T���V��
2�� 3�6�l��N|-���c�`��F�;$�$���$��yV*/�ȵ��Qb���>�ʣK�+9Agl����+������Rn�mέ뼷�����H��5�I#a�)46i��2�./DbOMUl�֪�x��8C$���'� |�Y�t|u�����w0}����U�Ő�a��������ZC�ݳ�>g�u?���i{��Y�l���@��D���%�����l�ɬ+�5_C뷚@Su��e`8s)��)F�����	n<� 
b ^�[��}�lP��T���%=2	�I�%aTk��P�O+dpx�u6�|�ٮ.��.Q��Lɢ�݇,�H�ȼ�����w����j4H�1[�&��\_��J:5Ϫ02<48�Ƌ/Ak逸���rp1���~��h.��w����^?��f�uR�H�����[�Ӟ��4h�q�:O+1w��9�j�6�-��!]�]�����R)$JG%q��A�WɔK�A�p�~��[�<���n�0�|�I'��lY�D�'���������|���Tu�-\��� U.=*%f��wm�Q���S�Ӱ�[m�+�.��t�$s���1;}}g�y���O?W�GhTG�/^��v�3�8cl�r�Wv������Y12���us$ \!���n�Bv���:��v0�.Y��-/��R{C��QC���E�&'�3� �(�����%�v���ϴ�s_+:'�4% ��6-2U��pSF^&��Z����$�std1[0�<�afϨ��˓���h�A���/(��T��)5��gi(!E^M��Z��l��ע� 
C�2�"͆�v�mcbb���>��3�WA��r�ʑ�^:g���h��X�p��l��1�p�|���ytSS34M��)	y�^ѥ7���A^�,D�uը6jA��ɣ�NL�t[_�{&���5�$�U�1Ә?D�[_���?�j��q��PS�?��x[D+�ľ�*���
9=�Psu�l����\�#�~�[h7�(�z���d��Jc�0�x�9�Ȁ+��5$Z$մM�g��44&-���r!b�~���� �j3Ǻ^p�	d�\��Q[,�5lL��2�	�t/<�~�R%l�m:94$��n��X*:E�X��HT���|/[4��GB��Pg��9���0�g����LOE.;�E��Pz���3۷o�o�P�Wj?�i�>�ѺA��Lu��-�ioo?��ə�k���-�ӓT�/_�G ��k����?Nk�����T6�78h�UP�=u�0��%=@�A�E�NZ�m�4)������}v٭6z<�)�"�~o ��*%ø{AnW��6�rѱ�����_���/�Z�ᢋ.RS���.҆�۬k.TA��]����x��tA$�yJ��k'Ȓ��������]�e��K�����������w.Z���iu�������%'�c���]�?��НGH��+����ݺq��p�?����^v�hE �T@����J�G����G:HZ�-�u2�A��#�ho0�ts�'R�$a������'n0TN�Ga�Ҳ��w��������֬�����ńe�H1�f#"C�+H��G��<u �`,��J"�0	`��rQ
���pm��o}�g?����7y�k�=��Su���%*Y��޽�?��?/�����^|H)�V�-1�w�w*� 6��6��V_L٬#�K��������A}L۲�͂�+a����4�LF�@d�F�踜L@��$z��f16֍T����I95V��/I�B�����j�����?[��Q���{�Ђ��Vt�p ���<UE<"�8Y��2񣈶�@7Yfs�n�����]bY*�,� ���=Vl�8�?���� ��_��e/��ۛ�+d�#���D���hG �("MF.��D�!B��Tr�P�,�ݗ������軄c57U�왖�Я��c�*<�jk��Ȥ��Z��|���[9Ĝ���  	��`��v�ݙ&��펞P�D�h1�s'�c�)=��h���_�/"�X�tK�]�-FV �`4V��YGo4??���ݣccc����Q 'idd�/ U��Tcփ;vHE�&�))0���f��c]� �����4���G� �T)�G��֧�z��oڴIQ��tˡ������k��/ M��a~)���pI7�Y<��יۇ;��QF���=̗e���ff�%�f�uF��[K�qI���d���" ����Z#R�48y�T�P�  b[�})�v����0΢H�'Ī�i�uGs���KR#�_���EYIG�"����O���`tQ����o�A8�<1�����1ϓ���Nv>�|!�Z�����N�V6�֡R�`fxґ�dFir�֬Ys�'"��=3�l-�,N��X��%'F˞F��!Hh+����o	�I׊ׄ/XX���|�������"�I�"v\ѕ� ��Aй�S�$�]z���R�B�qzG�ⲹ
3�)��1�I&���T:�����"���T��nIB�>X�K�o��b���ŎE&Ȑ~Ap�j���386�N��75?�u��y����i����b_�9CI�Ѡѹ��0X�t�i�?4H��ݻwg�5n���6=C��+�r{*Z	8?��:�-�!�@�js5xhM7~vfN�����k��u׮]K����{av�ޥ8X���������'�Յ%��-*Rkb�6Zr^H^���it��?f�JX0f����ַ���׽�]�z�i����_����|�(�]0_mI���"��uD����ƂG�wTf+JF�f�~p
���z��߸y��7^��?��e��t\~��_��Wɛ��UW������?��O|�����l���d��}�{$���{���ߏM&�+C�����H�oS�1�ؔ$�|%)��P�<�wڡ����P�1{�����'Ƨ��_y啿�[�ȟr�)��ŖB�M�Ĳ�V�Z���\K�]Ij�q,�v;���󣣨Y����)� ��M���{���s�y�\�מ����4L����?������+�&��ĮVp^8/*����F��1�������%_�y�3צf����[�`�������j*�
�$UQm�,㖮�0y5Rb�[��(1L}�#kI-����nEq`� X筘�m�`��ػb7H�"�䵲�t,4VG�2&��0=ό�w%לv�Y�_Q���tK2�TM�L�:��
�-���!eRT!'�B�a��E�����d��v�g[ܯfڅ�7�n1L"���$���ڑh>\삳э���
�m>�57���0[���^
����U�W�e�Je�,���g���ZS��'�O8�w�������[�n���Ν;S�!��)8w\GQS�|\�f����
E�gK�)R��YH���������T\�z�4"v��?�K�]B�����qy(�����&����)^���E,@h�%���r�����L���D�Ԇe�1��S��2c��=&�m,T�+��D.I(�H���j~~Qy���W�gʭM���'�T�/���V��* ,�x�d��$+�8��6Ds�������j��*��07X߅R�����ڜo��~�0$�ԍe�h�i6��0Lf���;w�=�h�E+��޽��@6�2����W��~�Rn���N�{5t��*sT�&��u���D�)EG�z�J�d[Ae��իI�U��9���dh6Z}n��d�?�����w�O���5O�&&&���b �n��,�Y���e"�QV�^m[썤�X9�9�0�3�,}�h��z�WI��R7Hɶ2b@�S���nKZ<F�E7rt̴�CBb�#3;C!�֕�V�N&l�Q��,�����L9j�8J��0#oh���'�޿R)*��x"�� aACit&x�a䭟u'�ت)W���"�B̌L2��O�ہ�Az5���>9��#W�a@���[��r��s��$��k, �o��V��+x�̣T!��O�ī{n�4�W�J`,p�qZ��p���G�������ٷ|����M�TK��{T[i�� 8ס�2�-kJ�0H�4ݑ~�Lt�~�X�H���ߟjցjdi�lӁ�'�F�\O���2 �cd��,T1�\%�H�|�ŤS�Gr
��4�_*��w���e����w����׾������������_ЪX�z��M��{�}۶m����g��J��~����kל��׈L#��+���/��H�\�L-G��r�
�&/�$5��N�S��9d�����&�k���ra�T�芶Z�5�!�&��(;����v�$?g*@�k��E�� my�F���T;�D"�d���SS'�|��A�R�q˭A�]��ߦ-���<x��k���C�/<a�M�b�C�����?� qt۵?�l��n�n��2¬K~�u�f'��t��g�u�u�]��W_��}wWJA�L�I6w��ٿ��g>����
�\g���h1d���Тbʦ$Ӏ4B����A�^}�m��t�+�����6�0�:IU|��S�_.����M@����������,^4�$X
4'�t��?�a�Bfl=aÆ�w���C*��[�Ȕ�m���-�����d��G�a��YI���J�1*F�}�ɉ�Z̨�鋯x�+�l��W���G��HL�w����Ţ4?�����	� �1Tt�2�v�)J�Y	Rbk�k%(��h
�W��i�Ï��|Ҧ�n�ᕯ<��kJΩDa|/�yiZ���.y�;IP�i�#�ȵj�� ��.#+�Z�4��b?^��o�ۦn$�p�� ŰW<�	�m�j`�����c����qW�<h��VC5HP����z����|'����(���������䔚y��xY��%���)������D�����y,<`���\����~�%���o��4������'�t�W��5��P��v�Ύ�_����G���I'�t�/�;�O��?c^����7�8*����,���-�X�ݐV�[�C��kU�7=Za��yȀX�ti�"�9�F�X@5���ԝ�w%S�YG��U�%u��\fLiF��7֏�i��;}j'���M2lg��PA���pqʬe�%�k�tu�(��%7e�ܸ"�gvm��	8y��C�)�����z�G�8@��ԁd��: ;֬Y�2�ʹ��Ii�vh24�<�a|�	ь�Qi�pj�3$���s�m��t	Y=H�~ooexŚ�k�.^��Z���k׮�j�;
�Ӽ"WW�[�"xqf�P�5��.�6�'ƝiJ�W��>�� ���Y�dI[x=C�@h����C�CV,��t�z�L�
�\(y�1���@E�=��4ϽHSY�����1p5���;R(K�"��j�PX"�;�雨�eeA���<��$BA �	$��H(
�1���K�0SR�J�LN�+G��5Ӳ5�d����q�y�]m��7{ofI]��k�:[�޷��Y�a�fXE���"q#�#�r㗛�x�<��3�1C���jn�P"�J`d���a����}9}���{���3K�����PO�s�N�}���]~oj�J�I��=���$˕��,ƣ�`Sj��zF��ki�rX6����y�h+�p�"�u6jX��)���ݰ\�}�P���m��� $�m��.�j`l!S����,-�#��XK�� ��O��{9��#��D�����KM؁��d�=�梁t\�:E�S5��|��5���)���}�JF�^��d'�G�)����꭮7����o�ʕ�w��@=�.G�f͚��c�����2U��і��&�iwO������g��aBH^���������ރDا�!�l13!�<��oA�!�����@ga³��[��<�-"qۦ��QD��9C�Ymф��0)��puM8�a@��˗/��eC*�D�ц�-Da����
� !IDz��R?��m��J|W>8����]d��E�k����moQ��SO�:oyM��O��O���������7���I
5J�c�3��(�T+��;�O?���?��W��I�8y۱���w�~Ǐ�!e�[�Uw�Y���;����V$T�.���;�`E�Z���'$*~_�5��䁩�C�qiKr3�b!,��z�RQ�jw,�Rє����Ŧ$̨	e�M4߆k[�C7o������?��sΆ��UY���?�W����;>�!E"<�	as�ŪЛ��x/��QYС�w�Yg�n��O~��>��Q�mn��}������m��Qa GZ`����>�M����7���~�J(9��R6@����w@`�|�[�h�{˓�6mhC
A��.���楗^��?G~�@��۷\�����~��T-�W@퍰𹒂"F\�	%ʁ��xS�^4��Ŀ�Z8�f���7 ��W8�sOY|�D��n��8�vᖆ�Ѣ�겢�۰d�h�����O=~��3-Kq�5Pu�((�f��eI�����+���wE������y�8�x�u6�ڡ�'��?���^~�j79�r�X�T̎*�B��6��+Ɖ+O�^����ή©���{��Yh�:}���{GF�G��a<J���]�k������!��)aY��������SL���~�T)3c[��7��Oq�@� C�`̘�@�}�hD@��ju�|�ij(i���[�1%k"F[[;,��	D;���uE��|�"9O�1�$%<��[Z��dL��1��E��$	��N�l�����5t�X&z9��tvv�ڱ��alI���ͷ�����oA�:>Y�u�7<K�T���n�U��,?������ټ[����2��]���w#�ް�0�j����i.f�=U�B��(b��<2n���:thZ�?�����K bm���{nd׮���|�mm��S0�=-���=������t�:�%��&DYZ���`SUԞ�bVV*�`�Tp/_���]5�,����B���ڰa��с�v�Jպu� �ˆ��~�y}���[o�uf��)�|f3�!5�����D���LLL��Xf&���$>�a����j �~59FE�[������n^	�J�ʣ��(��)
�;�݈�댌�
`������� �<1"�=H�M�7�C/Z>dU�����]a���Y�6��c�"ǝ�6/���ۥ8I=Z�z�c�hg5��@X{�����Q)�V�\��`��ڼUdYjkk�����b�z�k���?��]�����XwG���J	��3�	V��ԣ��غ��3��j���p|�+��r1�A�������s�7�^�Nbt2�i���ĈǶ,b˭��]��cS.r��*vc�lO�f��-��,V�=cc~&�Z-e��2�����Ѣ����KVt?�/���D^���\�0�d��,�%Y�[��U��\�бb���U��go��Ʌ9 	ӍJU�������\�^u�Uk�m����<��s����P~������'W|�ߛ��9��s�8�w��=��t7p���<Xq�����Re��U�M�`��J�9T$��p���W�@))vD������.:�h%�0lT|�a�coT�C��^u]��J�8��r�k@�,"�L[QDՁ��Z�sժU+�-[�re�,_��<�pjn�Ț;��D����:88�,��ӟ�jt��ן�����e[�ly`�C�\r���'8rd�de��t�+�����t���#Qx��6�H05@݆�������!d7О�j���نkĥH=郗_~���ba	@��?���!eD��Q�X9m�K/(���N,Na06~��xӗ�|sŌй�b	-_T�W�D�Ȩd������U)��R��@��BNk�uԎ�S"�h�GK�yM]f���ZD�z2�(��=Hl=V�H�[��f�2V��l#��4Z!�:)��/�U�`a�f�6m�T�#�nx²
��F)ceT!9vM��]}���^�
ǋ��R�h�9���s��bP�v*�u�����~�����Efx*�2'.�.`4�"Ys@}U%V]���k��Z��縎�zEs�,ı���~���^��#_��f�"���[A!�]���n��n�;h���6"���SS2Y�0���ko�̧?�:h�ʘ�_��H��	��S��K��*��R�&����l_��f2��_�]�̠����h:[ј3È����Y�h�Ѕi���$S��FG�Q4Ox_��W�{�9�u Z\�N��!s�&�x���s�d����|[����p�_������۶���������$n���jYDQ�QLQ�č!(�mu\�UF
�b������?���#�g��K{A�Im�N�R�XZ��@�a����6�p����L���I��=�qf�U҉QVe%�iZq�?RU�d-�TN�`��n��uH
z̎͘?5�%#��>v(q��M���BC��m�%>!�S�ۼ�3���𜎎ÕDcU)��6���bOa���[���Թ�Y���m����v(�ޘ���y�D�'*A5���aa�z{{�9LyY�B��iA�,2k >s���$t�Y*�]��
J������f�Hh�D�㖣�<�='H+W��+�TV����H��t��.dk�	��4�3�#	ݰ�t��:>�sRph�ʘ�]�@�D�	E��'h�򣍆DɄ�B�4ҏ(Ӣ���bh�(���m���U^{��H�o6�E`TU��
�)NY����*9~�(��*��N�J�^�m��"A}Q��E���,'h�(!��4��.7����Iuzd�� �EE9����D�\^�T*��l�Z�x��"RE̗a�b��^�����!'@�j.Wk~#�<��@�ecp�}#y9Om\�.%��#�Yx�~�Fd�����3j��z�a��LS�wd/�2�bV�O6���i�:L�,\�1�dؼf+�z�12g��a�@`�.t����?R[�٥F��'5%%��Ô�~�A`�ڵ��sυц��Ll�HL���A�h��O�/��6��h�K�h�2Il� �6&�/i�P;�ǹm�����[Ck:e(x!���X��b�� �"��hZ��g �;����J�G�X�9j�h(;�5��)[y+�w`�I��ͤ+Yb֗_�J�=�tX���ǒ]t�Y�'l�q�0���U�3C?��(�,���x���<$�0܃�� Dwheĩ\HPF�ue�^���Җ.˰��?�@�2�7��8�~Q�c��dЇ#�Зd���7R��ϋ�gE�<�W�*u�5�Db�'�>!L�q$���|I\�5�%�To�����`�9z'.u��
R}Nj[��z��aZ��1�CQ��=�CC1@!^Z��E+'��q��r�Ij�������Q���h�t��d������EQc�i�$�����*�`���&|�zuC��v�=��J}߇.�����'&N���Sх���[�ǧ.��}ﻰt&<�Ӿ�_:���9ﴍ��En]�Z�H~���&H:���ąŻ�M�m�:F�$�����`)����h���1yh⫥B%��<=Ŋd7� @6�ᔻ���^:��5�$�������أ�|�o��m>m�#S�6W�r�韾�����������&�16u$V��x��^��ż�M�9��`�毠�"_,�la="�����.[���_�r��3�<s�)k@ܯ[�n���[�<�َ&æq~� ��V]̂ԓ5���Lxck�`��b���f�0�,�B��Q���,d9�tC���U�B;$џϘn���ض0ߣЃ�=�b���3s��.[�,/��E+���V�Bn���b:�dL�B��� ���H���7�u�� ��L�#�=���7�ֲFz�a�
��X��U����|�f��Н�<��c��z;�į�ʶ��]�0J�R�,Cr�l�$kn�.�JE6ZC-�-%2�Z`�]��F�-W(W%���a�ּOa�X*CR$_��AE�4�QNJ]��f���S�,[9�����ԣ����h���mX,/���Δjc��nP%#_h��c���x:i�fم�%����hA{On����4�Z�gׅf1JӮ������Q�Zs��[S�0��g�c#Ƴ
9P(U�V��Bm�K:#�&�0���OLL��ߖb��$�`�0����A�Ga�c]�l�		��i	q^h��#�4��)���'����!ͱ�RB�E�a�F0@��m��Ut�BC@5��T*��,S�F���y�6�+�tt�)��"5��l4��I�A�e�9]?�J���m�z��r�
;��bŪ�O?���k<����GTb����e����h�M;bj0v{�,;�]����Cj��Mue�A�_�^G�
}��DU��8yE皕;GvT�����0*�Q�称ro�;���|x�~���?P��^>�l������A\ ~	k�V�
�R�W��lK��Q(��J���C+f$�$�G����������x ��ζ���a��ݿ�'AITt8�DK{[W���������6���Nرs��b���[$��Z�>$)��a5ǭW�:���]�����SZs�C�����r	Ƥ���������)��p\�8ub��`����G�� V0VH9+�P�q>@�j�b
!E��n�R�� �[;ZaMW��2�R:
i�J�'�X	�Ĥ�ڂd'VL�� ��C��hG�0��HH���K���4�dE�0$���uߝY\h��*��T�j�uˎ�5ܶBkyq�45��&;�����_1�I	|d2
p�^�*r7����OW�˝�M�)O��zp8QN@�����f�t�
J��42\b�O��~X�BP6
��}���j2����E5;ѫ�P�:�?�k,��JC�#��C�` z$i2��ng��f�!��	k22�B�K'ݒYs)�g�"z���R�3��!gs���*��1�W�,G	���4���}R�'_ ~h^V��f+DvXg"&4<�S`�-ŏ|��&��D���S�ʊ֜�A!��}8#���SX�F�@*/��汇*V������!e^ �{�KYCKˊ��I���a�F�z���Z�r�����l�X��u8�~���.r�W�டlٲ��}�'b .����?��r���7�������S1<<|Ά�H5��q}c���+z��Z�f-!��cr.����{�{���-^t���'>�1�~��Ȉi�S�n��;`��O�$Q\�hV!;���_뭷�t�I���i��{�\��%��q/%�)AET*�=���� ����E荁�v544ρ��F��H��l��`��P���l����7��Sw%�ΰ���!_+�>�p�����p�r g�yI����'��R��e޽{�ކ|����{��ǱU�U�
0�!�;+%�]���N��Z�E.1$Q}� .ݣ�I��O�O�m�*@�,�&��5�\}߸r�>��~����r��I$�����%
#o�$� �2q�)ĳGye�����s��v������y��yS�9��H�H��|�H��գh||��S��YL��H]����-��s�ʞ={�a��?�{�a|�>z�����_#�~-��܎�ZH�fTd����� =��r��5k������ر�G9p����`i-T�аPV �岭��{laAJ:�J�����̯�8�O?�4��V�S��C�����L������������6őZ_	��;��Wq����uC�`�uKl9L�p)k�a��b����\D�g ���ٟ"@��}t�]H�٬��H��m�IZB�,"��54�)ix�JE�*��$|�N`���2,����Ӣ$�����;�7��l%9��HH�4*�k���n@���
6����]%�#���Fp�y�wN�tG�Ӏ�R�[i���3"K�*��kժU=CC�����qZ������C�P�������H�<&��������5 X��p?4��I���G�Y��O���"1�WC��s��M���m۶u��{��Xh34~��Ֆ'mݺ�Ћ/�/N��+y�a��R�e����q^���?��Oê>s��7n����&�g�B�T��Sx�x�f1�EhT���*��=b�Щë:���l�]U���p3R��}�v���]�՚і���
�k(Xf��O�(#���.�sss�RD͆S����Cc8WF���6�E�ZqŊ�_|�T]���wuu!���EH)%�D�|ίq%�+�b��(q���H>����_�>{친Z}����ҷ�h�%�߰&�����WS���Djʉh�*" r�ə&�4[��6�_㊁�N�X��"!���vzlk�kYK?ga+�G0L.5���&ş}5��~��7�֫\��V�U|��[~4:[��.9�ܷ��l��K7�=���S�eݔE����!7w�։'C�����B�0u4((��ZC!��x���k\Ǯuq�B|�ź�
pZK�D�SlϵL#m����<�j��������u�O>�η�p�1m'��2�M���R��@À��q�Աr��C�Fze���Qk��N�xEX�9 �8���W�7�T1�x��ɉ�,�0�����c->��uFf��� [g�'��Y����|����ʚTa��D)/��˶�VfH��,a�$�i�* ˅ߐ���� �W2�^��\	�&&&+��s��;:�g����~�����߿bf+f�h%v�X�QB��Id�j(��v<�j�z ��(�dM23���(�M���j�`�5����E^ ���#� -0r��H� /�`�U٩�G���,�����uQ������e�7a��3>S���Z�MW^#�{�nX��ٲ�cЂ��̗F�����%p�*t!*��䶶ZF{�m���ibTT��<���%��0a�k Y��N�s�ľ�N37`�dzZgFǇu�h����Z"�3�99�ĉi|�˪ͬx�[5SU��:��D��X�%#�U,`F~��а���Ov_?(��9d�X������_���ʖ���ޞ}#��ՊD{ͣ�Ѹ��8�)�
���t���:�wl�0LT���X��յ2�I&�w@��$�4s�%Z�#��q�V�a,�#���Ϡ�p��1H��T i��Y��Q��%��jq �h���^�(	��� �#�(M�`�F��C��>Q�$���_C�|��\�1�ZE� �HW�\�Є�>����t���	h��͛ Ϝ�a=R��k0S]v���vG#�\���\������N��32Zr�֯�n~��� ��5�{t~��yR���_W���r�[�����q��+=�e#�"��U�I����{�ɭ=UC/�a��z#����ǆG�r��������4ǔ�����]s�s���r��.�aN�X��g�+X�-��#��s��
����^�F</���e��33�u���zhh����dǯ����MC흚���ʁ�;���҈'�5�*���s-D� u�&Fa�k}�ZX>Xwnt��.L���38��X���2t�'�a�-X	f�&C�
�I�$��	����G �?"�
$���<عg�ў(َ�X�
B�Q٪��f	�[2�����m���=�6N�,�T�e��\$���d#(g��N���a�\6@8j��y��"�2��M���`��Sc���]}م�:��Bˡ�ѱ��Suu`Պ�����g�g/N\��*9���/��tx������&! ǉ�K�6IKP�q	{.�x1��
�;
)H��D���=+m�8/�~W��f˱���#5v#R`�G��$|�qK���BjB}�.I�EA�X���a(ѩ�R9�U�X\43	5���s�q�f/�[f�����H
iIᏈ�"��i���0�U*4�8z�RبF5�Bu1�:�����p�%��d��zDèO�o_�c(%	U��������D�(4��h�����s�Ɉ���*W��"�ɵV��8ѯ��\μ�⋿��o�رEߣқ�1uP�1� c���j˖?��?Z}�y��{��4��:��ԯu�F�k*�}�+��׸0��󱈥F������������K�\�-���4tEٺu���	x���M `���:Y�`�ێ�+�x�������l��<�(�{�'�tB��
�k�u@���A�M-�����ջlÆV^G;���+	EƸ������=è8s���<&%i-�>��j)���:�W�Z���7 Ђ	m��g��z�3�^�������F6�lٲ�~������^�����R[�n\�6��u�B#}a)K�k%I�4C!�?>Sc:� JJ{�^�옂�s�q��6���0t��O�-�87mڴ��0����J��� #,���!����0�F��� ?�
 ϓO>���hٵ�\�[$	�<��*�fff����z�[���[�ώlhZV7�{��/w��=����Ç��#�� 9u�!�a�dq�V�t�;8"[��(iB������Y
p���m{Jń��e����2�ɽ�K��ַ���-Vo����bF��M�ӡZ̚���pe�G���e᱘d��NX��9Ūa� ���^o�_c�4b+e\�bq�����6�(�8M����	�q��gc~H)q�%i`-&R�*T�F�"��F	WK�h�N��b�sz�8R��f�'��̕�~|p$Wa�{�>-u,㨺��w �,���N\��Z�Y�,Z���Ꮜ���{�.�˓����Bgg'LPooog���i�ӔSD�eLy'ˀd�<���'a�~�?D�EfE���=+1۪aEr�"��KZ�OZ#֎Դ����(ȵ���F����E�^��$���v�i�ׂ��3�{� �j(:^|�ŝ;w��؋Q���K����q�lY+����@U��գ�{�(0~����O>��od�y���a�²��:�� �J7Z�r%�����Yg�u�.h�7� H��o�_ټy��W��-�����0���%�w�B8<�t�K'�(�Y�>'���Aڷo��@ll;�H\�~}GGG>���U��_}jz�+�E�CA�~)�*�,5�:t���mP�?C�`_g��O�1A�2� s�<�mw;2��qŊ�����}�ݷ��3�<�s�m�6h|�f͚�GGG��m�s�2�b
�x#��B���5��3cCk�������k��vq>��fL[E1�"�V~���ĈҼ����G5,Jw��sG���4�k	�-y�^�!q2=�d�F	)���}\��y��)'ִ���K���*�ף����!eӇ��(��7�֫\���U����.���b�УϾ��wtu����{��/_��]?�g��S�Hd,C�|7
�Vd�w���뮻ޔ�)N����M�QFW1�VUj�������P��{����C�T)��(0�rʪ�7��믺���S���j�
U݉$#p3:f��~ls#�� �j���L�P����#ņ����y����r�w�"�IµL��4�r��RUV8�As�ԍ
f��b���/��* v5s��Q� 	l߹��ړVM3�����/k��*z��̌ �X�*#��dr=�-]�����W��?�����x:�z���[O?�{�.�d��}����mm�p�*��-��:�`�0�����T�:���O�*&�R0	�Y��%*P+ZZZ�r4��C��!Y
� -��&]? p)R��թ�Ƭ�({饗�/_~٥��ڝS3�総�Z�j��G���>������۷��Ԑ!�;tH��#���@Os��l��j*Qi1��.iAOY��;���B��J��6ܲ���"��c40�Qʙ�,lٯ֫Y�u��`��/<��kQ?�/uw̙j��o��)��[ֹz��y��rev�����E��D�5o�r�n�.�BE�U��#<wa� t�H���"o�O[�-���=�xc�H~���V#�kษ��jZK�\
ed$cF�lFf.��'d�.`VtL�Git(�І��y�T6��j��O�����\5Ѩ��q/G�G9��s���dU��$@�؛�P�\�(�X��r �6�y�(r��z�,��57�ԅ��_��_�\iK�&�T���1.�T(IYگ���� 2��H��eMKQ4�i,�����w1&�����<z��ځ��vPV�]C�s�����2AnT+�KU�0��Q�? S�)r�m�b���;���].XVC�?1��V�޾���Ź�y��[�q~)��5�U�>	;p��J�/��Zs�{mb���bW*���7#[]��55lk͘�1��Vrj�8h�/[�}q�3OuJ��d�nM3����F�]�fMk�e_k������櫈�!��f�����x�)�o?�Ó{�������/�Ȕ�`f�BP:~�z᪾��B�������Ryd�N�v/y��h��c��<v�C=Vvm���I�Sթ:��	�����4KA(c
'H',�7�w�h_&_��˱_�&1��BT\-��Q|[������������@nff���	��������m�̆�B��!\�~�T�L [��dA�_����=��=P4/�ɕv��9XIOҔF�����B����xa��a�f�gg��٩��q�H��톷X�ſ>4}��vh^�}����r�&d�$5���y����~<B�&��"�}K[s)rLpi������A�BIJ(f�K�f�ݚ
L�VR��@�-/���j"��\����d�k�Z�xJ�Q���e�7z^΀�|O�5:�ău�[��.	:	0�
-3"d�EުĴ%�}�g��5�r��j:Q�GJ<u�W-�&�/0��Z�?����R���[�X^B��|��׏�����Z�r9D֤��h�����T�+����Z��~�������/]w�uC�*�F!�1F&��xc$ύ�����s�}�G@Σ�%(��Y,�k��W��Q�w����}C��uJ��	Y�������/|����Y��w�g�2x�*Q}d��d����G���N��	�H��RA)^m<9ꚩ&Ӹ�˴��T`�g-(O����p
�q������������(t-�O����䲀
 r �aن'b�M�����!�A_D�4@K^�j��Z��+TÝ;wr
賳�����o]y�w�w�޽{}/�&�cGGGEy!=8߃r=��e2o��%�5G�KɸaDq|�uLQ�(�%�������Lr,5�Lm�_�~��_>���]��?MR<���)K7���ɩ`
�,�Zؒ�����>��/�JKd��h��0�r������tF���3�t���2��Dp�W#��u��<��suŊ'�pjr'1I��n�g�+`���_xᅮz#�˸UĮ�}���L>()g��B�t~(dQVLb�q7�>5`-h�U�b�F[�K����R�����g��)��y)�0V���,�r��k.�A�v��/��0s���ZjLZȳ��Y7vr����bM�$�c>��I�C���c�H�$�0�_D�q@`GG�vZHׅ��s������fԪC�9���v�4��<�*%�͍��=6'7��������R<W&�Bi�ՙd�I-~2�	�b�
��=�1վ�>�z����-����0����sB_7`��"C�{<�����ܓ��6m�}���lC�Z�8e6�~�q�"s`)RY�74|����䓰"�����7Kr��G��,�sdx�4�U�h�F��l���w`�� �a~r�  $���dC!�d��|v.�ս�ދ{G�9��8���eԂ���O?���|  ��	��[o������f:ݶmH�8$��������C��>�,�2�)Z,Zp"�|a��16QY�ᯝ�݈�	�T�-��B+�u�x?6X8.�ZMBW�,`O5��l#]/�:�0������a`@FF�Ͼ��'�|������Y��zV��"4g�=��8�/���MMM��f?31���ӱox����Y�����Hp)[�ȳA���a�P���+ڠw���^�� C���;��h�bug���q�W"qT�N�:��}�Q�$���Z�����O�,�r+��q5���r\3w�7�٩4��MU����������3Q�SN��c{ެ�4A��.�~}p��K�F���������G�^��xk��j�jh�3��V��W�)�hy����
�V���w|����`��n�
٢SEU�����+��"k���[߼���+>|�mߵk���Ѓ�Ѳ����e`~�k��#$74R}Pg5��i��*�~�u��'_����|�c�HoDd��)��rף�k�FK� �����3�L��U��=,=������>�b����s���v8�A�ǠoJQ'۪H����J���<�����|^�T&u�$E�}�&���:�ޮ>euwww[踒i��J����Y2�	 �&2p���T�1����ԡ���b��53�����}����u�iz��\��uk��t��b��V,7@�2���X�����)�ȸ���jk�?�%5r/aS�"�&�LKddpm��S�'�򉋀�p#�#Z55E�5�@Dm�2�.y�;�-%}k]�=�[<�Ҏ��������h��2й�rԤ�A�m>� �$�)�Z�Ĭ�5����Yɑ�:V!�5��6::"Iu/ͬ�68�w���8lUC����l	��l5��"�.�������Ng4���/o�����N�+��j0S���c��ٙ�9ea>rC7*@�P�r�jc-����v�ֆ�b"��#v�ְz�!g�/�@�Owm�̬�b~Vȩ���1y豭�F��z������y12
�%WUf�qxz�(�)YZ"���[\���yh��,��9N�A�{�u�D��%�Z%��%�R�8�0	Ó�@A"Gv5MA-���>
��>�YSU��{���b�ʹT���IX
Y�Y+�A��1���jM3DI`��K�ެ`0Xrq� �lh!J���:�h���a���`�����au�.,,NLLZ+3��Hrn
�\mذapp��0}Z� �?��կ��#3IȊ��!��bx'FL!���X-� ���\�S�n��ۗ�����b�T*-��Z@�f����L#��hohm�b@K2Jef~~f�pn�2���jlC���O��zF�����A#"d>Az�،[��� �������}�Vq0D����0ĒUH���1R�-�x^ rS]�ف���>QA6����7#���S>aE=��m�t�����Z��0���?$�hu�50�5��Y�&d���F��}	����b��l��:g��������׹j�ƍ�Z��֬>&���C kO8c�ǆ'����Y7�-ٕ=3�-U�ja (7B�g�*�ttú5�����7������ D͕K�'�|��w:�|���{�'~���j�z{����Q)���P2D��`�<�m�����q��}='r��T��m�4<���v2;��"�e��],~�+ޓ!#�(v��X׏�
�1��X�H鍉�8莬*QLWC���|)T�6=ū3v�0�@r�~h��9v1��*���D�PJ8�pҭi*Hj����N�����gS<�ri4����t^�c�VER�0L&'�,D���Г�x��C��P��S꒢��������=f@I4x��xj��]D.��Y����f�K#,q�,y�9"�a[jr��T���z}(��/�#���bǳϗJ՚+���*X�>�9x�*֗����^�~M�3V�R��6���P��x�G>���z����]hkkuº.cT��tի_GmT�#���Y��@�%������u�)�z�y�x�;����n��sX��rުU��{׻.��,UY,��u����/�޽���)>������� �^a���1(j+�bEM$�(@��\����?�P$�E���Õr��h���/� ���ʞe˖�mkk��z�.\�P�A
b�[ZZ��*h��Ź�^zi�����:��=��Ӡ!u����桡�}Q;��ȡgesX�%�Hr\�x��'4�G��Lqz0�c���3=�\>�y��t-4.c%�����y��,����=�br�٘+]�nE+�A�*eX������=����}!�>���rh�6q�*V�QH��>{����mjV<Vُh'�aT'w�����H�TY��4���l������\,���'|���`��͛7cZZ�X���j)S����*�R����.����@e7*���Xm�qɛ�PH��;�#��ʩ��=U^��~�:�[�CC���I��_|q����3Ϝ�]��׿>7_����ڸ�"9�=��Gp��:j�sv�0�@r�}g*F^<<�<wE��*��%!�����#NB8���}��U��qJ�$ø�A�,�:`����>���<�-'5��]�Z�ӎ�a�ёu���6U=���t-q�!�>������T�4�q��\����~��SV�PZ�V��a�%lF��@n�m��J��L��m�s�����Hh�K�;�qw�J�*�����Z�A��x������ )=N�C2����z��Z"���b�XD=�u��09���޽{���ǰRwG� k�'�<��T�.,��o�;��ւ�����*�҈i^�aK�+�B"A�`?-���(��rH�~SU"��YG6����&Ơr���~Q�r���bԟJ�'1^�fs�H��1��Ri5��E,�a쫗��:�O�z�f ��g�0,ڻ��8?=7t�w�8��`������i��m��P���x�G{�s�<��j�j�I �?��OcvV+�3Ș7o۶m��I0�'D�~ɍ4M�# ��A'��9@W�aN�ؗ�e9�9fS�q�lD�BB�(�]����:���;�焢Β|!I��9�ᱷ�����qd%qD,�k�Lx�E��FOJ����,Ux<n�cu��Oq�먗J�R�X�蓅KNPӑ�Q|��#�W���!Ɠ�|��5�^(��7��+]8�J�	<+�2Z���
�l��nD��ژ�@�������m��N��~>�c�S]�m�P9uG��U�}���b�8Q��̪�HJ�7�T�#9"� N����?�	7��T�ې���ʛ����$'��-ȔI!|R�@��a
�Ѡ'�.��-�,8�-W�׾�7m���?�����fdY��?��?��_���|��K�H���EA[���������?󙎮!��)���GĎ����a��\�X&��`SU|g��=$�B
I5�T�>���H���E`�PG��f��8�:^F
�>Ɖ�7�y��++��b���Z����G�.6"�PPx�ȶhQ�Ty�W[�n�
����mG`�e:��{0�\0��^h+X�Fm~Ϯ]�
b��c��^苪�ʘ� ���l��q�]��D���M?0dː=M���4�V��?�/�^��Qg[Wְ"/�,���7�I�"Y��
�C3d��UZ����QZ�Y��m�4��=���c��r�\����o�hW����Ϸ�����jYO�S��U���G��6���dP++)c���z�gT�pq�����$���B�Fׂ����\��R�V���"f���^(L�f�vU�e�����X�(�|����J锓םp��w_vY���R$�diDs��眼n�zд��yhU>������Cdh�3���R������=H�����f4$�xd�BZ���~�W�@F�	,�3.$x�bA��:w�8��r�X���U�� 7<��Q�"C�����e�C��-mBF�k\q]	�-
�1+�ڙ��P+WKs�(���_]&� �&.����������a���7�(��o �Y�XrhꖈIh�⏌��煍�����@��h�;��0H��膢��hQ�DA� 쒾�:�Ҭ����b���뚎9����j�q�&��z2�z5�H����Q�Xe[���T2���	+�6��1k��w�����}{w;sX!@� eu:X���o���������Xb�e�E|Ґ�0ǚRff~1�ʠ�&׷ឧ��d�ŝg�q��7���͛AA/�����)\�<B�uP�m߾}b~l˖-��	�{$����V���"ZJ%�W�̖~�u�����C������RY|ہ��,�>ꁅ1����B�!Z%p�#s=Y��~�UH��5,�&�%��"p�}]2�|��6�2�̣jȳ��e�n`�2
�B΄��\�m�D����e�'�E�T��L�sK����(#��
 ���|�"U�64��պ�UW�)B��]0�O?�4���oy��==='�<�f͚��WN�whD7�����*>b�+5��==�=�-gm<US$��~��v�^���}�����(�����#���<묳")r��L����=S�l(EWQ,�0�C�ׇ}VtzV���j��K��"�p	&IÜm�\�P)�a2��~.)�>mj�G�������ʞ�-D�53�9����pI�w�t~6$8�t�1c�8"<)�����A*�Lē����<A�.���B-j(0�A(��^=l�
�e`�;N(;X�7p�*���E���G.�"०�XR���%�U��`;�����7�+�[�!G�s�+vr�;�RF���6���'%�B�̖��"�3��x��cu4��*�%t7�t���֊�F*.���5'P�Qœ}^��2Uŧ�*�óJ'��F�1��%W�6�(Ȇ��0�茐��l�E�h��@�q}�R[���r}@�X�NEo�������F%�"	O¾h�GN@;�Ƣ�7�֫_XI�G����GpZ<�륁e>��t�Ͽ|��p�}���M������w��|���9��q9�q�2F*��j �8RD��E�9��淧����AR�3E\�RR���E�#%�A\(�	.�(hç�I�0X��_Ԥ6�A���d�RH���2����Їn��w���V�8Q����/|�f��=���Mk�������}���\�ꫯ���N\ZtIId�h2)IKf�W�bc���
��erh�>,B�]Ek�mOMMU*�b�
\eq��RUb���A?����
�*Zm1a���%�����loo�]e~~�n,��D������a����ꃌjB|<�����F$���*;cz�Fu�$T�
��������诓�t��܅�
��覤G�z�����|Z��׵bŊ��^�`N=��b�8zpljj^j�oܸ��M����=��G_|��F��
�n# ���`s�X�*J��k;l���Iϋ�=kmmE�:��9�r�Ȳ��몋������}�0�T*��g2��0V���-:�6=|�X,b���l&�R�|_4�!_�4sןB������ݰ4�a�oCe������ �Fr �0�G�0��L�6={���Ow�Ċ@���Z�"(}�1�����a9N�ZXXh����|��ǎ�d�GQ�l%��P9�q�tR���B��3���2����>�g�9]$�����ᒹ*:&�y���K�i�U�D�I��,W#�0��x�{yO�D�ُ�����+4�2��'ǐ�<g�[ "��H劸~=:���B�rA����ny�X�0����,Z�лR#?	�t�%% B����>�3Xӵ�t���&��	��j����Z*���B&333h�aS�@%�nݺwn�g?��L��+eT��řJ��E�����o���!���pU�`�S��Z����	�yL�yT����Hm�o���,oc��Nd�OF���p�MAI���L����靴 ��^%���Xc�p�X��k� tvv�tu���n��`����XA�=��SЀs�L�f�`�����D�� TCa�D���h�B9WK�����w���h���l�R�d,Y�`�7�Y����d��~�\kģL����2�c̚�.G��� )�Ӧ��5���c68�ļ�k��5��M�*�LdK���Dɟd��KQ� �"K�	��=�GR&9��$� �@e�M���j�KsR�%x��t3M�pT'���:��!E�����'�*��Dr�"��g鸥�"Jb4B
�e"��:�q+I�,̗sG�zN$�͙R2u��LE�
|,�F��W)yc\k>��=��CCS���ab���Z�^��,�L�M�8
Q�F���o��6���'��a5:$�c�y8�x.�քE�C7�5)J��0�~��=�6X�ޗ�r� �dC1p2��6&3�^��X�.�P�,�a?������g@�a7@hHI%ɾ�9g[_��W>����k��=��ʗ������>��Jl��|�_��������	dXƕG��m5�����7l��h2������b�`P�k�` 7p�1��)K���NN���!�j�>��� ";�b- ����X`�H�b�"���������)ٶ�x�k����g?�k׮~����D�<?0�Y�0~�_-�ǃ`@�W�����e(R��d(	B�`�C���y��86 �UDX�J�_�\�0;�؂��V��������[�6�R���� �L��=B�G���+�v���6_?|h|���������\�{�:�B���Ԛ�y�z���L}QU�r���:"�X���X��^��B1�X���g%/2-�ŎS8*C���	!�$�m��r�蚤*��^��xt>��P���j�R��Y�re�8-ffCC,/#eĠM7@��3Y��4Ђ.Lt������S�����y����gm>5�Z���Wo~�5'���σ���=?{����,�v=�� �%ҕ9G��4����U³k#c�2���픧�z���Y0�)g<��zJ2��.{�/�٩����}�H��A+:��������{��^|��A͹���|���;��/9 oe���b5ޠ��
}���б�r�5�y>.9UD���N���N�)��R��a��d�O�~ v���w^{OדO>�{��R��j�]�M�8�\�q�vXm 7z.ۆu�T�r�؍�`@�����5k�ڶ��\�Wn��t���/�N�MXk�.%�>*RD��RIA*8��ިe��#c�Yww��s� ��s�ʣ���Q���%����$�d�HT�4��XRr�c$D��X��+9!����|��g�	kWI��8� ��m���=�����r@�?��������{�5+a�-�]����}���`��˻�S�v��
�
@b=��DÓí/<�
��8D�6>r�kΕ��`�jM��L6�����!x�R�a�9Mc��?�`���nh�p�n{��y��V�u]�uf�9�\v����S�����ఝ]w��0V|"�|@܉�*z��xTʽ����$QbE��.�p	93zDʥ��C�C5����ȓU���ق�S��
�0		a�8�48 =�db�^��6T/X:��ur��lYO������Y�q�# �&W�����vg?
���=e��l��o٧��J�` �Z����uh�w����l��R!�R��wYw��}:�֭�Jv�o��5'�,�{���%w�n��p�|h"B$��H.2m$*ks~A��s�J�eja�^nř<��(�2Nǆ76�i���Ҡ����k�����
l�H���߸���A*V*�|!z�o���gY�TT�8Z���gN�M ��xT�U�Nji�����r=� ���)������UU���w����6 �軓u����}�����-��u��������.�L7�.:�qCh��Dp��E�"��Z\���c��R�Ι��Pj~Zj�� Nf�)���ݦB;�"eI�癠�H�Q�s3A# I��Np�w\y�U�߲��������oy�{/��Yh��{�m��v�u�AKl_0�{*������yg�8�#G;ᄵ�֎_��WZN���P�<P�.������T��P�/���;~R�������$��58�~������0@̷��0�\$]��U�D�9���c�k���x�)�7�tl��/�@xƴ �`	8]���'�t�5�\����c�=6��w~�_��;��x㍟��'�xg����}M��Gp�������;�5 �1��O6c��J�}�3�Yu`�|%Lr�y7�Y��O���{;u��y��I�����OOp��66-��0P6bKLl������}����G?*����1�]��;�����(%����իx����빠XG���-���=5��z�����Y�Ka<_��	�#�z����gf* E`�+�*�ӒG�;Pv�mۖ+���L�������~ OP�49t���᱙,��8���m;�8��F�MS�k��y+&:�E�L�*�>"\*�.��61��
�V�ƶ#4i���q�� -�f�bDgOX(/6Ԓe�r�dUȹ:V������A��^�|����5@n���={�n���ۛS�}t�V׬:qdd�4:�@�o� Ԓ��L!�y�]d�@��n.=��;�<i:���`�֘UT�&����� �9u` �g/]����.���B�(@�g�6�h�򘳯g��F�����	�ߋ�؏-(/N4槦��IKO?����uuu�X���x��k׮����z�P���T�ׄ�%�8d�Q�Ȅ�@�)jҀ�`!~<;R�V�jcGEq��C��Җl��-K\��ZJɰJUг(��.X������@�F�M�>{-[H�7���t�	�8R׌��ԋ�/�uCN
4�6n?�6��d$�SK�T
�`�400�iӦ3�8�_>�Q��)��9�$��qk�����	'd`-�7n+U��b!�#�P1��3�ɩ���"��([�I��ЗE� ���CCC3v�5�)��C?�]�t\��[GW��N<��&?��U�<Sha��l�2��`eb�-Y�єv,�<�*�䠈4)Ũ��k�|��'���Z&�N�[EW���uTRM�,ѼH2��]�ǹ��yY6����Tj�e8J��͌�����������a*O��g�J�`"FF�OX�r�:q���eC]��ݾF慾UN��8��-��'�0x`��Ri1�+��AQi���U��|衇��Nءj��H>L�~`���M]H�X�H-?�#�l�W�[���=v*v����P���?~޹o�>"/��21��p����a��z�1�:��_}ϡ���3�/_����qک��8�셞�YF������?����� 
YS�ј�����?���������z��c���'x��ʀG���2�x��_븼BĔ���{��f�f�O�{���=��Gjjq��xc�E���(��9���g�f!���o��+Ʊ�m����W��}ltt��Pd�!�bz>JU�G�����Nx��7nZ-Q�/� U�f�����W_}��o(x�	?�����˿��?��O�"����S����_����������+�����c�$x���(�.�7�֫\�Pu8N�`ˣ��x҉k׭	=�C�l����e������~�M���·�����}���s��wE������o���s9��|]S��{*���V�M�;�wH� d�����5�`aBa���
��ŏE�7b`g�`��Y�f�;��W�ڦp���@g�Y�9��XYҬb�Q���_��n.i��{��ȵ����^���?�Ც����cyS	Cwο�5{QW2t�1ʰ�ѐ�#,9��y �7~�H� Equ�,	�Hc�"q��P�\ۇjJ����
���!�C��uM�,�-V�8�NC*6�h.��h�V*�Z	\C�K�i�EdP�P�i���nT��V�ʿ���4���}}5ٔ@Wv�)�I��k��t(�l�

�ˢ���0�g�~�{����Q��X�`�C���./�QY���n*���ޛ�[VVg�{�p�{k.j��*��(� �T�hDP�t'��N'��8��Q���MlcB'55� �
BQUPE�í;�3�y��k��謁@�O���˩s��g��[����we��T����^��+�;S�3r��`|�)F�iH#�XM�p�8����nz��f�홇�bߎ>ph,X���c�cg�}�e/�dѢEK֭\��8�E�L�7�y��r���$�G�z�<"+�BH�|_7*����j�%W����L�:�.X���AH����n�S�XN�Z��j���Y d�z߂�K\g�cόO��S�,Ͼ�ӭ^����P4>]i�3��|p0�x�]k^�jz�N����¾�b�6�A2N�H��i�e� ����>��z�E�Ǯ��߰���*��3�[�!�s|b*�/�y�,V�e،�U�(h��)��U`�����[	[�V��J�����*Ѐu�@�{�A��8=�\���B5͓��d�YB���s
`7/�ڭ���.\��,'�%������l9vh:�)�5�֔��'�pݿ��X�޹�ܸ)83�6|��Zj�J�ws&�0$�U s���x�@��C��c\�h��W�rj|,�������xR�EU2���Z������`��mך�d����Vzz{�T���V�B�j�m8%�&gk���C7���Kw�֫�>�f?�"��`bH���\�"*2�ID�v�Al����ϩ�ҕ���%uFz��T�dx�v�%��va�iIڬ�zK�vڝ��"*G�&��O���Q�`�cSЙ���	u��W����*{�Y=��k�� �B�4p+���*�X=v��?��O:W�hdp'&�P�d&i�T�J)�M*��SF�wb%�� � AE�ovf����o�U{+n��Ƕ{~Zr����lm�ٮ�_4�g�>�
��#��o>�Kif��<x�^wQ� ��!����2��@"|l�p�v[q�2V�U�����tm�1*N3����C����N2��tmE5������~VW"��Qʰ��"��Om��m��1�>6u4�J��R��|��_q�e�i_q�U_��ע$�bDOzf���ӳ�ˮ~�=߿�R)�Z��Z�W_��_��:`�������������~���#�A�j�f�!��t��<������]��U��|�ͦ"����������n���ox��^�9F��&yǎ]kמ~���*6fAz:�QS!G�ިWʶO�kU8}��(t�ħ���D�$�EWh]��g�Y�)l?	��*�%���%�%n����m�:���m�v�j?��c�]vy��x��n�ۿ)�ʾW�;<|��Yg�U�����%��u7"&�"�v�M7]����^�'�*F����O?��O�����P��Ӛ3C��R2k}����O~��x��I�^s�kn��V���Em���?�7���g��^s�u��* �<���Q*�ٳ����K�,��;w|�[���7<%v$��Vd��3�/�����~�AN66H�W�L�4&��؞�LOu���"�L�l�<�-�o�q�Rz���ߋn�#AY�e)JDD�i��If��l�E5�|�."� W� �)�a�x.	��-�}��ĸ�7{����䚝O9^G�����E��)@�#*O���F�Xt���Zm�Q��5#�0"��E�r�:B�'���Kqʴ�װKi�7�#����.�3�{�l�_��,�JmX&ƚd-G>:��)Ҵ��#-��\��&n��q����&H���\,�������j���wY��S�#gAH���%H��� I΁�Gh�ד�;�9�����d�&D�u��Y�$�L}�/w2J��D�� }�N%	�_����8��c�`�3�2�;��cH�2�hQ.B�@7IW�K�j͞F���w�w��_�,�nyvv���s�9��d1����<ܳ�.^��>=�{�)o�*x#Ah�
�drr2LQ�T�.[^�(D�4�ɨ������Y��D`ފ����9��۷���I����� M.[�	9�&:J���)�k6[�Op�R�s�@V��!C�/WQE���-[�l�@�������xf��'�����4<�رc~�XI�;���=,xxR�u0��*�y69��K�%8�ʝ8��E7+��S�n���Kv�~ty����y-�XxS�Cc��͎k�#�*I5�Q����Z&4�l�r7�< LB�zb�e�W*�J|e�JN�^k��,2"���.<�"�(���J�F�hz�p�iK
�>������>3-6%J.+�h�9�"t�M����uj��9`��ޡ=���3���{��[�e�q��l�(e��+ylN��P��Bbyd�[
�,r�pf��	mc�x-����-f�;�j�Oe&�NRK�8a����F�M$<�Z�FE��l;���`E�tM�Ϝ�u���E���z�໷�8WvC���.����tX�R1�
�Y�I�CJ�	׏�k�2��\*Xc��ho�+Ze�r�.]ڜ���bZ8	)�޾^���$��AHBo���6�b��0�@�8�I'����h73za[)�z��uE��80H��%�c�5"�qq7�gog�⹋`��q����c�F ���ٙ)2��/����=)��+/Z��|�k���w�}7��7n� K��|ZY���ԧ�9�������y�/}V�^�շ�]�\��u�]k7,#ی&�>uL�#������>�����߽�kh��,D�G�޸����4���4x��6�ldψ�;�H�:��"��V_R��+E�����JW�J�]Q��%"/�Q8Wb@�Ђ6~N��Z��ۭ��s~�������w���.��#����ī_ݝw޹{���hs�嶅�H�0	'7�p��gv�{ߛ������=��(Ǭ���]?��G}���� ��}��N>����;޷iӦ���߹�+G�Z���oӺ��w�C+H������O��m��F�ɲ�4�/�{u��+_���n���J���M��#��$Rn�
H�њ�0Y��������`UQԘq���;Y�z��X�!���N�V&�\��:���
0WΑ=[|*)���رe7�d�V��K��,n�>Jw(�����G�'� ���
���.X�ɑD�H�������S7�f�SO�q2�,=lB�����%7T"=�]�L�Tt͝0a�u�+U~+��?3ɴ��&5�X�Q��r�TA=�0�
6��u��y�JI`�WՒ��J��/J�~�b�ɷ\v\�ZUig�����ʅ�5�S.��b՛� ��"85�2�5�,İ{{�ڬ�p�E��
�YP���juT�ڎn8՞�01�@��J�:�f4DϪy�ֱ?T�K��ĉ	��+eG�5���I�ɚ�Q*�i��@
�Ve��ت ���jY�U���ȵ*�4�^;ʐ~a<��毆1��=�~8�j�u(֒����b�Ӎ��`�q��5�4�z�Ԁ[���j�FcQ�L����fu��j#��*�[�~-�P�8y�2��f-�F��~':�>����Y&=u9�6�\WϒUK�,Y���C/l7f�&�±�ū׌��!�r�A:6ݬ�m�5ӘV���V*U\r�Z)���Ւ�Z����mp^K8�3i������Fmp`�����Ѣ�F��)�Tn�K2,� ��nn2�mIO!1�u���u�-���24��� ��a���t���LVk����u1��	�X�O�s�`(9B&+ڔ� .��H�N����=X�ߵ�Ȉ=/�rB% ���=���P�v+���	��E�&��}?5��H��Y��U��i��,b҂Wo
ǰ;k$����\���
""-����|�i�|��k�΅���;��}���Ű5K^��lp���V��(���,�{��P��ox͙��d�ةѯ��V
4�xk\!9h�V��J>�ldfꩡ���5[s4�6ܰg"�}�d����&`m�9��TI!a�E
,~�-a�B���r c�	�D�*����z�z�J5�T �HЀjZ�T�H����ZI�!y��2V�2�#9Xa)�	2��)�`�B��q�Y�!Tڗ5�/!0Osu M!�B@�.e�..܌�����N�aj֖��燑o��d�4�%��k�ɑ i1Ƨj�1�nZU׏=�2�jelf6LQ��:t4U%�=��S�a�.��I^���XQLֈO3�k�������WP�*���������n�6Ss7K��ߑ|�O�Alub(�9�����o�v����Ķ�6b]����oO�N��G���W�&����d<��	��m��}����<g�n)a;Pu]�'d�Q;�t��N;�a�nG��X�["9"CK	fI�}���6:6���~z���uۋ�����H@/��?������O�3p���1;s||rrժU�	���<���������Lx�Z����>�s L�(ya�h1�
�q����{�@
HR�h�^L���9z{��l���ګӘ�&���}�+�NML~�Cz�����p3�H��G�V����9rd͚5�V�V���pɐ-5�ٲU�H���kV-��w�v��E�t����K$���������������
�Ա-)�Hcf�%KG>�鏽���������n�*�|�mgoܼa��XS,FC,^p������10��������es�~�k����SR#��T%hG��qʔq�d|��]�I���l�μRC�|�VF��#B,^���8����ؕ�ђ���s�+�V��*B�=��]�u���2��ԟ�*��-Y�q���d�.f&L�>p��.��/Lijh����K�Z�:"?L1e�-`�߮8�cø�5#hq��b	_!>͇��<x�s��4M5u���?_�s�}-ٹ�GR�O��%��z���9묳�����`dْ������"2�zfgg�|r�hҹ,%�}#����8M�Y떑�\�b!mH������\�5�?�l�2���� ���6n�H��<0>6�(Z<x�\��ygd)��p�H��Oƽ����y�{���1g%�����<ɲFFF� <�IE�u�N��KQ�I2�${�5H���TX���������Q#�߰a�J�l ���G�����v�Ⴁ��+W���m۶`�b:��m_�;p���w|��?����a�h�==X ,ޒ��Eµ!��8�%U�3y�����+����s�a㡇:��Itt���窫�ںu���$���o��G��k�t΢�A��y^�V�y���G器;π�ʲ�A�M�-p�"�ғ��ӵ��i�5�a��+W���/�|�gf͛n�il|J־\S
u��f�|�������K�3�c;�z��@��h qj+:G�p)��R�	���"���ɺX E�XD
�u3���nV�y61P:�ozM&Ͳ�'ZU�J�G�5q�p���3�.W��"U�e,>;��Xx��힕�^~B4*�o�Em��t �H�\V�0i�?7U`-�k�9w�٨`��@W��/�/�`(��`Z��J���q6V�X�������lzɃ�a�o�`�4���� �,w�2�&�!�.�QP)��_�`8�������OՔy�R��Vy�E�X������a���2��b1��c@�m�?��η8��9�̎ƹ�	�t	��kc+���@x��]���I��zw��w���Wi�<ӨC_���@+����f�j�(E�[���r|SO�!�@h���رc�\r�j�i~���Q�d̖���99u���`�Y��ĕ���ퟚ���D�I\-�ŲX֮][u��=�ob�������9�Ո��˗�hJ��	�"S]2O)�ϳy)]���!���٭m�20nI�k�.��K/�T�<Dr�L@�R�a���~���	���b�HrRA�Sn�������>KW�cD�=l�w��A�󒗼�ܱD3����n5��B˖-$�=��i��������<ޢ�Z�f������~׭ı�����<������A�L�P��H<���� {A��꾔웂2��2��¥9������9�/�M��BV�� KzR:�+� ��2L�Y�bRn����~���*��vۣ�u�O|+Ce�Ν;ɹ�>a�N2���X���>�{��#�a�؂�P�Μ*�	.��"ڐ�qzs�������� �u혵әg����}�v�u��%�J�N az~���~�QvP�r'S�֮i��L�W3;�S��@E�/����w�3���M�Iu6?�vRP�v:'(,.R�)e�� ���Eɫ�b��&��ŭ�rla���ba�ț�E����'�)�Y6+���z
~�̠Q�s���Y�h����z�A-<�bif&QFE wh��U�Y�Eo������݃7��;"q:�<t��.���Y�q�JH��I�PC\�a����+���P�p-N�%�a�F{�՘����7@��1e�"/��Z%���l���"'�X"ￄ�Jd�7�Z�F��*id��j�v�w�t��ĸ�p�Y�T\��g��^�3�>v��P��l7��d��K���#��M4�$s�~��7S���v�\�(��]�Ơ~!CO,Gv�,c��"m%�5#�m�4!�tv��WM��5Ҽ6��4��!$(���O�7����[>m�q+HiC�A���Q2��z�q`}  ��IDAT���(�Wk��"�CP��2H�b�+;��I�V�Cs���m�Sq�D	�*�6͚��t�z�$؆j�*��r�����ѣ�S�O��ў�58�V��6AŴC?z���g���?��Q�>�\2+Ffբ�T��藕8���H����a�h��H�ǋ�]h2�DP&C���'}�r{{{k!�<�i��� � �)����"�����kQI3�˰�j���NS:�w�#	�B��KFOةS�Nl q1�TS��b�hy+dY)�/ăm�9�%N���"Cs-��l�O��4�;��u��N+
#pj�e16��lA#9�سD<@z����=o$Uܘ�'�d�w������^��K�I2b
8��!��	r!7� ���MCM[-�$^�t��E�,X +,�ɥ<66F�Mmbq�������j���c_����~+��L�ֳ��#�p�Tdჲ�y�4��ֲ69��B�T��N���(~@Z�e}e�x[�3�0ǆ�ڤ��z��O�s~,do'������Ͱ필�!J�K����@~z�jv8u�-��I$Iʬ��_���K�(�oIV��*�1�[��������Fh���X��)ቁށ4�ɧ!��aD��V���L��Ljq$�@�Ԏb�Z��
銁���� =J�$�I[)jqݾ��?�|0��L�@�l+
�s]/U*���o��_0ȕc3��pXn���[� ����ǎ�:�.Y�E��n(��{A�;f���7P��9�Ƃ$F�=q��`����Cr2}���0�cH;�-'�m�?����ĺzw:S�K�����M�"U�޹co�T�.^/_��Hr(��3i�ep8}���$��G����L�ȇ?z��߾ꪫ��H?k1y8��~�.;q��O?�����˖qE5�n��`�6�B���r�j�ZoO/��$���w�>��={/^|��1�>���c����ϲ��y5>5�����*�����5r����Ts���o$�_T�Ay9$�/(MtC}#�c&h��%Ѝ-͖,Y�A ;jP-��#o���,	��Ė�X�J�5U�������W��U���r��Q˲I��f�13;�����tÌ�
��A_�9�����yV��;���J,�C�vO��F}X���E:���2�\i���f�����x����{�����jީ��4O>�Ϟ��}	��x� �Ԯ���E�u5�*B�i�;����E����,awI���8��3��iD��d��	�o�`<@M��Bјj�OW����Y��	�n綈��y�Aq_3�����Z&�S���y�Ug�A{�L�?��c����_��͛����c��������l�D����Thr�去GGGg��2��	R�}Z}���l�'�x�^��}�
�`o��v��#�Mr�����)�ĤFK3ͧ�~��G�8~���l��;ځ���-�js�!R��^�C�ң9�?3�y�1H�F�g ЖS���I�/ y�r��	�r �D$ؙ�	
2�A�
���A��h�ؾ}{�ZJN�Z:�aOXY��[��>��d��q�Ƒ��sN�Z���k��qh���4�k��J�9�Uf��h�}�ȥ!f��V*��%x�Z�������ڵkty�����E'����x�ݻw��g?���f���Õ�b&F�~�-�ڧf&�Wh˧w����ߨ�����q�[`lU���D�Z��q���>����Ǟ�������ַ,n=<19=55e9��t�*X7�}6�8�����E_ �F�6W�t�̺�4�d:e��f�C%�@�3�0,�;ʘuO��m�W�{'/�\qurk*��a�4��9�:�[�� B����?���׶d!�RgW쿓m�n�J��➋g�)c�����R@�,.%]�d.��NV�"�\QfHx��dfj�ܪZ�4�4k߻�[(����vШӘo<c�uL��s-�HG����iq<͖_��#�D����A�91$'�����6��,E`9 ���NH�b�r,5��L��oE>��`�S4�Ҽ�$<��4�?�W�)	��`��i����V�oW�n�c|d7@��UȒ�#m��د�g�IG��ڡj޼yr�fˣU`W+�t��t���>�$L�@��?��!ԅ �Q:�a��[�h#=f���u.�ڭ�W�G�9sy�_|1i�G�~b�i���FS�J�c۶m���w�}4�R�]�x����Mkv�5�y��bs��A���� ͂eKY��|��M�W�X�b��駞zj��S�M]�t�3��jC����|;o�Z�~K�Wi%S@�^��|�IR����c�|뭿����)�����W��U_��-���������7��;I�\-��]HW�-�C��83z��LiB�e�~idh�i�r]-J#���Q��S��~��<� �CJv��7�W���w��3��������n��&���m��	t|'ԗ�t�+yQJ}Ga�	I�AyVu�,C��P�1W��Z�P��{<3I�Q�s]���$�\�li��$6�N߿[n�����7��%ژ�k����[o����׿Ey�oa%6}��]�M�}���'�N7B7�p�7�q��G}tÆ���8���f�]-�Z���{�=����+�!m�Jt��>)IZ�s��#��j�{!��~�!,�]�v�N9�V-�N󷻻Lt*�$��M;�Sc��H��^}W~��+�DR���N���:4�(&3�RŴ�f����HL�nkj�+��8	Z��Y���_�$j�����)e[l�	sNƍh8��a"�n����Ԍ�����y��h�M��ʐ�	�����4#բ �-R���F:FCw� 	b[U�l:$���w��C���+�Y�Κ��Y�C{��d�TR�z6��F��n��%�
�f����
�OM8'j�əZ}tl��0U����R��j��#�g�w�4�;��$'l
�C�BS�ݣ��@d���0�>mN7P��@��'���x�jQӾn ����l��P:b�]��6r��˲N�[YA�jV�An�xZ.�6����n�ܲIagI���5�<�`��ri��6Ӷ�ԁ#3���˧l�<2`����em0a�LM�*q�]"�V��/Md�eQ#��8,����n�^o������	��ׁ��Zs�Q��z{�Wa���JV���}�'����F����4
ș��x¯ѤZ2�S�_�/��*A�vW�p̞6D2��T���FsW/�W��%4�������)��d���rQ�ޱqY2ฤ��M��щ��^[L��i�H꼶ϨO �J%�2� ��<`P�X	���t���ʏ.���j��O�`k>�l�ғd��\`�u���ȡׂ��z�}b7˷H��F�Ӝ�[ЭiG����"�#�N��)�'�W͠���J��@%t{��6!I���"��WF	r�&��Ve���{�!����-;m߳��'��M�Zbr�>���lӮ�&�*3/j��p���~D�֮����'�Ac����p�Q��HE	
��YA��$�q�E�'��}�:U�(ICNg�e"3�'��l7Päa�D�L�}J��y(]z�6��=s���TG`fmM��7��i[&��ѲV�b��s�"��9��}N�� ;Q��0l���Rq�óӴ�b�p����47��L�k`fW��M�k��*�8�1J
C3\[�i����k��h+Ԏ}�~*&1D��J��3�[M�]��=::24l��TkW����Q<%q���T�"��7P��x|zlrv4�ڱ��R�a����ˠg��'Z�Y7ܪ�3\]���ڬ�8=��Ԁ�v�~rN[��)�{���~H��I�� Z'Af�g���W�����=y:J��(����sC�Y~�.
NQr��&��2m�ٛ��g$9|ҜC�������x�k�J6p��B�Nɰ1�(&��ls�pȚ��=�G���?�{�S���E��N�̍� �������	ڸ[$=�0�H�릥�\�|�������s;o�6��$�lܼ�׼���oW�^��I��(	��-���6��P�RTmIn�Hz�b0p�$�(_��z��
��\�ˊ��ڏ#Z.�g"ݪ#��f�A�u������Ә�gx+���-��B8@�;A3�D�I�gie��!�o�k׮��Ǐh��y���jq;L<�޼�_�n����-�Ϣ��0~��P"��Oj��G��f��j���o�}���hl"����}��lv�~*�V5;���P�_�Z�G���J��S��uT6=U%�,�p�2��)���&}��7�,݂49U���+�i'�"��"�HkMx,���K���vƁ���s �k��c������:��8)
�]-]wX䵲J$��/u\�?����q.+�(/�4fŕ�TuJG�]�|y��w�y��ݏ<������;�<R�`�+���hbbbǞG��G&��h���`�_��+dm�v�m,X�dޛ���+V���2p�6����{�{���{z�C�ͶPq788(�.��Q1�s�������ʢ̯HK��"	*>k��1�p�GD�'�D�!�\�\z76�d	QL8==�27���DCa+"��k�uF%e4mx����o~�i��߿�3�a7�?sxx�������zv�9p�=�[.XQ��]X��<,�o�B��tp�5kV��]���#GZ� 
�ٿwϞ={��>L�֍y��)~9������ j�nG�H�����4�S���'C�B�L'��&��;]M��h0�d�7ovj��"�T�t���u�Y�-�w����۷�L�o��ȱQ�*Is��0DE�ic���z�MS(v�t'��,ą9\�����!�������Qs�|�<�2��@��n�I��Lծ%&�\�S�GuA�
�N��h|��t�G4ŨgHr��h|c�t����۔9Iuwg�Ԯ�KSr*��J=�&�`�G��	j���M�pfR�A����n����-[.�p+�ʡ���5��6#�'��߷�.U-�x�}Z>�KkL�j-� I���_*sr�N��"+h��VąOR��w��׊d�g�PR^�n�|X]Y��1{t�U��B�;Fͤ���d���U�&�y��H6}� ��Os�q>�,!:G녓��IM��srD��(�$%�2:� =O~�����C��2d]Z��4��	C�UK��O�豳T�얒��b_6lN�g�	���*����VNٻwoG�]_vٶ�n�|�`��y��\��r��2j�r�-��v;��*9Ө��%��rWYZe�����w�/ڼy�%���x-4��
�[�<DZ�99I����{z�0A�`Ϛ�� ]��}VE|��	�v/���	%fѹڲe�~�>N��~x��m�Q��o����ѰVU���6mڄR�X�a�Q��o����_����T7�c�Q��\c��_�F;�;�;��0Bw)�w��o6i�>|��\�t)-��9�C����)4_���eqf]�+��v��d�h]�8��p�����s�����t5o�X�՜5N�MbkŽn��av�h��/�߿��<�Y�O� �a�������=8v��v�T��z��/}�ڷ�Z��|�`�ɼ(s5��6�A�9��-��}�G�����U61y����<����۷Ӟ"ܭ���g����ӹ"H�q�s%^��|�_�ȃ5�=�&���W��sn��W���2c'��ڱ_E#H��d����6��MZ{����l9��GwL���UTH�q�4M � �&�S�K�Q=�����M���8*���aL"-�5X���[��ֿeD�V�3פ�VS ��.j����N��d��2�U ԉI����	ۮ�7.ّ���
b��n&����l�� P��L�( ���Y;i�ni{axdlh���0��f�i�o�a�?�c'��C�^���*[u���Y���ڥ&�
����	/P��@��C�}3�mi����M�cO>E*���I�ARq�4<���B/�@Y�T�  g�Nɥg��$'&+�n��"���#e%�#`LWh>��u�|�6tI����A�L[�/,E��e%q��๹��c��i)0>q�j��eX�F�!*$����j�Z�lOz�R�����.0�Ώ���z�Uv=Ӵ��h��n�mg��4reܹ���PRsf����`�k[Q�֚7��,�7S����+�}�)�'	k�&2�t�\�8
��,�Yo�u�J��z����>��ٙ��l��zV��O��g��&:��M�'�I��Ik?�R#D}|f�Z-o�B���?��,M��z�M���N�3f� ��DS�3o!���D^;���0Aރ"LUuL+҂��u���<ŕ1�{��8W�s_ag(d��<w��oQ�3��Π]�(Mh�22ۤuH�c�DA�"��qM�@�IV��j�^c���XJ�@GC��Zs��Z%DUT�~���4f���E�[��`0}_��H�fP�#H�Dr�� �z~fq�l��|��F7*��v�N�=�{��q�f�Z蠭F���4-~o�7R+��)v�<�NmP�J�`�:hU��)C��ff�
�׬��af�R����ײ��z%�5��Az�"=�M��I�T�M��v+ ��q�b e1�^���,����0 �/FS��/m*�}@�j.�X:�lJn�T^���~+e�W�I�.[
���:-�N
��a�M~}$-����u�o���Ǐ+&��e�Z�j|�8TV��V�ݠ{��
�@���L�����	��`I����TR?۱�8F;K��m3V�o�FJ�u�͂�F��QǪpz6�Txź���Rۋ��?r��؂��uk`�&I`h�ѐ�=�޽��k6k���&	i�*MF�lR�i�5$�m���Cän�K�A�����Ҝ����ZӀ�Z�=���{ 𣑡!��8�;��>W/1��]Y��4L��Av�;0!R�<N��9��tjiY�$bY��n>�̿�˿���7_x: ��ƹ�*h������͊k�y�ǭ�{!)������r#)���Ǭ�)I2)��Xj(#�PM��׿��߾������Ϧ�+QG�PZȕj��w＿V�������0�H"#�4;yk���Q��{�ާ��鉱�n}">s��X�tq����P�� $�q+�����W/v��蓼QjQ*�>��-��(XaHr�զv�����K_��o��'\�Q�F�R���ٙ�#Yr3�j�I��
��h����(w�D�$�iC!퐚��pKK2�jE�fV�z�˾��o��_��� AZ�2P͕l�.փ>y�X��~�=��>4T��9~|�Wk����S�=}x�.E7V�^SJ:�CWA>Ю�������ov<�z�C�N�C��=�SyA�Ȟu�Q�	�
���jN{�x�7�bUيe���]��N��њ+.�4ב.J�bQD���(��ZQ�u�G{�g�~��Q&�@$^��~̸�5;-Y83���yi �&̓x�m�e'�M�'44�ٹs����O�$ٱc�Z��\���"3�������V$���g&9Ν�&'�o���޾�����ڷo���Z��N��7m�K�{�������y^�V���vծq�1.�TJ��T���mCF�2ٓg\(h!o�1֢���l�67�E
B����:�� �[2���l2y.��bG�M��8���zAMh���m4��j��ŋ��̛?~��@ښ5k�m�v���?����f���3UǏ�U*�ʼa��vOO�����s�A�*�7lX�v�w�����u�c�=5�������ի�C��O?ݘjӴ�,AB��T�o�ͣy=
.��a�*�7թ�d�@eȆ�	�)��a������#�3d�����u�]�`�P�di;#��E"�����X
U.�(e�b���i��(!YǥҨ���"��tp��Xs�ЩQ��<)����terW���܃4Ũ9dL?�W}��}���0������.۱�Ѭ;����Ns��**L��%%�0��&�����g
D3���Y_��3��LN�lo��G��'%����Ï?�8��p�^OP�4/�L1�F���Mcs�/Y�_�e��̠i2�VV��I��<㡶-3�;5��sJ�P&�%SG_"�DN�'��G���J�T@���\xt�sl-'�35�(XZ����k���f�Eo+xwbդ��疜=����X��.���ӦMkW���#�����W���_L�$�G~J�m0�����%����.�/ ���y��"��Yo� B���1�ZԔN�A�aҩ�|�uW� 9�q�1!p�]�i��v��s���Ͽ�<b�;�5����>z˭��#�4!o�4o�-��"E�5�<T������Azj?�������Ȃ�L���{�>���;�> f^ip�rQu6�x
�y�������ݱ����<��ߤy�@lR���׼�C��G?�ѕ��|��^'�k8d<ش�X�H��.(�c)����]���(����P�qb�UW]�b�2���/�|���h]������8����?HWx�;�!+w����<��1�HN=I��r���� �<N������׼oj�O�8N�7m;	C�}�RF�uO$M֑@�̓0�V5Ln.�r(ݴȵ��-�%��k���>���.[��mo{����i�:t04J9e=Q:d?�+L֯��A����釾�<::/	�&���o�o����\o|�9�G1R4������?��?�]��o~�������7������ݻ��{��e��3��Fh�����v��n����~��Y;�p9U�8��[%=Y&���NV�µ�b����vz2�B�=ۈ��HL�,�{I����ܞʧz�$l��-Y�qzHZ�(1RSA��3s�C�j�5�о��c���&��3%�|T^ƠZ6��Ɖ/ �N�RӘW��g?��ђ�U'���@H��B��u��\|��+����7D�=�|��'_�7 ��9|�lw�#]�����kkm��n���Ȋi��M���'�gm���N��<%@��Q�n���;�>��,�xU9�o$�֡XM&f'3n�R�U-�5T{[�894�G�j��N��'�%�>1ٶ��2�ՊMƹkV��~j��8n+,��R:2�H��ؤRi�g,�[4� �O� Y>:K!�f�.m�ϱU
H2J��$W�$J��|2@�f�dR�$�A�xG�|�s��NR�W��Go%JE=�fێE"]o��ta�p-Iڍ�t<136����d-Y�a˖-z��;1���3WL�&JB{x�bۼe��I���=���x�G������/K�m9��b���)��o[�r��V}vz׮]ǟ|��,�`k��ͳяhĂov�����_|�[.��ҟ�����O�֮������W�Z5�}YW����#q��἖�dGn�p:����`�(�Ѹ}�Ǐ��~�����]�� S��$�*�*P�t�0a�?��X'��Ghӓ�C��%�i`R�*��(��������]���Z�dx�њS��C�����"A�M�LՌ����G�]D��`B/W���j21�=6�5[�����T� E���f2Ǐ�s�6��'����,�4��$o���!A��K�!ABIz��eZ���ғ 8��'�4�SS���O=��;���K���}z�f|�� ���e� S�G�7=:-���{zl���;9�9���W�v��+����&�m>N��������q�G֞F���?�e�֭�S����n�*9u���c�J�1J����[-���ͯ|�Ր�4���?>9St.�I���I����_�dR�֡�G�gD>Xܣ(I�H���9�=Y>lJ�	�1�	�tΡ�M_EV��{͛߼t�z2�����ħ���n[�t����:�����޽>�����W\���e��k�;w�9k�ҥK�-^Bӷ�/���{��ֿ4¦9\z饛�o�q�����Il���;�nj��� �O�vt�x��V����HZk�� N�k�a{�\�����^HcP�ۉi��#�����~|���Ӎ��.'%pէ�����I�_E��PYӬ��ʽ��fL5��D!�[����?������_�q8c�`F'�����L{ƿ�6y�6"GW]�
���n��N#�8j�Ac�L��b�=矽�K�S5��E�s�T��K��h �r�uR�<݉��Ͻ���|˛������﹟ȵ2%���>{��c��u5�nn�J�o�+�J��s4�$�"�%��Gj����鉯��w��_���_�⋷���|�ߠ;LP�h�����W}S��7��M����t�_{��>��/|��_�����Qڠ�y�>���	��`�04SyV�H�2]:a��Wj��V�YN`#�����R�ۊH"K\��w��EF��(�ә
Tj�8��T���y|嫷^z�e��~�K���;��y�ݘ��=���km �XP�����-��M�u4�kF��=�V4��Ƒ�Z�D��Y�c��t�d��-7m���/��k~��_�r�գ(t5��������=������ޅ�?CO��k^�g����K^B�<��K���_:Z�y���z��d��U ��٩j�?
��������8�sA��I=���;R�'��e�Qy~u�\���*-EZ]t������a�V)�hZ� /�t2\ \����|++p��P5���[Y	3�댪ϔ9=�t"7'1g/X��|���N/),�����˗_t�e4�w�����##���Fm��8�r�v��==3#������G''��~�_L�����Az1͹�F�PQ���Y�2��|����L�tH�A7:%O��L�$����	.+EEo�%p%��hsDs��G��D5�ògRDTJM���T�̗�I>��ض9��k�o)M��:,�*۬���Za�j̯h��j"^`if��;��"D�]�K�qW�6��<�3m#�;�}� rd	ͅ34D��tm����ܷo��G-ZԳp�D�g���U�E13Ӝ"ɲmL��L�$��km�~��������U]�lٚ�^�����^�a&����IT֭[G�����G���W_��O���n{{�G����yyS���_���v�6��(��7v����w�R���.����}��m��2��iKJA��(��N"ɶ-��e�)��A�!��O�+s��Lf��խ��.E*�yb1�Vxe'��'�O�G"{.���5�̛��$w����D�s��;m��R�NJŧJN�����|X:=m
?�8�xGF�Ht��;7���J�h�S����̀8�4I�^�����,^�x���8�f4���/�Y�M�鑞����Wξd+�m&����x�ʕ�Ȣx`��S��X��wthȮ�ӕ���w��Fv?�F�#��4C��A�Pe`�EԂ�d��O��4%a�����=��&��/K���I�VZT㜼�.����|:D$�N������͛7+�***��?�NOO:t���Q����~򓟐;
F0��h173����֮]�ģ���C��t�g����#�+.]��Kd����bL�L�p�9U�zI�^f�܆.�K�r��J��U�9��4�&E�:����?��C���#�&������J.���K��֬ͩ�=�����#��9ìA�<RV!s�Y����j���7.X��6z�j|��	efyʷ{��oDB�� ׈���E]t�}w���r�,R�8)��HnU�$��?���nD@O�K�N��t@6�D������K�̧���K��/���;��
-C�aD����}쵯}-���=�f��o��?��w��o~�����4���n�="�v-'�f�+�z��J�[ -�?��5Ւ��ֺ�u�g��^Sp�r�
ͦ1���1��n
�#�r�Y��e˖�����-��.C�r��Cմ���V��O|�=�zR���s�X�$��Y�8h\��kg�2ltz���as�W9�����і-}�ߠ]�k5ݒ�zh����|�#�~�����N�ѦM�^�����i�U2H>y�/{��_���>u��D:�Z����|-�x��H=����O�P��`F!�m`�9f�,��37��%�"i�D�-���E������U��c2[W���
3K@�0�όQ@�k�k�el �m�����I�8�,�՞��΀<
��+�(�,�"�\�(��P8>-o�e����Z�� �*��9z�~��k!��42���$�n�����׫^����W�P?���Ss���gmy�\p�7oB*�-]?p����^5z|4UɍT6����;����.bX�=�6� 5����qΒ"C�s9��::A7�����S�19CS#KbҠ�&/�bqk��d�ʯj=l���i�9t���=s��7��ݽG�>3z�Y���}ɲŪ�X��b�i���9�p�9[.~�ᇽ]�5�sHP4e�JB�f�yv��Dm} ��5�E�ga�K��<e��l�h��cp�y̜��o�a�ƊV��[�Y���]k�ȉ���fd٧z,�5ЋW��5>\�f K�r�R��PK׬��:l��.�J�YD��2�З������O{-���(6?�s��6h-�*�'z�����n��4��nKH.��:�`���2�U�d7J��2��VtVhON��t���Zvlv��p�n� \^k6�]b{hY��Wq�C��g�i+[8-;�t��cc�z�>6�+�s�qx��u�S������i����<բ�.)�`����y���h��G&�]�8�Tj%�ݜ�,{��m[/��od��f��g�f���M�O����c�d��ԁ=sw�u����]֛�pdަ-ȰU���է7g[���'�զR5�N���>��okY��Hzɵ�L�
uq��c' ?�e��4b���PAX�4�"����f�T&���u���I��l,6�d�L�v�����]L��nm�$5�v3�p�֕���JO���.�P15Ӧo��t��[���z��Pδ.2U`��]����c~��5z���7a7(��c%���0���4F&�:��2��X�o"�=HF�ghF��8e([�5A5���~$�Lcf�k��םA���gO�b|�H�og䒮 ��f�wǎC�뙩�ʒ�4^v����mݾ}�7���W\1ddlffMOϹ矯L�/9m������L���ߴ��E��[o���W�j}	c�ОGC������[Z�>��=o8��bC�d&�-�H5K������d�e)٬ �i5-2sѼޏ� Ͱє��j_�wp�~q���Y����P%a��o)�&r�Q��/�&ζ[!����.Z�k�Ο>�뮻�
]cŊ��3\�Ѩ<���T���Zi�G����8�}Zk���o�[��z��Ͽ���LkŪ�dL/:sU݈�ѹ���0��vf�v�8H\3TB��R��u�� i���ֲzJ �*-���L����j��Pb�{�V�	Ʌc[m߯7Zim��B��mƦ*ak��$4I�p\ފN����(z�1�7��N�k�,M!_���q,A��V��/X�m۶'�����G؞}{Z~kvf*K�PM@&��=��mB�Wb���p@�> �� ն�jߙk-��Wl\��Ӹ���*��G�F�U>c�.$�塇�`���a$=?��G?���a�aO�#�R̲��J�g�%W����HIp�J��m�1�ĵ�r\e�v���Һ����/_��}?毦/�˿�կe\IŪOs{ْ
M�k_��o|����y���� 斍�ru��B�(�3/%X
�ŕ�'%�:)ߜߢ�o�����L@%WP�E��I~E�$��L[�ڴ��
��%Ժ�i��=��
c��[�(֭\�Z�Tg6X�?�����i�qօI��N�
�Y���w<N��T�$k��eJJ
�m&%�@����m	�������̟!(��<�W^u�7��M��Q2?i�����;�{�>���&(YL��C~�{�s-��}MuՆd@�8�;��/`w�߁���5���8����)U�[qw��94�m�Tr荛���~��ۏ�|��*S� E��W�ڭ��c�N�i��@�͖S*������G����'6n<a�N�
������o��w���!&���y�k�|��BДy�b?1L�M�9�n� �,�DO�"E���y�Q� L/B�ݫ��a'yws5;�+wv�I�"ϲ;���?����o��D4�<N�F��_q�5w���(��q��飏>y�i�}��׬Y�[V�%;�j��
|�!��_�{���*I�޽{7o���׾q�0�I3���~��^7m��h�҈�,;"�7Z�p!��Y��L�˧
�e�?՜0�?���-�`M5��g�بE�L|oM�h�e�@�Z"IT.�1/^,MfZ�6ٸ�9�-]�	O��&�j���jk�s@l%-�	�"��M�Nl2&�^����R�!�"S���Q$i4�[����Å�˕�2n/̈́�	I]=�J�A�EH?�{!ؖK`�
������+�/���/��|�F�HN�V��ڵ���:W
eܰNvB�e�E|<]�4!M���\p]�Z���!Yj�?��w>�o�>#l!��E�����ɤ�3�:g�y�;��N��u��i������ӧ$�hF��fp����|�"�9:=F7|XA�Tu�8�Ç?��c��̛7��M!�Z�D��?FW��/���b1�M3��%�ѳ�D���Kb�k-K�S���FȞ��v�X��E酤�ؙWseI��Pp�"��bW�3�K��Z:��ly��Ua�ț�b̺��ٳя]^M�}A���e��EGi�F:Y2�^�hK�9�4�?�0��:�0H�h�'�e����D�\����RFV����������0ϟ_��Є72]F�D�5Ӛ��=&uD��(��N��q��D��iT�1SA��{X�R�17�dD���07a�e�� �b<�1��P歅�m�HZ��U���芜��YD���$Տ�|�o��K.��E�aÆ�jO�R9�h�]�� O���M�)�gm�رc`�ɲ���%K�*��N��uX΄�_�_p�G�T$ɪ�C����6���J� {�[��F5����jK)��:�����s����5�dc �G�[� @����^4D��N8��֝���sϝ{�'h��OIQ�v��#��_�K���Sf�������j���Q�BOXr�Ӱ$7ơc;��^�0n���L��f	�SO=eZN�|��n������Ȏ'���=�qi��%O����w�F�[n���8���u�Hj>v<0\T��z;��zwg�~�Q����Oa{/��DƟgW����遢�b�@���4;ʟ6U�j4�gIyW������_���^{�[��V~�8"�$Q��Dۥ�`��YF�&��>��'?y�7f�X�Y����)���>��O�ə�����2
0�t?,�P^�n�)�����9C$Ul���Y��>D����f��B�5m6[����#���?zW���Iˌ�z]����w%��I��7�~��8w>�����4C��ʮ�y �{��G&�S��O>�'���P1�q-�Z�J����_��O��Yj|�?}�����M��0�"��g)�|�Ĳ����'��9�r��z�!<�ղ���i�/��P���Y�*&0D*�8���}�g�����u�<R5�[4ȩza��2�O����������f����G	o?���~򓟻�ʗ�NT+v�(�a�u+���t	e���`�C��}��;=9^� {���x��ݶ���59~�l 1����;x�U��&ق�W�]���������w�U+Y�x#8"��\-CsT.L
Z�OX��ra=@��{^�qu���l��Ԯ��}�p1+Y���KY͑Ԑn��Bmoǎ^۷L���r�kW4�1`��,�pԧg�+�ІƷ����3W��ux,X��b9���t#3H�Ю^�4�r�$���Vm@��1��ͼҝB� �[mZh4h�M&�4����V�V����&�.������ۦF��oh���V�ϚF`h���5�+_��u�֝�a=��t��~/E���?w�oGu���3��ۯ���@�ѱ�q	`;�yql���~�K\�8Nl�[���ر���1�!B5MF�^���S�L�y���=�$����7?���h�̞=k������S�nڴI����OW�V[�Ӄ�J8<�U�-c����w�9�ԇ�E�[�,Ή�	x��d��䮝0��L�i���b����υ��ϟ�0�mj�w�~��u��Z2o���X���q�K{��w��6�̲e�\V��ou��ȋ%�;#��[o�86�h�`��/���y[G� �+�g�{�1\Ө�*��1z�\;h�%:���3�r�K��Q�2��M^bD�*늁EN��;dx�Y�K��a�4��O"��J�`����(���7���9���q�P��Ȕ!�}7�M�N��b�Li]%�ֲ}�zHM#%i�� �aJ�@�zL�� �!��h�趍�k��P�I!>��G7���;��m�YI����"�9�[i��&�+Ziu���f*ܱ�T��{��>f�B�{��58��U����b������ V�Ǫ��[6+2�ρ}����˗/���{pfjos����������;��l����g� �a���%aW�`f#����N�8J��xc��8�z��eA�ڞ]ķ4l3
T��&��<��:a2�"(���\:a�Bx�~bX�ݡ�"�Z:
lj��H|"�򅂃Q�U(���][���К�A��횉l�R��X��+���#�����vx�,�ה
b''	�f�W�D�zk0�#��jy`�P����p�� ��z��<xp��t�m��E��8~��������ɉ0��h��`�!�]��/u\�C
J8 ��(y�k;m n�slC7;�|���,`�LL[+G�������%���e�'�v�������x`Px��OL�,�m�_�������?�9�ܦ�� � B5�-��!��I�����?�W�J3GR��Ĥ�<^x�X��b� ,
�+9Q�<}D�G �B�2k�d*�,J�K���&�(��c��xxA�l0��j9�W0Ȑ||0E��5��65��}D���D��9��ϐd�&�fv'[��t��-�)+��v	�:�JW-���sJrN�0Sz@��b#�gK�EqX,9#�m?j��/]�؟�fR����Ճ9֒��aC�^M�#�y�b2��ja����u=Ţ"�Lq�h��
��¢�P�9���0]Hצmp��Z�A���l�����t�M����SNY�zM�0���y�]�/|ᢋ.:kͩ"��}�{�_~����9�Yy�o_v�=�\����w_Q�uU�s ��[n��r�ڵ�=�`����`!�!yD�oܸ��w���}}}�_W�\y���z�k�z;n�alZZ$���H�ŮPv�p��|)���_�YK�#]��x^EIF��;w��c�}�]�&�S���g�i��t�I0-O?��ikN�f��kШ�x򱇿���[z�q6l��1e��Q��/�����k_���>�	�P*��ѱlx�Ys�Ug$2s?�Ԍbǎ{�o���.��`|P�� y/���l�\�ݻW���	�`�|XM�����:u�)
���R4Ϩ��\��nĞ���Hف�VHæj�����l����mW���vy��R�@eH�a/�3.�O�w���$s��e<�,��9S���s�:�NW1<��D)�f1_�oH?U����f�զ�*�~��Z�ѽ��+�;�3p�H���8s�\������ַ�9�,@A�4����n��w�����������d)����W�T��L��}�U�-\��~��_|qex��h���
�f���M�?_`�x3Þ�6RS�.U�*0�={l�=���	'�y�.�����]T1� P�彟�4`u�n	�\���a��ۻ��:������K˗nݺ�P�4]��O��۹s�h���X��FZ8j,�R����I�CO%�h�	
�*$�-P�D�an�|�'�m��s�y֚k��U�����΢�V��=1��R��H뾈-ã��ǚ��Q�\Jsa洮�����r
x0t��;��pG�L�fk0}v�r����v@6uZ� ԅ���|_[�����e����}u��n��jmN�>np��잡����c�=��#���]v����կ�v� +�#o۶�8�@��Ż�d��V�w�y�fZ#��ӊbbx�V�� ��<f���������/|l�"N�3��LQ��Q��c�������Cd�m`��D�, �(���i�2*V����8����3�<#J�U�`�a߼N4���{_xᅰ�<�n�?��E�͎��i������O�C�n2!L�n �L5�<mc������@=��cp;.tLR�E��,r��Ya��2�%�i��VU6[�#��>�RFĒ��F�}-�k�W�DY�y#(P-�fm�Ѿ��K�cAW�dh�;��G�_����I���1�PN�C�\�{���JWVr�����Ǻ�����Ğ��m��^�3��cR�VHk	�c���A�� 
V�#*�,avM�I೩�(�r����{"3x��E���b2�8/^=���0$&eAr�5�Q�������MK��	�ӥ�Rd�?40��}���V�`	`_���^��}����� Y�a�?#����+�\H�Ȥ�(��p���f[�s/�;�rN�VŘlMI�������At���npv��`�8��h�;�=8���';��O������֠�1������/��]w�s�)�٣ ���� ���.v�-�]q�w��~򳫯�lȫ%m�-�����eǽ�w��?�u�}w_w�;a����#�s�w(f���WbI1�`�w�}��~q����Ոmt��z�&S��+�,�i<\�.h@�5,����#]g.,�R��^��{M��\2�H���F(�mǶtç��G>�O~�������TaJP(��I�Y���w���������4SD��.�v�C���}���V�J��(`�Ňt�?b[����)�?��C��^RеE��/��ٱg����MIm?t;~�}�Iǯ>�����>��c�לqv�mݺ�(G-�i5:�[�Rl����:�Z/E1�5l F`��n[�dz�����P�����Ue��]�*�M�%�y�b�G���.Ƞ�u��{�/���W���<{�$���+�^��&n� ��BEa�D�)Rb���W���Ӎ��XT��j�p�E	Ӏ��V	w83j,b�w1���5�<{�T`�U�5��j�L(���9�4ݙi�c���U�B���)�Q�����vN��F�؄Y��U1֜Q���\�����|��﬛E�<ZӳEÜٻ�����޽�5;v�PO����e���6aڝ�i�P�TjC���3�lC/�j����`���O=�T��(Ν�b��n+X��}������c{�$��4Eo�^Gt:q'��U����*����w<����ٴc˞KϾ��}0�;��Q
z�>$��'A�|�����:1�s�._R�͛�����Fr�\>�s.��B]ї.[�n9_�����-�$ix���k�|_��~�R��G����d�!r6��6�~��e�B�)��ԐTI�S
v��A��4���(,�n�pu;�S}�9�(D]ՉE�A�i���2��@�BV��v<LY7H�BY[�K�%֟Q��f.�e�m�i	f�\Y������Jh�1Zd+&1`绂��)g%
$������r	=)(ޝ�i'�p��_��5g�͌�	|z�� ��J/"zz��`�
�Ƽ�A��E�lOvN<���������ܞ��~w+@n70�[��$b~�d(�6\���؞}`l�Cv��)S~�������:���*�~3��Mg�w4�D�=��
���I��P-=�a���`�ܖ0HVk�S��$��f�b��I�'�nbՒ�C��?Ƀ�R�U��Y^L809>q�kNZ~�@�������ļb��,<�c��M�qfg� �Y��	'��V�	z��@��Z��}��o�����Fk���j�2@�3�8ߦ8m;�����"��G����t"�W;��D� Z�H~ �d)�
z�E�ģ�af[3$L،BljgP�-H�k�Z'aE* 53�"S���X��	�� f���uEJb��<V�D��HW2�'Kw�{�.z]�V[�l)\��c�]�8�l�ҙ��R�(�DP'%Nb����n���G���.�H]ЈY��n熮��2+��f,K��c��u� ��kfba��bg��A��#,�a#6&P*�^���D�t�r_3Ģi��0��eˇ]!h))x/N���F�P�V<|(9��c���l��&�a6w�6Q�=;�غ���Q�sZ�w���9<k�bY2��%`�
���R�~
/YwE���w0Ð���Y��MeU�X�%�A�zߨI�D���y����-Nܚ��WJ SA��ݪ���E�ߜ8�g���=5���H��W�N����^s�5W��}莢}�|T"�U��8Mfc"�馛>��_���{�Z?���V*����[vl��O���ϟ7��7����\V�T����vۊ+W����$"���?��3��~0 67�_%��*#7w��LF�YNy��;Raw#&v��b��0|�?0��ī쟐����7�������[ny�{�kwܼ�(}����\p�:0��Z�LJ%�99��!�x���.��.�z��Z)�j}�B�؉쳤��s�Y�^ P���p3L ��ٟ������L�����Tled�MN�[���S��g���������[�*]z�Zm�XM��&X��9��S�g��m�6�5c�y�y���Pi�	��0:���,��9�]�������	�1::Z�ho"�7�����o%Ś֡J�}�s�K �Ȟ�ȭ�=m�]@ �K-\��)B��ՠsZ�ꎅbY��(X��m`M�P��.^$1'�$C��먘��sY���HmŲ~��	qփ��:�ln߾�?�f����cddv��T�^z��`��\C̯u-�N%�S!��BbMJ�jM3`&K2f�����![M�����?��X�r�"a�[7c�� ���j '�V�P;d�����s�=w׮]?������4��~���z9���O�!rLm�n�؜��<@�;v��dК"�+x��>���"̉��(Mf�;tɦ ǻ�է0#�Q���^�{��<*�m���Q,�,9�Zd��x��Q�t-�$+����F^.̉E��d���HE��2|�N��s0��$
��Y*�DU�NY�l�������EJ�sJ�M����v���&�}���� J�>�����8>>~����"KŢY�&7j_�G���ŋ�
-���闿�y��o��w���e��`���c�=�3������\�/��A�����44m�����:���pd�,b��-���:��3aJgv�r���	s1�J�X�I9�OP2JR������楨$�:�i����&N���|O����0�\̴����s�g�u�ӛ_��q�F���հfa�K�.߽�����Y(h�y.���x�����r\���3�8�13�/��/��A�f�c���*�6l� ��$�,Xo�*���8�%���ղ)�F�2~@0����A��vf���3[�Il�)�Q@0��]�.��R�ߙU�����ɠO����}�ǈ�NU��R3?]\`��9H�����Ca�������}����ګ�o��sv��ܹ �w �@D��!Y5��qO�4��j\X��#�d�Wi�k���+�9k4��+��\Ҝ��:DZg焴�uM�pfP���4~�:a�W�Ufx:��P�
ʁ��g��^�_���R�����iQ�����x�i��Y`<�(�3�G璬�a�[,��חK{Ub������9g}�o�Z��Y��w��Qz�X����4�!53-"4S�ˊ�{�*Ғk�^%��GcP�c�Y���P��ia�jC���4mϭiX(	�l_�O?����?p����%{����{�����)��;��ƛo�y��}����ޗ6yNg��e����T���t�q�sϖ�����	#�a:�s)����%c�"u9DY-��#]��QvK0*��\��99e�c3��@��ZT�.a�5�f`���¬ݾ�w�����M��+���R�oϞqM+'��^��O>��ɫWk&/%�{a�0��.XE?�d(xa��F���~��H�u��;r/>�yB֞�ah�'�GL؏�߾C2K��� 5q��?�� !��1Տ�Ƚ��u�ng��Ej��wl���V�?�4�ݘ�WS*U�/�)�+`Pb��$y�� ��?0!/�QV?��b�WA';&��i��1�1/���V+V*�a�'1��;9��x;v��m��vl;D&,�%K��M��犈���8~U�H�bS��*(� c+)m�4���9K��Y���;.�D	��ꈻ���� �˒\�����4� �l4ڭV���WO�h6�Y�SՋ0����&�-�2�,[�u�&v4"��I&�T���g�yf�VӐ�ʍf���ܾ��g���N��$Z��,f�z�����B=�]
���j��#61�(T��{�`��j�.$w�R@�#�Y�mx�
m�e�۵gtJ3`�w�c� ���
�-������<xϽ���{�E�M���{^�lk��	�n��^�h.�[�Di�O��h�X�q|X�K��{�L�G%+������h Zp���T��<c���������Nو�TRP2�_F��$%H��߿�_�L	�
��M;�r�R��-�U�pq���Y%I "6�D�lh&��Ϣ�Bp��'gvQ�6���>����v��\`�p�iB��dl��⍺��R��90�c�alZ�#L�n5a��{X��A�WETU ��@���(�b�1,��9дx#t!�7hGMXV���;n��h�pk�0���,�aj��S*i����w�۱e3��0�Ys��)�w�߷�G�x�����V�6�x饗tU���;�gV�p���RAC��ThY�#j��'����C�������>ٹ�;�Ý"�-,9���U����K!!U�� rƒ�o��U��,�n������i���YyԀ�:ю�Vh�Y��P6�a�/�xeMsff]w���mc�س؟����ӣ/mi��HJs��x}f����o��{�~�p`˶Ţ8�ol��'�m'�O� ���Q���Z��D������T*�M{~O�t��'J����Y���2�#*ABm5(^͎S��͢��������#?��R¶)��uq��%S2�C��D>7�s`�jJ"�����R:���db4�@���Nd�-Iӱ���,K-�
��&b�KϛFd`q� �+�ϩ����=r�8bnwIq3)'��Z"�`�.�W?�Wں	E3���m1�N���$����%��Tc��a��bn�|x�	�h6���f�%�/�~P�-6&F�]	w�$E�sd!逸B[�P�'Q%�}�f�S�P�sV�C��a�{D���5:g���� @�q�v�ϓ��抏��N�(w�����k��6G\z�U�:���f�"��ys0l%�qr
�$���R�V�����#�h=F��e63��p�	�~H���3.�Ba��Y�)� ��*n����C1Ϡ8Z��k�]1Y���⿲|�E}�#�馛�}���:��^׭_�f��}�H�"+�^�L�ы�Ċ�*U1��p��F�<�ȹ�f+��+���o������ի�o�Mj ga�=�cQ��@+T�%$�|��]�{՞	��e�훑并	�4�}Ń�Ѭr�H�elQyQ�OI���I�D�T}��vZ-ؙ���������_��'���;������Q}�S2K�M#6���XWGc���G!5J�˹�%�PQ���J���R��O>	"!_X�T��oݺ��T��NL�� �`������Ȃ�K�63X�UF~����70� �/��'��5 ���>�
���	3\I�Y�B�B'�K�c��j[m���w`�ŀ�~��[�i�4 e�޽�88N8.���'�j/&b
kp��|�H��2E��9��Ich�.��R��r�`yG�(��!��B^u��R���l��Yx���cmF�P�}lrr�nrY�V�-[v�5נ�"� �w����8����Y��p��\vd�cA�������Ie�#'",�`�鴘#*�j��Q�h�	���c'�#l��ǧI-`'�Hƥ�}� 7�����z��o���,�چ��rIrsKpNkjvժU��`�&��@z0hS>LUÈD�D(�& df���������{zz�V �a��Qɡ���C��R�
��(�9fw;YY�aV�$���G~����&�.�I@��;�aFz�i�1��y��$�0RV���`�c�����Z�D(&�������0Ϟ�@cƖ"dj���םµI�!�d���;J���V'��P�CQ��1�����j��XZړ���{{�8v��� SML�._���R۵k�7��>:>��SO���s��,��f�
L7S9z��ӛ`z2h������u�р�ȡ�P�MD!��H 1���d�(e�ll)�]@��G}��enp����k�T��֪Oĉ��J���Bh�۶mS���`W�5>Ω+��MY��?�|���l3j��ʻ��0��2��Q"y��9m�d�L�����Aʲ�P�f�*�TM�9u�ۿ�C.SSg�<\��/\�x�'���)!���{��رc�������X���O�	�Ta�〈�#vᛜ ���OX	�ydh�6RS�f��aÆٽ��6��'�j���GA��E�Ն(+�^�א,�}���ܼn��-��/��b"�(0�$���m��"�.�Be�E@+�I(8�5��+ё�ͮ�\����q�@S��8+Uby��;��
e%䔺�ҜߥI���'����!�ʆ��7w����)�8<�˺�D�������˯�}>�c�!:��;�.�8R�v(Ewd��NR�
(����aX^��f����7��I%v�#!Sm<����>��G7Wm�5�=�{C�:��+���~��G=��j��Nҷ�4�җ����ç�}~sj��hx�����O~�ӟ�3\̆Aܚ�Dש�U���z#�U۞[5u9�-E�պf����{12��g��z�������>-��"+���]N�6$vT���5��k
���2	��5�[���Y�uwV��y�a�ux]q�e��8��u�A�!�va�kR�5'Ǖ���B�������ÿ���?��%+�tK��U����V�E$cc*Xr+[7k���j6+�,�8�x�9b1���a�C̅�Q�(r��B�I����|#��,|o��L�m"nv8+�T�tұ�$��;� ���{�!O���d��q�`��g���_�zfrԶ�U+W�|�1�}Vju�SI__i��%ccc�M�u�V�eC���c��[o���_/�\6��Ã>eoW*u���cn�k�����f@ �LD<55��3��DNY�[�S����t�᫔�P����WRg�h�$4��q���z��qb[�.BUV��6z����d�4�����`1��ҿda�%p�f�BK�}ˇ��;������z�	�M�L̮�����I϶K�>8��o7&v�R��"�A��vzXH*檩�}C�U��JM�%U���m?�"�������tѢE��~�P�@.o������љV]�ے�o�\[Q2R�[�716i������1{O;���.d{b2n۽f1�ɐ�zubY�鱃��pc� %!7ə�Ƒ��~���I��SH[x'Z? kH��u�C�ͅD�ؕ<�����%f���W��7�(���E��U��l���ɫ�0ьE���>Z���jb�&S��{"��Q{kJ���k�;��`�� �<j��Uh�gw5�D8��Jzl��z6!G-��T��z[Ðz�{"�|7� �Iw�:�X�a���sN؈�Q1�)%}10�/tl��IDX��檮�|Rw $@Sd�1�hpqx�(65��	ʪfa��Z�� ��״8)��d������t�?3#�=�6��E�u��z�睰Zu�=�<��Vmp0*+��S��5c�%�t\�P���J�bb��OZ�gB�U��UK�1 �̘O�n�,�H���S|z.�;���S1u�G6����Ls��0�������0��O��C&�p�7)_1��"�-n�
M��QF�@�4N��Lv��᠌��6���ý�{�m��l�Ɲ�s_6T���vdk�)6(D��1T�Tr�M�1�0�^�A(�
` �F�<P���$�
�N��E^cz:01���sV�-���o�
���Ο?�z������wԝ�����1a#?��$k����la��d�@���^�78���Nk��yvc�"j�Ȁ�[�a�=%���$�_�o	�D��K>il$������;��wW��ɛc�����ܛ�͑Ԇ�P�U3�gp�/�$���FZ�DeR8�t�J t�I)������=�9 �2��C7��4l���ل7���@�Y�Q�*�(G�}F ���ĥ�)0��+k�drS=n�J�k\A�b���97���Td^r9˦fo����s������I�9����B����iP.����\@~CKϤ.���OF^������2��ɸKaU/e9)�e�/�
Y��!�o�P�3�N
�����*N2��Ὀ��PV��v��HM�H���<�z�u����'K�,98v^�G���mw��n�	��կ"��ǯLEa���?M/aN� V2���������g�B�.�Ξp�]����������7t�,�N�#�,X��f h!�����H�`_Qy�<��;�{�$g����l'�X�E�g���x�+V�AY���?��;��;���u�]��	�Q�bŊ'�|��z�k�L�\�����e������kE]]���n�6h^�z�4�ԅ��TĴ*Q�?�V�l^�SO��m���^���(���s�>������)	�z�ŗ,\��΂s�TC��w0Z&�C-_Ȥs� ���`_�?����v�;��$�X�=0����`3���O?�W6�MK�*�n���K�.M{nГf�>��1��2�q��a2�:�v��-*9҂|q�V�D����G��)��ٔK�|�l�;��Q7��?���z�,X��K5t��ܹ��[o�g0*�s5�D��z�'n��6���ԺG�"� |�d.Wd�À!=�����M�6y=�U�V-fax}S�`�jz�_89�YI�A�5�͑�b�+v]����'�^���W^�~=|c��������f�Ћ})�����W6�8�{�+J���82�����P��V�qg�e��q0`��p�~hҖ�tj������xf^�*�Y�8~��5��g��у$e�|}NS����
M΢R�H�Rf���j1Q$uġLK+�O�q�`�����peW��t!?�������k30��b��0;������$����W���y��02X�YT�'��iX��r�ٙ�>�2K;���q��w?A������sƛ^x̱+�a�E�8�1��kP�Ǚ���p�մ����WJ�Y4�1���0����ę�D��R�L=_��[G:�T�Js�y�\�!��,q�;��z�L46ES��>��>����jA�{�l˝��А%��6+�p�8H0���\��N�˂��Exx�<��N�uS��F$�{X�������K%k������)���9_�x9��ux�2��z������۝w�y�v����
�0��.�By�!(���짰�����{'&&��������/�x������/�|ݺu�@"⚝�yXV�a�v��59�V����u��<�Ӓ�j���a���+�"R�a?��E��)�9		B\%�<�{�UƮ�|�_1.���R�u����%��
��!ADb�c���TXm�:b�P�L�8��E	�V��:uy��f������^Ț���S�X��C{���Ŏ�0�R.u�	��o�(�3�S����8̚�$Y�����B��P�CKR<�3t���5�On #�@�؋��=�cN�ϣ�}1��x����9��S^����^�~�3�f)��<Z��k%�W;"0 B�R�Ћ�V�#�Qz���?��ǲVx����<�u��u���65��Xt%ݔ0]�S��v����M=�.�U!��y�׳;FRm�Ȳ �EC,�fG��|�_��j��J$.ؖ.E���A-�"e��l S6�4M����5���MIWqj��O�ʻ_]�4+����ޝ���IԪ"d���Z�CG��`%nw�f�쀽p��\|�_���/^��:�� ��i��r�}�?��W�][L����04�m�������][�i�uHі|�7���+M�i'ԄI�X�!�B���vd��X!�U��!��-�Q�S�hC��4�)Z�P���c������;���_�L�_zie�9�f��#���|��(�qP.Y������hgS�l@V����L�i��{����@�-�v�?���V�\�l� �ڴ��g��z�����$��x��k���m+T`�^��$��U�Q�&��%�!�c���Ή�����qXAp�u�S��"q)؋Iʺ�`�P�Rq���|� /T"G��^�N�,����^y�	��*ŒL-S:����G�n��O6vn}��b�T2T��\��U��A��q�i�׹U)F�v�C���cC&��K���/v�M�4xk�e��8�Ԑr���e˖MO<��b���!�=r:J��R��vG2���sF'w<�ܥl�����;mOcLR�ZM��]?j����{�=�2�i�Jٔ{H��lt�:L�$y*|){8o�f�� �ڮ-K�!����X��)���L>�a#�3 -ix�q�QX>�wD��Kyb	� �KU�"�����@�-��DD(,siC�%}�0����4.ad�`�W�sť ��M(4+�I�-{��^�u�1X&�OV���3����#�5b,�^
9��{�'�~�ݶ��i�� #�n�b� ��ȇ���fLRk(��3a�$d�-9k͝pS@ȱ�8�:��܌�.&��BQ��(j,jB�
1`��$��V�|HĴ��L���~��&Q�[���ML�IT�����^L:�@�(6�EŴ,��@��u���p�i>�ғ�n���2�S�/^��h�����M4g���Z�g",��6�"��{&��n7Љ�I���'����Y�~jĨ8ñ��@oBB�!(i�a�O5ǧ�vg��A8h� H�=����8֐�J���X����DI�,ɶocE�D��$U�!�!�����{�"�H���˖����}0��=�	t���;#J�����C��m+��b�ߜ��n`�5Hb
Dx����c�,譖Ao{��S7�ڳD�1=f��c[0�+w�䄜�������A�~���Ȝ�fk��唓�rS�>�)�)G�X^a���C�
Zpv��u�0� �W=N0K 7�S��h!��s%`yҐqE[ł�r�̔fD��ؤ��l`�
�W0s=�,�EVqBX�90bd��0N�}��/���Շ�BE�IV�0�ZP�Z�&yӜ�����@�x_�y;�,���(ul��Kg��WK(b��'�
�r?Z�U�f!5�Y����S�
=F��VO�^�^��|�S�R5ݔ��9�A{;�"�t�r��FE�F)��m;��y�%�̡b�퓙c:��	�*s�l��nI��QSw�G?�:�t:+V���ܰa6�"��(XV��vڛ���u����]*aC-$�j�y�k~��իW����{��KD��6�i��K~��m۶j�*Py���l���ba�ɳ�V ���5ګ�Z0���zT��/��T�Zc)G�}�N�#��Y�.�:��R���ʁ-8���N�����Y��y�7\��;��/�2g傓?��|�[���7�q饗�K5��(�8�O��`�~�3���c7��2>�������k�!nʪg����)�%ʇ����E�r�?Hּ�r�u�m*�j�f)�n��V�XGt:؄�7�SSS�Vk����b�V�����C����m�300 D�Ku���	�[��[��j�+��>�y�\䝕�`H6l�u�\��C���m�`[D�lhâA�U"�m�Ol���<�"ۺȵƹ#T�@]��R��w챘���O�L�ٳ��_<p�@<��]Z��|�V<�=� ˲��9�"��y�ND�|Bt:Y*2�®Ξפ�.l(np�I��K�Ee�k���H�""�MM�H2����0����|:D���Ф��ʓ%�%VJ��s�A$��ɛL+Z�Y>5canM&I��<>�$���Iڬ��TM���|�K=���7����_M4��ELGrz@���q�l��\Uŋ��,�ۊ���<�<T�,żF~�8Nu�a,��O�(�V�����W��b��PeE�|�<lͰ��� �d����]g$]��e��6M��u�,e.�.�IJC�R��8]T}�ZTd�!���K�	�}%�z���t�o#)�u����"0;�
0�S~rr�db֜I ~�=����тtg�GbҎ�-^�D7j⻫�h�B{}z�AX��^,�Y�i��kqu�a[Xj��u�%8�)�����$sA���A����MU.+:=�0�m-�e}�ݸ*L8i;�<�ɲ�Vi� W�H�EW��w�o2&Y7��1 Z�r��FÏ�Y��e��% �۱c����8�fƂtY�Ur 
4��F���
�ej�%��4���	�&Ƨႀ�P|\�:Ɖ֎N��b044�jc'FʅD����J8�[̵�K�Uw=��E��V~$YcOg�#-D>QZʷ���ජ�\��C�����
J,��ȫ��k���L{d1c39pK�ؿ�,�Z�)�N�lE��2�Z��h�g�R9�s�N�d��f՛y�h�!���N3!3׶��[��a�.���9��K
	�v톬��3O���u�L�s�
#��@���V�b w|�kN#��|<9��*KH�l]� �h��.�J��ƽ�THw|�W�4�uHR������/������q�c�� $欳��ɝ�=��'�v2j~��y���܋+��蚇|Y�O����GQcS�۞�+9������,^s͵��܎{������mc=��P��(�j�M���_��w�z��Z��������F�n��{��h�llߺ���~�e�U�%��p�엱�*��!o�l���Ʈ��<��vQ��\Kd��Y�C��8ܹ� l�#��/"%`7�q�Z:(8[M��Q�٨��,�qܱ���UW�t�M�T)X��c���������]84p���{�D�~�3�?��J�z��7� �&�X�ݯ3�`�Z<bjgR�sJ�:W!���1-HB�(_ ;�H9=�a�H�'Z�>T��$���ā�ى�V�h��}`��V���&&f@��dh���Yx�[~��J.^ om�Ȃf˞��*vCR\�W��W�?px��T4gf!�m����W	�r�I�-i��-{w�>��Ӷβ��Y<��o`	���oN���@�{#��A�� �����0�x�Y��.��r�A�t�`
)L+"�HAg���0�ͨM<Vt0eO���=�D<	cΆ����<"nQsqo_UӶ����7o��
���!���J��eU$���m���bO��b %ҍ
V_���.�_S�M��O��c�i����|WҪ/=����� �-Z
�e�o���5�-8����6oٲ%��m(FUV��#D.c=R}Ǘ?hF�F]�I
8	����[��`lH���0��Ċ��f��I��`���(�~T\�/ W��X�`��Y��a�-�|�f�r�f�XIH1��f^���WE�
Ř��_��r���V�1'L���>��OOϰ/M;��
�mV2�
Ȭ����	����O�{6�*B���f�T�-ש�'!�r�<==1l�B�a,� a��S���(�'T��:T��[H�)�d�o��d	Խ���i���ZG�l�o����0m���v	>:�S����&{`��KK�J̓�wQ[�0��.�נ��L�A,��yP��"tEQ�6�N� D#ԍhˊڿhYX`��`ޣb����X�x1 ��{�-d ۶���mo+/_�d��o���U	�]�Cɧ�ųNA�^}�Ν��e�����b�=ֈ}J������vL	�)���p'J���F��_����1�&˳M!��C��8���:��O�C+���"a�����բy�'�oh�n��nblqc!f`g�Dø�@�UlI�%�<?L6J��ޛǀV>h}����)<*�T���K��-?�ٽp��1���$/M����q��g���?��"P�����KEc���z�UN�*)��z�m7a�<�裣��;��9��]}���K���ʩg�;��5ϼ�;l'��X�]��N��Z�Y�+p�X�&���\{IW]n�q~��x%������LX:�Î`h%E��������epk����_rI�h�رG����?���S�O�aw8 K���Z'�c�+W�����eMu=�",��7�s�w��(�������?�1��P�<�H�0��r�1?�駟>��s��^q���'ť�#e9�9A/vW�%C)NZ��ç\�����j.rФ糗<���v�pë<�)����p\���r��>>z�G����tA�8�g�5]�P��o���7���?Z�p����~���]���a�*�~��kׯ_ߺ�֬Y26�p� $\�x��n��ڵoh��n�1g�I�X(�fȩI�yPNҰ�$q����aus6�#.<����J_�E]�ӻ���͛������TL�gŊ{4?���תXT���N؈qB8�����;O8�X��2��/n۵��?�9�-A ���h=��o���������}h�����4���`H�'�n��7���.�(Q4%���a�g���EY�M��P�2ʜ ����n��\�!:����4_���	{�Df��2q`�����}�;���K1	���p�s�6����\r	��(˰�R���6�j2V�b9,1���O��j�s6��W�8�ˮ��f�m]X�E^1�+��X�J�߶u7H��s]/#O�y���)~ql/r�gG������˺�Z��'&&��Q���gjQ�8r�v�8�+	���LNN�)���"���>VL	u��8%Z|��7��."�%��D\ye��az4���W��:p��bp�^<�o�>::
���ݍY�-]���r�[�!�.�W�����&!�h<fF��RF�|�3��`��}�4�`�b�����~�?M�عc��	���.U/�}Y��bm�v���Ѝ�x^0/"�Jy�0� �&-�S�a�s{(�o$W#��5��ż�a���,l�TCŻ;��q<�����X��3�}�ve5%�D�P8�
�VC1ۚ��P]g�M�q���\���*ן x���(�,�.����Ƿ���Q__�l��P4>�,��W1`BRC�߂���u�%0����b��W(����_W�v0i 6`#m	=G��!I%��D�Ƒ@Z�jߗ�t�.�лV���j��d�w���̒���6��7]���;I��˗'nIY�ʃ���!�4��c��X|�c��@ʘ4�k$*m�[m�G� q���H2i;��y[���l�7� �,ԬRr
CW�Kѕ=��qӲ���Lo���9ݱ���y���Q�,αV^|߭����~��\� �6�RPk�ZciΗ�J;M<sf��yI/�M���q�7N�b��Q������*�Q��d������)a}��Y�����A<�������銈ӖG��Kl���hA1��u���4�t���ԓ�X�)�|)�����S.���]dQ/����t��˷Fq��}�P���wl^��<��9\�P�Q�p
�������=�\_ƣhQ�m�+�`n�Կ.��߿q��U�V+�p�Į�Q�T�2�Ⱦ����}�S0�	�1䇺뮻��?��?��g>�K͑��F��\v�e�(�vp���x�I����<�����Q,�K��Bcn>�j�YI��.2g:����w%AN")�mY~rC�#+��;��:R�x�E������Ըa#����K/~���ϖ-k<ҭ��z��~�<��ӱkH��z.�y�;��f����p�y=^�`���a�a[Z����צ��;�~��92�2�����4�ߙ�����=S_���?��_���l����3N���>�Q� �k:����\����\ȡI�&�
����ك=.�/����R�K/�+��
�9S��`��c��e׬�����ۍ<��+�x�g����_82ݺ�����o|�5�]��D�tD���W<آe�+p�I������H׉�-�=%�m��/S�:�ܘLU(���+��Gr��k��mS/�':��d0���*�k�ͯ�����;�����^�tםw�>]s�91,f���^�jÆ�Xۻ�i"�j����{`�("�x�c !-�hMB?A��2���s���D�}��V<�X�$�(tk�a�!���&l�Tk7ۨ��i�A�L�M�ͻN�l�`��A����K$Tdy��DSӓ�F��j�{�����m�%����� s�������KZ��r�Ԙ�M�D�C�:T#��q�zd�"��(�Cl4�$�+�DZaŶK��F\w�v�D�����'w![d"<��Ť_��_04��~�*1�8���$��y���~�CA�4�]t]+ZI��BT�LA�.RC��
&�)�)`'F�H��Bi��p��-�G)}B�lZ��6���ʽ=��o&,_����~ɒ%� �0D��'�u�RA�Y4x��A��Sa������gFg�Hq���u�K��U�5�&��V�9�j�n\qQN�T:��Lc�m/��~0��@I`�%�	X�Ģ�@%QC�X���h�%�D�$Y�/T�"�������>�H��Um���Ͻ�<�#0�1e# ��V��̂U��;�i��E��`�|�`�*Mk&��	3u���c��Y���~�~�1�*��@��ݻ��j������p٢��319nj�[�W@���дU�f�=00P-W�N�hhDt���p�eK��+ŭ[���Z�p<��j{a02oLikf�	Q�p��NN�G@:��*�%�OOO7�&fq����k���RWkp�vY��_,�/!N�׏�m��)��a�.�i�]ϛ78�L���_V�U��t�5��Aǆ��[�b�$���8�t�@1+I��E�?kup5)��"@�n�|E����g���F3�C�Kf1l;��~� -0gX$ӎs��'�w�Ec��I���O>���ӳDq�����p�%���Ɠ�=��zzw骆4?R�GĞO
�yJ#N싉�3�7r4K��(VIaabj����4sOP5���gQe���u�#�z��!�^�h����	��b��Ao�dsV4���Q�a���6���"�S� �F��T �w9�9t驸��[L��y�G~ ��i��R���*�W��x��1����ٶ��1�(�0����M�.Z��x��0��=}`��ȧ%iܛYA�Ʀ��ؚS3��S3��'��ccM~M-:�fO�o��5Z��IS3�
TݨԪc���s�K�+���k�x#E����fn�K��B����,y5{#oҡ�F��DV�w:/<����oq�������Y)ot����So|�o=�أ���|�{�?���W��ݎ�h
f�GA�����n�ʍ?��`v�ثC�^�,�D3���c���=��å��r�-�Mv�7~��_��_�8��k��:ɇ��x!�p����@�!7���	����f*�O�D��O]��XdP*GD�M�5*ô�+�r���hW��A|&��<���pJ�g%�R��������q�`���5r�W��կ|E�la��.ޕ���?n�`��L� �;��3?����|���y��ccc���V���S���� �4]q�N�,��oY��G �ٶK�MLu�`Di����C!;]x���H)���}$��* s�?w�z���/�����'��i4�QMô=����㷽�Jؤ8�>���\��"�]I�>���}�S��|�v�ڸ�e�V�x� ��%��x�E^�����w����n���/5t�����'>��+N�
���g>��O�~���1�؊���PO2Z�`��������i���s�
{>���9��]&��ń�
�4��o~���m/A�96~J�l��}��}�EŶ�~��I�Ì�I��:VO�4�	a�ôf��e��}�y�^Z��)F�GI�O%�GU�Ē��#�Y��9���Tp���L��+���D�Z!�s��X��$s��u��\�+t?;`���TƊ̥+\7b)�Q����JO�Tu��ґip��Ȓy�[ɿ�v�� ��D)�2U�H���\��d���1�Y��>��1����S�Q�Cx�@�Τ�=�{��4���hyO9
)G��'�,i��W�\��l����Դq��#����N��J�3�RL)���Έ�j(�F�],b��=��w��u� B�ޓ$k.)�i�
wfqWA �9����<�0>s�0��Y��`)� ����2؞9���ÿ�XȑFL� n�����X�s��Yq -��]H���g�
�`���k�����١Hv�F""�b�,�v~M^\\�������/��T�Ac�%(� 3���x�E�8��h�5�`̥�����͚��b�lfBZ^��,$�T�ǍC��+:L)�����ШL$��%]�T���<Txn��q�s]9̋:�����'''�B�m��{|v��2��8����ۤ�T�zВ!���t���L�Ē���gf��:��J�5U���K���*6w{��E�I�6�E���P��<vė����rr%��I^����BD�xe��梪i�B-�e����=aerj{K1�7111<<<44Ĺ� �`{��{i(�8	�,���5۠R�z���� CL����CV�:�g@����'�[o'Y���"�s5s��# �Ua���+�4���}���/� ^�&JOO�Ν;�}�;׭[��SO]p� �l�`����n�w  Q������3
���}�-���l�.�ʞ*���w��^��s�='�>�(1R��җ������s�9����^����>�g�^`8/��7޸f͚� sK���P�H2%r��J�iE�Y��|������W�� �e�����d��s���0κr��NUT)kў�/0�?�!~x@�.�&�'!�#��������'?�	��[o��ꫯI;���LJ_J��q�=������ɹg�0[n��a�mߕ��}��֫��uU��q�c-�m�)K�4��`�(�h�s��0�H����$�k��~�$���%|�..��|0ePF�,8}�$$���D���Z΄��*ų�\8��ND��x�0"���_��+�e��R� ���o�$�����]Vd��"SU�]���iA;�a���������D!_�����1580e*D�mԆb>�P�J�8JP*����`�
_8:Ѽ"r��f�I�bȖሆ�H&�����n�X�KS.B�Vrq'�C64f���1��`���w%g�J�_�f7z��3T�HC����++�X�"�[���e��`�)�^�qKء~"� p>���<q=�T垡ϛY���'6np�i�P����`,EAM��e�>��E�i������j	��>mH����myo8e�A)L�����`�/��|���$a,�裃WS�LU��ʕ���A�e�"aO)���E~�!;�[Ak[`>>K�aa�Vj��b�� rY���4�(�2�4�L�È�(f�(%�@摒����ãx��C_X�	/�	�� &N(�?�Ծ���q�1��B��5�,`����Y�)6��)�)�q74n���\O�����if��E,�U�$����s����ΰ{�ԠA;�L0G�4��&ƮӜ�;��; �E�|��9��,�>`ÎBSS#Y
�y��-������sT�|H�Q=	K��<Qc���g��%%6b���h���F�+D0P����zd5)!,P&��5�!�-$]��l���U��3���%�r;N�\�����
���x2t��d,D9�D��R+�J�	Z&�R,�^�L<�{�UX����`__���228&�7_�
��_�s\��D�j�:Z���t�`䕂Y-Z0��S/Ã�P�6�j��E�����(Xqny��s��U�(W�3~W��a�O0���C
6�-�3�a��BO�6#.-K=��h�B����-]���J=~���&A�Y�ȚkM��%�􃢀MA�
��ŘGdRTZf�kD	���\@�������u�`E�HF��҂ť��'*��5�~G�L�F	^�vsrR+�_��.^ i�<����:@�0��&�@C��UXSH
Cq}P��ZNϣv�2&u8/ ���L�8N묺%��l̇���g�E%�Dđ�Tq!稫�͐	�L�eۋ��{��t�	<L�2��;����~�����ף�7,bt�� ֠
'Y�b�K^� љ�wm	ٝpU�L�>2E΂?�lgVh	�Ndʅ�jE��,��{�f�U����U'v��	��Fy$F��d!�Hdc�a��~WƗK�	|��&�a��L�MF��%d��H�G�&w��t8}R媷�����]��������9]]�j�k��5�[ȁw �Ӆ��[#�e?��֣�9vr���0�7[�q27\�9��x�Z�٪=>>�r��_X�y�C&����H��`�]�����vb�'��|tW�c�1X3���&�9ù���z��;ңh�3bF{$�a��Ҳ�l4
'�rޝ$���k?Ex>,��h���\鿫����}�w���_��W�E�0J&WBo�PW����_��ػ��ӻɰ�ƴƙ�*/̼(�\c�zN��5+^}�:�ng��B^�HM'��V�g���v���?����?#�H�����%}������ox������m��Z.�Ef/{��^�K_��l��S��oZ�Đ�TS?dX5:���Ԓ��*tZfeT��Q��U�^P��&�� Xu}�м$�V�M�!���.�H��Z��'�>F�9���ZAz�)fȥ�:������.������x�e/{�{޻gq�����ӎwm�BA����o4�޽{����n���P�i��o�[ ��#�̄�D��Zca��[��k��`���i4�������k���B4��%Y�]S�E�xC?xh%qV�Gr����V�$�/�A�zb^���=%���fX���[5�P�i�ʔk��k~Z�\"9Z��'���/s4!B��Y���� �+��:VY�\$��<�*D�U�AN�9b>ϑb��G._����о*bIqr��s�0ei�㴧NL�q��Y:<3i�����b:U%�.�� #�e[�ta0��t[�VF���J.L��+���(�"��-)kI*�*3�ĖL�[V�������,����L'��*60�ɴ��WR^e��=��ХnI/;��=@s�fn�ٳx�'EL����\��k�}�h�QR�T�J,��%�Yl����-��Pw�a�L�CG�ء5쎱-��xz��*X�.��%*cr�I]"=�p|&,�w�2a}��q��OM����G�6��-��_|�aʌXR&��,4V�L�[��%ETR�$�I����8�(�dl����R+q2�BV�{��P=N�Sl�r;Xf'���$�Yq V3�j�b^��>a�eN���OJ�f$�qk����ȃ�2�@B��IB"�2{�x��q�99�s����ͻ��.2%��__;|�����b�G�E��u��mHo�4XJ��1��Z�
�|�O��|lllA_l�ۋ�f����1e�DU,1;mh\�Z�J��!��/*�I�����U���N�Z��g�Ք&���Ƃ�)�X&�-2�r!P����F������$r��������%iOU���ɩ����(ƒ1�+U��Sݧ�[�.��əs�$݊������M4,Ut,!�3h-w�"ZL\�2�����*�G|у~�(y	������'��5$a����L�4�Kk.��r��z�cT����(����J�ﾛ�t�%�P�Sg�q�u�2�+�Ye�λ���>ʲW��(-LBX��>M�T8G�r�t������c��?��ȩsl?�e��E���W�W�����{����$#���Ќ����������R~њ�Q��lÌ�X=�c�������U��H���˖m?B���ŕ]5gQu0�+���T�sX�ӟ��7��M���'����v�m/x�et�Z4�Q^����W���c�����<����Z�p
:B9��J^���]]m1�P�7�u��Gao����ߐL�Z+0ceH95%(�zl����窑��)�$��m�)%,sZRVȇ�~T_���UZV�����\�F�J�0��~dI�\��Ġ	�5�[+���J���~�9@����������&�f��3�S��\�4c.Z���e�Bs��F1�����v����3T�#��h���Oj��u��/̆��Wǥ	�v��&"��Cku�٪9.)h�p�{C�/�1���+R���gI�:��#�����"cj����<�Ho4mԔ��;V�q��-?Ki�CN_��f"]*�Q�Ѥ�`�!@�#�M��8E�UȶO��`�J���N�&g9���*0@��-Q[ѥI��<[��kER��q����R�Q�9ʊ徊ś%���a���~���7�)ȌI�B�J�J��[^}�~�X�f�c�g���AXKY��Ү�Όe���b�p�L��6��0�;)�u��|ŸE꘱F�fwN���|X���Cc�
p�d�\Xkr���,=�a6�����$A�ۡ��Y�� f��&d��A_d���J�D0�{˳��N���D~��Z)��p	U�S$����qC�д�����Omw����>�i������X�~�`72���u0��_L��A�|�N�ʫ��0���K�Cég~��tQ�ҙ�4� �pnD�Rӯ�`H͋�pc4���1� NKw���@ru�C��=uu��`�ŉ�!����	�'4��h]QyL�8F��x5N�n���[zPw������ȃ�;�/?T���ah��&3����Vf0>����Kgߐk ���(�dU�;�T4Q�/�D�i<���wz���l�@گ]3���YbXfjDO�Mٱ}�#;��U�u��`ȕ��M� &yQ��Tb�#TVk�#��5	c$�@U�
	��X��"z���/�k'�uY�_��Љ#��p�1�N�h�������{l��\�&�D�~f�"fH�C/롡��LT�ጧ����aE��#�I3�7S�Vpm?$��p��.���~�#��&=="�w�y'#�T7�S�~��|�ώ�E<��k�X;�o�O�{�4�㹜FH�,��L3zY�0e���Ѫ�X�!���k�&���Y��5��A�[�31�^���XI
c��@h�������eK��%�Z%�/�	��Ȋ���*���A��si���D���Cy�c�@�C�x�Z�&�}�r9�Y�tI�:*p<N���q��w���w���|��/ys҉�R�O�5��:�޷��%٪5�%��d@�H5gE@��5����i�fN�A"wǎ��������ٞ��8�MˍQ���<���x�I�O��]�E��+���~R#���94�bUbQ9�� i+��?�� �?��l��������/��ͯl޼����>�����v�Y��B[�]���25����,�,�L��y0��9~F���]GI�#z�H�\�k>�,?����\9;K�V^V+��hL�b:����!=�s�2K6�>��S��An%N�'�ØX��$��b���PrB��,w�AO:8"�8w���|���Qv9X��>ec�LPI� <3~��H�V+�֗J��$�L�zM����u��%KKK�ǧ���399�nݺs��@z�|ǦM5�`L�\W����o8q|||���B��$�T�`�0/x��t=miP<�x�޽]�]s��8&�+V�����t��4ֻ�L�޽{a�os���.Ņ2H�]e�,۱ٽV�*?@EvWb-iP��8_�(�-���l6HB����G�.<H�+-o$L�����0Mu�Q��\O6�!4�U�(�[��,�Zgg\^��hJ�R�p� ۼ�A�M,OzN�la�kS��Z<�:���J����4"�tľg@�0-<�0�&	*�)��)��zݮ���G�.��'>W��3K�xe��(#!3)�G��77��aL6*g�hC��ymR����+�|��W�"*~PٳS�2�?0�r�q��SH�(8�DGE3��D�	��J����0���RF2ţS\C�=��r�i��+���+�/d����I�Ƅ�x�匴�Tj�(R�bx3��q����FDJ��5Ԙ�}�%�B�l�9�����A$~90�%�����$-N���4�Ԍ�qBy&�����Q6ط���Z�*;�O�b�����upCe�X>�@NgH2�������Ċ#�#��&$a{������Cn��F�v�E�0��3�'}�	�.-X�̥|8ϙ��'E�b���!�<��*,*hj�WR��;]�+���t�������"F���	l#]�٠��>g(qu
U�hk%�V�uI
����a��H�^E'.������`�h�A��|q&B�u/��i�9�ׯ���,=�>�`�T)��j=��u0@���W��$+��"��t}�FN����ɟ�!�ʔ��|��}��'Ә޻�QT:����An���g��ݿ�.��J��I��S9 Ó"R�����kÆ���pD^4Z��w�o�"@7��Z���K���/8����U��Z�,����p���+������6%L#b��m�ݶi�&�Ū�BP������x�)�\���q�Y��w��裏~���N��Ob�'�$w���ԓ��O⢧rT[y��%r{�����=H߬v�"gr�yR�1�5��Iv;�����_�?����-�@��8�ylY�a��~���A�^�?�B����c����\'y�'�0��������)[�	7��d> �66$]��K,��BE�Wn����`R��˜�Nn�*�ʋ*���u�ʌ�~ʉYA,qT����s����J����+*���<O���󦫪<�"OF|��lk�9&D�Ứ�8o��B#zo>��[�����{-N0	��,��~�ga�ۣ�5����N��t�<[X������Qw()�W�������~h|�+.�݉U�[ٶ���=��+���Ӣ)���q�􇽩Փ�����wz��� Љ޶Uc�1�3(�3�G�=~�9��ʳ/~�������p�F�w�ygw�HT��憣6\�җ�y�<�����ޙ��Ņ���,�l�q4��L�aB:dP�]ݰ[�&�"zFP��Zb��Y��0T^i~s�R���i�E*�A/�/u���C�t�s�("!Ҁ�-b�ՔA����<4c&�64�\�E�����ų(2�J1��U�3�h�/�g�v��1"v@�躓cm�ZZmR����?�:"�<FG�$]�v�jn3�{��̐���4A����qW����YI�	����7&��ns|�r�v@��	�&X�z.je�(kP�ط�4 �- =cYg�w��#^�9�+*Cu&X9S!��RRc���z͢�J�rMͳ��N�G��m��c�\WTOh`>��!�V�	���94�YN�W֣��:Q����n�*�i?�5[�]ٚ2sT#�.8��n�t�P��Pn�ײ8�kv�$��L�]۴�)WTQfS��\���	��=�"E+�7�̄ �E?���6��[#�ь�i�g讚���z�P�&��A�4E�ZKA�ִz#�&U��ؑF�~���d�σry02� ٦V��vn�F?'�4Q���*N�ݺ�����L�<�m�e�tO����r��*��\d��@�檨��փ�͋<���s�f���*Wi�8�Jz�C�GCq�%�ƃ�w��eR@�?���N:�>6�>"�>>r�fZ�x�f�Ī�0Y����CX���G��L���ؓ� ���Е_�^�����RU��� 9����ɚ�K���&�1��
@�F�B��p����c�cՐ��#C��n5!�h�%J_�6��J��	M����?�a.����n��A��e�-ì{53gj{=>��7R��]4�L���LC?p����j�zk�M����''g��|<�ߥ��}���ɱ����B���g��[�e�A��٠šk6ռ`^�t��	sX���( <D��x}f��r���S+W��K�Zm���;HN q��-���I����u�h��3��d��<���e��O�n���j�f/���'|��TK���?�{7�1�M�&N�vF`�N�����H��HٰHx%�-Cs��xG�*�4�S6�����������؄��O��Mg�6;;&1��Ӥŝ�nc��C/��S7�F�Gr韾��o}�_~��5�����ض	rc��i�Gx<g fת�,#��C�����n�X��|�V��Z6v��V�y�?a�~"mP���H��S=f�d���޺�c�+���:�����\s�7H(d���a@�� d�
��8b�O=��s��g0ȟ`�-�G�1ڈ���8�я�s/f��$�OyH�����K^V���Sy�*f-s���"r/%,l��|�p��O"A�xP~P�v؟]���1�4TJaA%��H][��k���������&��6��4�#	��ٳ�p�6t5s���l�X�v$�~��o���}�sO~�i��w=�mo{[���{���`	d�,��+]�wЙa¥�󂠒�f��#��`�ꊷ���O֍������� dkG=�$ٱc�Ν;���]�ض�L$����G���Xǅ���8ɖ���B�Z#�Zx]8���2��!�W|,�톤��O�t�dh2�� [zz�Y�������.�������U"&u��+	K�+C���Lm ����d~H��O���s$�����K�ﱗ���$�����?���(�� 99Sͱ�rz����Rs���t��J�Y��4.�S�FhJ�h�,>�t�Ҳ�O��0�zJ�II�.�D�ZH]����2�@l��� ���*D���J��?i��LXZ���&��η�m҉�WF��g�Hh�m<�t��$j�hG��Z����5��TX�x�y���j����?-�w��OLH����P*d8�yh؍z��J��9�)��!��CQ}��4)EƊ��"�&��:���ӥ3g�8:x��;c���d9�#��
Ù���-^�@�e~H�0+#gԌd��*מ����
���l��6�x9S��e5Ӡ�y���+�
�"]܎
?�H �:�L��SOF������R��m�k'��Q^�C1^J�j�/���I�V�Y��\�U�*(F�gH�%�Ͷ����A�f�N-��D��L����`��� c`�a��$5K�u�bsH9�^�|�|E�5�:�&�E"�ltQ�ɡ��x�%9t��o�x"3{��u�E�z�- ���~���.����\g�����*C�T�K/�o߾<�<��\1�z�5>�=�;A)q�.G��<��:���k����Ty�4<��g��Tν"��R�� Q��e��f�᦮)��@�;�?��k�����lh���`���u�{��_��� ;�/a�B�TJ�Q����寤a����l��R�S������Z��'�\��x���g<���8s-����Tٶm�ujj�~ݱc7m��z���:�,n-�P���k�~��h�.ݧ��ѿ��w�c�'E\HFh��<�͞�[��W�\��$���-�I�Af�K^�Z�y��g�}����_����_������z^��J��O6�#�+�~��{���)�yQ��E*�&_����F教q{Wġi��xi����I#4��U��(�ˋ��ᔖ9�����n�U+2�є.�=l�m�u'ĝ���d��VR�0����Tnr��;+���c0���m!�(�*[#�(�������r�~�GK"&(�2]L�����B"�V|��
�L�Z�jۍ2�1dp��a�Z����ߴi���Տ>��57�Zkb�N8���H��[�za���p�%3��C�Z�Z }��Q����Ǧ��=��K_rY�?�����.�¾~�Io���m��ξ}3h�Y�-�>'L�i/���O@9
��}���c�0#�0B!�Zvs�hOL�MNl߹c��=�~��T�co� �q���&hMٮӜ r�07hX�0�N!�i�0Z
��&/�:I�F�!)�L?��,h9a����O�c9�Q��g0�٬���r Mz�Xc�guo�(e^oA���V"
��]ęZ�/��a:���I�Y&�,A�B��C#�:�Y�#qZ�f��DT�;���X,�͆��U_������R��i2=�1`%��-L�!��U��ۍ�vLZa��c���fZ��Oz���	�P�%P|�}�CR'���˽�e�ei���<�5ݴL��W�I�=��s��Q5��I�ZS�C��cа���s3�1B�h�wӴ��m�EN೥i����?h��b�mi5�$ւ�f�R'��nyqd~[S]z���C�̘�&L�~��D+jޘ���,kB��47P�&�e���M�.�H�~C�N�(X�ј]��y�L����&4�]kZF� S��%�n�5>v�OUC�����j/K�t���F���f~-���uM�-�F�P�c�?�*�BO�-�l(c-����t��³3Tr����C=�#�pdZ6a{v��X�&��
���fpyC��Y��N2"��͇l��6�&^��H0�>�2\�H���0u��nä�"����
h��EѯcS�ԙ{�g	G�۵�.S-	WL�)��ǈ�m=�TO�I ��!{b��P.xfY|��I,	�'E 0V1�&8c R9�8b(8�u�z�������?�q����Y��v�����$AL0�` �N��𛮹�%������� �Q����n�B�����B�c8vFs��
���	Q`�V"���֮��d붝k�8b��#��%��/��Y�!8��trrr0𧧧�V�#Q�{���������
քe��g�I�����=t�G�X���n�Z�vպմ��u4����%ܲn��c�?�;��������G���M�ZMo03��1
'?'=�䔵(��I���[~�U%���t�*Zy,gj�ZPI��Z�t�f�'���8���귝��aUs�h��۞b!Kc�^̌�ǆ�V/ּmG0	i6R�(��v`�`$�i�#�mfzB����.��w����7\xιaFBQ��{EDt~��0�o�տ�Z����7h��Ї>�я|B�ٹl����-��߶o߾be=����G��z����^��W�������V�E;t�X�csM�T��H�¶�(.[M�����>��������/~�.��7���_y�f 	��v���l�n��P�Lz��w.��A�c��p�k=�Q��,�~�I�tA�Ԣ��u�����;m�:
q��� ��J6��-1Z���"�|�X���!7|� ���3���։���Ĩ)��~���������������l�֊�[�1�p&8�d��}��g�ꅤ�<����o��|%��j"MMMu�Q���ƍ���qW�aÆ����8��h�Ͳ�O~�W����œ�+�8��O;��_��p����޽{w홑��~n^P;�p�"m�<�����?LO\wĪ.������;�z��{��A����l޼yf�a����(-8^�]��L�O�$���σ7|��*SW)!�+�]1��Ş�l�u����P8�����J��Q�	ғ8+�:WE���(]Ƹ�hf���\~���-*#+�����#���Ã����]������( ���l�s/6�N�9cE�+��!�<@���p �ڮӨÁx{���M�t�F��L�I�R%ա{�0��WGq���(�$�D+�J��`�+�y��"�4�?v�*j��[-�����'� �^R�h[���uC�Ԥiccc+W��]�j�*�g3��u�C@ӘZ�l6�	I����tMQ�r@�%�Պ�mqNN�Qm�0W�v�A��nx�+�?��^�g�a�}g���Ú5kd�^����2����+W�޷V�o�L�I˗�E���ܪd�i||<�a�&��0�)���B
G��d'��
i��)��5�z&b/�d�����P*��Y�Y.��-���cd������.�I10�t��x�pT���Ca�4����g�y�Y��߷o��9������oĴ�}�c���{0:x�W��pI�\�Z��*\��^��<W��Y� ���3_(��!����If>����߿���~�o�֫�u�^mii��{����/�ZwMȻ�o�Ν>����g]L�c�=~�5�������M���t�{z����u9!]y=r?�㨁H�:vM����X����K����<���_�B��.�eG�^�Q�0O�>�x���?���?���p3z>7d��(���w�M7m�r����=��,,��}N�t*�m�=u�^�������[H8(�&�ɚיg�Ixl�}�}��x.\UJ=Y��VJd�}����;�(������?�����9n��_N���f7 ����aE�B��.�Hq�$M�(�@�Dh��&�z�|,��o��o~���?��g=�W.� I�8�|���Q8�w����S���w�".^4�zMK��3�p%r5�3�QT6��߱"�6C(�[Ra+���y���ԓFWc7��U`-��f#��/���\s�s����_��(Ξ�����mo��'>�{��{_��P�%�,B%Gࠧ<�Y�Ku��c�Bh��#{�\���ӕӮ϶1�:h�� Y�+*(�+GdL���&����,!G��sx��*��4Fn`�-�I��,����i��''�h��^�Gkl��pu>�_��JU�)ey;1�T;�����Z:��6��do2A,F���{$���I۔)�xmi�HmӃ8tPwBq�^fɇ]5�@q�-j$$��W���G�#%�OQ�U�grh��e7��8Jp��x�rTU���5��r��m5BCݵ���~��}���3�<m���z����O[�Q��[Z�\�붙��}�t���l��z;���o�fL�)B��C��`�s�,[��H����ZX>���Xr9�Y�<�x����|��f�� ���{��v:��No�����`��-�TXeH��h���4�"�5*<��i���L<ΪM,�+���m|�LTR!*P���;\����ԫ�\���251��L�-|VyJ�f~[����~X�>c�T�B<�i���$�{��қ��3K�2����ĩ����>���q�ph�����]�;�:�|���I� 7*���� �~��73T?ɻ�E'D�[��"�-O �g4�e5�:q8��q��u�>N4���D�jADKT�f��-0&�E�L��t�*y�uK���^?��<Ǐ�(:J_��VM��e	�<��[�+�jq��X�����;t���[n�k�q+���P�E���,ѓH�w	��5����&UVw���M��j�a���jǝ��v�%�2�&m.(�ei+j�NXKZՓp����]t�
@��FA-O�O�׋�����ZҤ/��=7<�x���z;4I�4�7������n]e^��A�4��dr�`��
�V+u�5-cԭ-�$)���']�����H�.9i�Ǟ��l/u�4��v#�	M��̦k�qM� s�^k8uьJ�a����oky�����&i%�Bl/@�-$�d)�w�߆��hK�`݊���ͤ�[�Ҩ���%)-sd���,	� ����Nݫ`��dv��!��h~�ۜ���jO��X5e����'��t{��'�C�QhB���b�F�V�E��p�䠪���8�R�m"�V�28�(}��4��]�w	em<��K.�Ĩ��F�У�s��k׮�Q:/�Z�v��4�0���|�|�Kw8���+Ʒ�N�������;��l�9���?�|�O;��K^����%BŪQ���[�\�Z�zza��d���ꦎ��+�.i�n(���9��R�Q���h 훖N8�.n�V�[ܹka�}�ƍ��+֯_O��ҪuGE�^�<�ȏn�s߁�����oA�o��$�NC;r�����=�LO?�}ow>�����σ�m�A]�}��m[�|������e�b��S$=�L��'�8eEi�Ij� pҺ>�Y�]�i��e�����VZIjB_g���^y��.�袷����G�w��QB Rc���ݾw���,y)5�"u���n
�Ƅ���d)!���J��߈H�I�V��?���=�y_|饗E�*�2����?��G?L��/~I������}ӛ��jjd@�q��?��7��3���K^z9�.�����zZA�W�T�D���I&#Ս+5�I�;�+r+�R(1�z�:a�PYkrS�+1)�M��Ed2jm�+��8�\�\��Ƞ�F(�=�����e�}��_H|�{)����׿�٫�u�5�^��/�u0Y&��$��FQt+&-1�QBj1܆�y諩_���k=���|�iA�l_�I=Ӥ?�7�1��8��u�!�,�(�I�Rn!CѐB�hR��	0@.�S���q��-��(Z�̖�����P0S�"����A���L#����^P���&ZY^C|/����*�P�:���r���e�6�������[��DR��4�b	�.Z�`Xs���7���E�B�S���m �(rm7���U9�����?𐎕v�y~)0z���X�s�1v�1;;�wnH�����̾}���5��h�'�H�	J�e+W��;7#��}1	#�X�mONN���I�#ሣ�>���7L-)�JA�3X���{�������mۤ>�Ž{������q\��nrގa�_em"�EbΏ���rV�m�E`�[ծ,���1jy�rd�IͮC6����g�uu.]Y�((�R���鬤x�_¨RDT�!�O��n�2��Zui0�1��F�2�,,,��2W\�-�j��i��FP���D���ۛ�߽{7��N8a�1����{�����t���>��͛7�PöW�Z�?� �&��
�<3mVD�
����JV���4�����ҩͤ�J�{'����oIT[Oŷ&�D:P��<A)ےw�ZX�..--��j�,�i�Gn!W.�]Q��x?����gXQp�<W���x���RU�u>=T�I�=�s�TK��D^R2���3 �̤�	i2m���X�9�P��=q�d(�먝47�Ba2�����:���Ya��v��������:�9<��*Z�U|tF�(�c�MXmb熨�!�Y��J���B3�t�����Q`r�3-�$�N� U�Ӂ���\��Ҕ]5�H�d�4� NMLL8A��J�1�h˂]��Q��j�rc��<Ǟ�!Q�plz��?8���7l�H���-����
"�D�ٿo��P3H���۷�r��#�sLAonn��#������?�}��.���s�y��h������+�$���$�O�Q�.H�@?��TI�ʗ@`.4���q�
�&ⶭ�Q�f����>B�_|1���＇�kf�Ɂ��l�ޖ��V�0U2']���l9W7�p������uG�|��F���������}�ݗ&y��o��ǆR�i���l嶆^�'T`�I�;9
��Q�#��S�c�tkB��`� ax���?����s�}������6�f�i�h����������Θ�,�k�b�����v`��P�81s�1�i�o��/��ꫯ��L�ח���|��^�2��L	/g)����	9QY�L`(��8O�D]7��o�4�W5��%e��#~*)�(�Z9*k����Q��J�+��T�z!}uj5dy��$��� �fiB|�ޑ��Uڡx8JAo}�[Ij}���]�bRcd�(�+�����{������5k�d�vV(Ԑ	�l��X#6*�=TW?�����k�q�#���<�CD���` 9h�.8�iveF?J���a�~��EHc�"�#��i�)�A �VOͰ�e�*�i�uP�I�Ra �\c*���E� 	������E��(��W�X3z�dE!NU�=@d���("��U���.�^�]r�l��]��>��\�o�N)�=�����s�C"�G�m6��
b�'I������L'K�Rt� T�����2�C$���n7����!)C��c-j5�*,O~�Q����z�c��)%�#�u�E���|g�]wl��7l�p�Ev��@��v{ף[�߾�]�VMY�M,r=��es9�&�m��a۲O;��p�n�����y���/�h�-[����g�1��xtĕ!1fbJH�g�ċ��^B�3�f��ei�ض]tgf0�F����5�+R��hP-�u�ed�����E����-vf�B�f��
��twL�0�v�#���X)G7YS�DW�v.�'��/��eu�����!�噢F�ƽa���2Ą���h��뎄=l�E@H��pY���g�v��.�첾�^[�`��Dܒ��_Es"M���@�6�h��"��_��W�<�����j�]3�t�f��͛o������z��덷Hl˃�\s͎G%�O8묳���w�G�﮻�ZX�6V�����r<ݵQ�Y/uH	Gq�Y�4�D�B�z����v\p�O�}	�u��'}v����:�صH���ޮ��U�زe�u߹���1Hh~�4�"`�	Fk��5�dLK�46��$II�o3�ga�V�wþkd�p�E��н�K�.�+�z���(����Fw���]K3�ac8 ղ>�]T�������!HDȮ�HK��SK�Ȝ�h�]p�����wl�M�&�beK��D�,L�Z}�	ڕ�]4:cE�J!1S*!�t�F����!�̶W�{N�¾��vo��.�.$^0�@��!KOWh��'��\�ǰ�s��q��}|�yo��U8�3��F؇�;�����$6L�<������#�`#�ن�
���\��}nN��K6�{��d� *.�)�[q��E��屨wM����Ez���ih�L�������~�\�A7\�ܹ���Rg1:��qF����a�vH��dz�L*�-���y)
�v�)�@Qݫ]�Y�*�\_K�1|M,J`��]5�/���_^`�5�����ݤ�s�]Ԓ�m8���a�#���E���~�{��ދ_��s�=w��w�v�m>���G�{�3o�������s�<�8�^[�z]|`q��e�Y&���qƲi��4K������`�(/]!�X3k���!@S�=00�`���M�ܖ�l
6�0�v���	)�`�.�i�LǴɧaqڒ"�ްG�G�B�A<33?�g�ƛ~�h{��7a�^o0�������ԋ��z�	'��㡇����=S�L%����-��V8����>4�_�a(���Q|#K����DR).�Ջ{K�;���g^D��C�9���w��]���C&}�� ��4��k�f�-��ᨃV���I�N&mZ$�P!z<��9�,�w����ˏ(N�������/}��⤢�F�@�k!`��u
 �$�c~"�����U��J�@�6�SH��Xe���nq��{��ޣ���*b�m�a�0e��҆�(G�:�����9ªb�2��@3h H��n:6k1��CH�ڦ������\�寿�e� |@�z�O�ޅ������Cy����կ~1d�$͜Z�����*o�K����w��`��<hzqX|d��$�\@�l�5ӋP�N*�!.K���~$
�5�Τ*�)PG(z�ԅ��r �����ie�W�XsaM݂޲Ҫ$`I�j^�����;ՈV,�$īh@�!�����c$�X��De�J(pE��^��q�4�Y�I�>bsH���u�D������\g�({�2޹5֤II���v
�V���j6hIK%�@F�9��`:�>�a���	)��He�M�o�3}�����E�i�z�iΏ��ig]�zmٙ~�@I[1IXs�Z�b;����hUuA��Z�6�/Ex"�/GqI"�!��w�%:1�����"���~��l|b�M�K�fK�%)�]Z����*�*�Ar�*UQ>e�Iء�bJi����Ţ&ZņQ�I�H"�O�u�=0�5]X��/Ukh�J#��e:�$��llN�x����K�!�mh�.N:��O4�4�3%���4X\��zsE�+�
�e�q�q����ׯ���|��Ԟk���.kO���*N:�裎�я~�f�M�ڎ��j�P\��pbaA��M�B�f��M�%֪ޢ�`.���:� �Rbp�9R����X�����٣�:J��a�z1�蜕���d�Y� d�����
�8�!MD,D�⨆�k�9��(����gK��Ŭwz�_*�.��(�zY��DZ&]<���}�ã�8�,���*6#isU�K�G\��_���4/=���J+�3q1�qA,$�=t�6ׄ��r�����eJ!/y��5q�b�4�F���UM~�{�d<*b�Zk׮m�}x�Gw��5��A��0F��v��GEx�d���@�ֽt^�r�K��h���y�y�Wa-�R�>11�M£˅ 3�Z�Y����-���/�M#"��8�Ծ������|��Aq�ָ&A1#���Zy��"T5f��Xh����\���o�>��X�b1F��v��v�[o����ƍ�0:�c�,,D��ڵ��I��������C����cǎ��9����q�AG�l�L;���1-i!�MV�?�C��'��8[�÷ZHD���Rt	�2�����g�l�?�)`��Y�2Kb�VT���ŕ��D�k�x`�����0J}����M�}�G6j���s����d������ڲ;���%�G�j��:�U7���(���32"��4];��7	�����.�Ke&U4�{�~�M�Owu���~���hb�J<&s��ڶm[�O�B�����~�C���i���A˹��*R(7+��T8���6�}uVpQ��4n�{Uq}��)�2h�1���+EqP�eD+�L��u'�%]L��˪�g[E��&nJ��u��0!x��^�V�6�s-��m�
8d�$�̴M#��׼�5������Dš]����$��>����zfВ��,�d+8$c;F�8�$Q�yT��=�*�6-�,�;ښ��w\R���w�u�Y49�:�y�j����ƪ����3s3g�q�bw����z�7�z+��<V>��n���<��O�ӗ�֯ù*1��ƣ�F�*���>��7�Ͳ�_�����֑��,#�لU�~ͤգI�ѕ#���˻b�h�*t��pT��J2Jκ��T%���0��(ʲt- -�W�,�>*)*�%��3�Q�����w��ʥ�^��+����>��Jw��q��>�9���W>�A�lS�5k�ޙ3�8{qq�PCj¦3N���=�l&�F$3I�7�Z9�JH����*[:���$�����g�+��9�l}���=L4Z���.?<�3^�K��s�ٚ���]�4
I{���ds´G}ܪG�u9y=	����0����\��h�α�̏�*=�-ۍs��d�*1���$�b7?]�[:����t׮�e�x���	�}���i����]9��RK6����i�������u� �g�?�+�4q(4Srˈ�*0�qt�VDS`z�N�٦�h(���]�6~P��VaWk�:�M�H�\��a-�P�ɂ8b�0��Íf3C`�q%4ˁqw��TK��V�9f�sZm�`��<�i'��50��[�*����G�����wߛD�Z~���Xo)�w�����nz�k_;q�q������%��k�|ի^�����͍��쥥�����뮧�����[�l��j|��h�i7��:b�32� ��DUY�o��M�r�l�H������סV��L�g��v��q>�P�g��hY��k��߹���8�<z]7J	V�~����[B�`��� ���Ŷ����9�5��D��ƿ�1"��;��FN��aNV#��?6	�4�PY�2�:�|/k�L�	#_Q�IL,Ey�F*	mP�D��ВA��!5+w-�Q���j*w�{�N��t�ǆ��C?v̜f�)�u�Ʊ�|������<s�d���׍���v�?z�����TA0�4�S�׶k�Q?]bsD��#�բA]��{.��وJ�,J�{�mX6��<���8X�d	�_�C!ˤ]���"U��Ǖu#+��h����H����ð���׿��3�tVMҕ=�i$w����Hoaأ�5s`{�a/_�����t���RB�[��fk�֭~�X�qbL"	#)H$�#�B�q��	�2��K.k��̙`������tɏ�(n�����[Z�<��I'����\���6��z������~�x�94�3͟z������M�Zڝ$����;wlۻ��s�=��g�^��ܺ��]Ϝ+��N��ƤŢx*�;F-Z�ඩ!/ C䞏]���I҉���'���:������p�Y466�+c�T:�V���ܮp�sq��o�i�	R�nvH��=���No�Z�bb��I�[���c�=��[�:a�/�PS�	]�&W����|G<v4$��Ua�����[�K�qp�:O��*��0�W��]:�T�n:�^���R)�I,Q��ЕS�hJ:�H�Q��|I��Sl���⑪��L��tW�ZM�Z-�{�FȖt��/,4�-�MH<��XC�a�X��ή(�2=qlGc�ni�^�v�]6a˵VX��"������F5f�Q%˲e -K���2�C�c(<H\@�
/�gU�܂�Fa�l���Ep^��M
p�H�`�b$�����=7N��(��˯���pا�H/E�FN�����А���x����rQ���� �׽8CT>]�y4D!�<!�<�1ʨ�3����>~���nS+I�������&�� c�9��w��}���? _��@��u�}��|hI��<M��￟T�o~�?���Hq�D>8�G�f���=����>��XE��ַ^z�e��ַhm�G�v�LIq�����v�&�,VXٱ��
_e%堘L�OUMdY�bV��@�g�8��JT �[P�E+9w�;�z�9�Я�R�<���cӟ2UXt�G0�+^��o]uU�1F�Fp����ީ����x}�6�Z�"�?�ù�������ժ��Rkh�;�M�W��UaD�ݎ�Z�;VXͲgff�OGq�1돢1�C:s��ܹsv=��ÙS.DNsy�@�J
oP7�vy
WnZx���8�B��#|.���Z�b�2mB���!˥Ѡٺu���$FnX���$W�A�2��$n�LtD1�yX�+��c�Ε�T�\*}e�`9��Q3!D��G
���O=����N9�6G��#�/�|�x�ʱ���7�!�m��]��w���g�Gs�J:��{�����o[�9���}BC����C}%D�N#]��3�8��S��VӃ>HW^r�%��z*�"�k�U�V��?�|Z�`)���њ�Ĭ�|��V�'��Lq6{�įUj;��	s ~���h�/�YΘ8�����K�1[׾}���lq��8����U�H�.5�R�����
{��g\���*�C�x���@5фH*��C��6s`^�z�@�U���|O�KS�39�j ��^h�6����L�rցۆ��+�A/V�J���'�� ޕ��b���ۀ��3�-����E� Dj,I5���v9�G*t����D��99���!��]�<��_�6�li�F4��uQ-I�*���Yit`�hBS���b�L��
���"c<�*=I��	�`PD�S@b�N�5
��ך�3���,�x�����_��=�l�I���z���p�q����wu�Q�~e/{����젥�+޷@ JV�Ph�q���6�2<��#�t}��t���O�[۷op�V��ɧ�.3~�<�47
*B���N��U&��<� �d� �mz-ր�@'�ܖ�~r��iτ$���W؝Ǚ<#��"���Q�K%4�B��&"C�Hy7���s	n���C�l��e�g�F�k���rtL5?�����E��詃~$Q`h�a�)i@�NW�Ր��Ǟ�ؔ����&T2���h^��A@��?�X�m*UTI��:��Q�6�i-�>%`֞���X������!�G��8Rl��U���hHA�'D-��4=Ә�C����z�,��Vfs��Ve|�#9���^мL��U�5:OCFSH:Y���	��ق�.`��^S)���TAI)B,C�e���q��.h���mŢJ-�.@�TR�D���H I�N� ^;Z���E�ݭ`� �����Z������v����n��_�5�������<�k�F?�я����>�??��K.:���U�[���?x�W���31I��1��چ�'�~���/���G�k�ڵ=��x�2�(�3.y�V�'������ħ4e���ձ�v�	7�p͗����E�x4�@ax�2�\��\+�+�d����[�@W�F��gT�>��ѲaT��Uzt:Bl(���:K���
`���$Y�b�9���{'~��4J�z���W��O�? ����5�i�vJDz�{�|��k����[�����UH������G�����Wo�~�"g)'���|�yGr�L��L�b$rc��ކ�0[^�������=o�}$:'Ƨ��<���3���Vwƙ�vw�;رc�ٞ|��{s��у4�}`�]ݯ�W/����N$�q1˖��T~�}�p��X���Y��4S˸������r���5�XHSf�����z�LH+5�	�n5VM�h�㚆d-R}�DP����z�������Dg���Ǩ �U��(:��X�U��
�:t {��U�d�Й�J����*Q_�	y�Aϰ�����Y�$�5����Ө�rqm�`u��C��II�6��p��!���ze{���c�����.�U�Q&WL;�Gw�}��G׮]K[��N�ٻj�:����j�#��ZFGZ]�y����9��e�����o��N8aa߁��:뜋.�����L:�ńk��:c�	׳i�{n���6�u�4���a`�Mo��r3<&ǻK�`Q8Sr+�n�D� 5G����Ŝrk�~��L��ilh����3w��8����w��n�m���yM3�N�fE��U'Y+��4)ԷJB��`�oKA�x�|dq�tu��)���N�������I�V��|-��=�i뾑�Ӑ>�zk��)-��߸�)�1?��f���!�Ű�3j�zc�� #��z�YD��ҵag�����BF�Vk튕4ę�pu3UY���2�pk���f*��a@3�!Tl*���&�r̚e(��a��Hz�p`[�d��j�����TyñC�!h9���h�ô�g�5٨Mxu�@Q���H`��8G'Ƥ��L��<IF���L_$V�=/yƐ�Tƙ��~&8V�!�vб���bGG���7���w�ȓN�yŌ�<[x��K(��Ƒ?�,��ښ5����������R�|!{�E0�@������f�ǽ�5iZ���m��	�r�`�/�xh����J-`cv�-�!��	��K�1��y�M�����~��r󍄗v���ȶ�^��oΊ�][�.N�'4�{f��+��ZI]JK��g�m�u;������{��!���y����E�r�o��o����h&l��h����+T#�g�ȹ�3Ɛ:��4o���8
�칤wX���K�!m���O�ך�Zw�Hw��^�[���
-��i��x�F^��&�w�U�jӀfQ�U(t�=G���ٹ4�Q컆�U�VR�!�3���Q��s��[�=�i�t����|�.vL]�]�zW6���Tˤ�5�p��z,��:����\E ��\N�C\ZO에k�$�QjY� ���RL�ݱ�A@h��;�[�1+�NU�$M�I�G�nd�gP�2?;a+��hf�@u�iBԙ��Ro�]o*�k����mA�-d��!��:
�覄� l�Х�����$�3��X�Ƣ���&6�����d	*��D!%�]�0��@B�;U�/Q��U�U��4���&�_)�
V}��s�C�4p&�2a$�(���4���6<�*r=7��3Ж\��%`9�.b����4KC�S����fȁ��[����yt�����h��Z��\�?��/�:�y����$���x�)���fIt�y���'?��o~���_�g�uu���ӟ>�䓯��n���L5�����N���_���>������ �bC��T�JVE�=���f'?��N $rꦛn"��ꫯ~�+^a��@�'��E�sR2e�F	V8J"Gc%�R*���FV�,׊f����%g��V���`u�K_q9ńK�q���k�s6n�x�7�v��]���+�M�y���c�9��Ͼ��H\�y��g�g�.�����o��]�~���I�����!8�ºg^�h׮]�s��\�ߟ��J��>�3�������J2��[nI%-9E�X�~}�ZIZBNj��k���Y|�ƶ+D��:h�b?�����'��2�_�`��*�@�h�|���l��_ZZZ������^����Uҷ�j����Rk�/�)��ڵG,��GH�:݊''zO+Lz��+Ja�l#�`��]bQ^�j��sL@�!ZZ@-��m�ۚB����&�`�/9^�$B�������䱧�.N9dw��$4����cccԁ���ET��YM��x��r!����ҳ�>�>Ӡ�vۏ���	`������w�sĺ5�y�k�$��=������L�*L�I.y;،��0���r('t��7/���0Y��?#�ucYX6�|���=j��҂�b�AM�2��٨�y��c�dv&��y��Ƽ�u���
`2^L�Vh�EN#�:GSX.e2�5*�; ���?����]��zS�4��\Ժu��:缕+W^{�ջw�����:h��z=A�	:�:���X�E���f�nWCnX�� �����}�DD+�%�!�nbb�+�0Ҟ����	�u����-&�����e�ߧ�0C�A�Kc��J�v�e:b����ʻh�I�$�	��eŖ1���N���o^�ڡ)Z\��ę��Y��wny��Hl��c-�eǚ����΁�����(vtТ#����\��qq3,Sx#�{&>@q7%ǮE��V���e��X��)J��=��i"��1Mi}�qt+������ݻm۶�����/�Sb� � �V�ő��q���۷n���c��^���5��u˖-a0���KI��m��V���w�
VI#�dy�w6X�i��������0�U��kM5BL�7����1����Ņ%�P���Yfɢ��u��jr�H��+q���#ኔ�)�W5��g�M�%��{�}��;uߡ�n�Q(CШQ���Q1qH�9EM^��bp _�_��gEAA��"膆�n����\�����s�'��<���k��S���{�������f$���^������ل�.M���B�Y;��Qݼ|��%~�Ð�Q�pn$#څBp�k��v[�D��=�:|w�N�#�I�>�E����_Q"
 B�NG�<��6�F�J�m�$&���uI���iHk
�L��zq�s/1�O,��k�_��<�)��� PꜼ,PfG�.ю\���I!��D^PtS�y�Uv��k_�bG'$��OU�^�=DC(S��GI.U#�4JڥB)%�#kx�gi@�x2vO��n�Y�G~�P�����Cc����]�B�O�����
d-���+�r�������ƙH�Y�-=bXQ2���A@�	X�U������W��� k5������)*W��[1�Ph�����J����s��a�&o+��Z	\�(��0� �T�9�6��ѿ~��[O;w����El��ي���z�_��mS�Mc���0SX�d��B��ɡ|y�#��M��PJ�m'��<�|���t��.Ѹ\ɹa-���D��R&�He(7��Fꐬ�H�3#Ӝ�]��w���xە7�}��Qf�@L�A�ݯ��f�W�94����Y� �\��+>��?�i�j�wb�7�dˑ��~HǫӞ�_zd�4D��z�;:U�'���~u ���?R%���ݒ�PU���U�>L��lk>�|?K=�4(- 9���mƔ�>�<��t
�P��;�X��N���ʎ��6)M�+iqI�i� �y����'�'S����n"T5�R�F%;��*�8@�n�w��K
YBdlr�_�|��6|=նl͠�(;��$��q-�jj�FFmU��T��J/H��L��$����MZ�ҥ�8U]+� c���`ӓ�JIq*��<d��t����C7Jn���zFi����"$ (�,Vyה�n��Ġ�ሻ��m�־Y��*�������{�c��v�J(7hӑ5jG���9��$%�$�M�ݚ�7fKYRU���rl���;�80;=�eT��b��5?�U�Y-m؊Vc3c�B���K�!M�,�˒5���4/�.���mz�xR��F	H�)~�*��$�e���eZ�t��SuSsi�;QPq�@m���}�݉����f��YJ��"��n��*=�eZ:�T"@`	��p�lg/L-׈��D�c�JRʱbd
�� ҕ0�;S�fB3��4���'0&I��erf����HR���@&#�(�0�FWm9~ll�oߞ�F�5Z�~�Z- �������O2N�0֓�B߅0�\E-��K
�'�y�U���K#�V��%:υ��CO#��q�*����[BKm�\��)4d���§P��U��
�R_��0�tKM�:݋u3Ґ��>�N X�!��-@�Z:ki�q�`٤}�, Un�a
�Lw,.W����Kb�HO)�����+Q-E�Hy�6�J�%�TC�u���&�3C��:.U�=�r�`�]V��(U5��V�g�n���)��hO��UE����ryH*�`t�(&�-��'�1��fٮ�N�z�ޞ�����{Wn9���=�ƃzs��]�r��������4 �F�P��=;_��3�4r�033sp������,������ �Q�m��to��H�e�gM�
����;L�H�i��Jb2�j R� �I�z�h��b0��?Sځ�6_�M�Ἥ��6ͱ�iA��ѹ��]0�����DpLQ��&Ԥ�g�a�s��&�4������j��0.W+IȳWۈ\ r6IV�hW�Zu�<^�a3�J
�TK���6K]kp�/��0��SI9��8z�s�Ȟ��QM�˝:�.;n6� .�ʽU���H�~��W4��� ��tp*�
�ˌ�rP	�Qj�h���H�0=��܄�%���E�mF�� �-��2����4��[a� �LLZ+�#�m�J7�"co`r�4�ՙ*��H1�t��"���	�t�<�nS%{_�B��[���ta�E�C�}�C�u]>)f��ۣ�{�C*��`T-�'Dcy4t�"��x��Im�^�K	62դ)�2a;JwK�Ђ���1ث��"��q��f� 5�Wj��
-�Ym�5K�̔���R�\�{�m~J�����:g����1Ҋa�%&�_~9i�K_uya*yWB�>��,�&&&T�9묳����W-��4
Na�ڵss:#��2��-�M��Ep��P
&�����}���H�hK���3RcӦM�=ӯ�ZKf�I��CfL>��v��G�Q��3�ǺH`N�D^���2v"�4X�Y>g�u�y&1?��E�2]�_��C���_�����x���}aW�AG���;����?�}@�Q w!7��X�ϓ
b�+<?D?R�k��zc�ӑ��Y�X�N��  ��IDATn��N�� [��6	�� �/-����y��\�YqCY@C�ld�E]�1~���b��|��=�� %��������n?= �ڞ̼��D�'Y{N���8p`��D}Q��R�-[�-[�=fOr��N�����ʗ�[���u�Z�X�W����ƨ��!��e��/�n�.HW޻w/�) W-i61�|?��p�4��f ������ܵ5/Dپ�V�\�u�ֽ��4&��s��XOhqIS2S��v�]�Eo�i'��q��};wʵC���-~���_>4���=���~6��-/r���~��4�q�Nûnh��^����=HQ����}�~f�I�-$�H�iUh��=)Ty\F�6�t4m�����nwқ�L#ǅ��f������]�>�O�B/���� c�#q�$]�C�D������z���V͐de�;B$K�����ӈ�,;��X+y�[�;���"�R.]8Ah9E�k�Y���	[O4z7�tӓ������t�h�̲.��/x��ߺ���{b�C�]�uJv�F�NZ�p��9����?F��"Ő�&ѵ�d�)9�2&�+�N���mxtYz"?�����\�1O#l���r?��l�E���r��t�4!�V�:}�:��n�yzzzY����^ ��r@R��*�*��4��6=*�)��7��N��l9c�~�`U��T����B��-\��*Y* ghh+h�蘗�mY.!:��\�(��*�[�����%8��n<��d&+�q�4��D2�0܄p�xݾs���ENU-Ѭ5�k��)%�֍�6;��ɉbaNUMM4St�[o��j�ʕ4S�FS��}�����q���|ScLi[
��Iʝ�q�WyE�e�g�.2fn�f�N���2���:�S�u�P�}�)3��V��1��Q"�^�n� �M�՚��<���dy�k����ХSo��w�L��������X�`�[����]��5]�F1�OGb�{��=�?di�Q��;�!-�t+�z��[�D��ƜY�����8A|0����dn�f1�b#�x��e.�*�~8��F�
�N1�� �ܑHM�$��I�;�f��>8�d߾
m���ؖ�����ѥ6�vg�!�^����\CF�#���K���cv��:q�,�?��a��$��45T~�����ǉ�+#bd�����1��e8~���%���XY�&����\����F���1-<��,�#G�����ke��̱r�Be�o=�����G���ӛ������T(}�{�;���X$!����k���\G�D��,N�V48 ��O�ɟ�-r�I�����Y�)g[Eǫe9��yn��G�!y��.lU7E�`�0!�	��Xݒ?�h�E�����)�\�ne��,,Ѻ���B���(�E��Jrc��bjq�����K.��/��/���߾�/�C��}�]ݶ��-[�����	��f��G�&����yǾ�}�N�Q�.N�R�]�ua��C�c�n�֥�"�E��!Ƭ��M�@��[�.�7��&E�i������A�9���j�B��$Ū��|	�G�~��
$]�94��6Y3�\m��B	�Z���L��6��`?��KŹ���&�����d<�tv��23�{p%����ħ�4`lGEՇ��%2�mS���4�����٪N�_D=*�2� �W�2?�@�A#�B�|�\z��H�=f���O&�K��AE��Z�0�f���8x�	����l��H{E��/TX*a)q�PPr���6�u�m���#�6��9ϓ�5���&7��u�6�ر�!�K��FG�0m���I�L�(��Y�Zu-�¶�XX,eY�L��i�,����7x�v1z}�^�ˣ$J��L,S �Q@jK���Ͳ[Y�r�������k$c��R��O���j���}�Ry�Q�	E�C��LP���{$�7\��� �E3���V��H��8�HƋ0���/��tdfA����$q�OI�V[iA�Z[�<�qվX#K��P�D�V�4's=]�_( ���=�S��OX\6d�V������7�����dI'����%�MX��!��n�m9N��"���Q1��c�N/�2\��&eV�aG��b�/7Пj�d��?˅J3Nh������f=0\�У����6��ՊR5��=�����W��ԺfŨ�͸eHΩ��Nʒ�v�\0J;d�ym�)
̃k�q���y5���Gt�EmqBz�b���aj�"�2G�<(�fKFs�lj�s$%�9��Ԫ���:�h���0e���]��s�90�9�����<P��8c1p�RQ�N��E+[�]�N�z�^����EæJ�q_����( h�#n�k�i׼�Quŏ���"��J~L'Q�hmIH�݁j���B���P��v���O��ȁ�H@�]��Q}qN#9Z�"���1�]��vX����g��{������Tg�LroIR�G��a*&�N�^��M��3X��X.I��5�0~ɫ#�%����qӅ�*��47MI@���T�(]Ȼ%ރ.s��G}?o2ϕU�<�E�A�^���a�(�h�é��4`_%����"�݆�����*�F��FI hr�s3���dt�6c.jE\�,�Cz���?U�����	7RzQ9h�ʸ�-%�+U:LwK�Tf���ke]����>�:�N���9~F�dr��.��a�+ѳ䗕� �#��Y�0Bd|�5�S��H�@�B�_���%
��n�$��LOq�5��}���ԏ�=!\I��]�Zq��I�%(2~��|��K�/��5=~�}�c?DU���k.{�N:�$�WQ�����f;��>����Y�9V�Ք��]��ݶ
& �S�H����&lu�-����H�N��;�dU�ڡ��I�X4��u��dO�̑�)o��u�d��)�ho��#�6PIy�1�� �J���S(���C��F7@����?�я���*�/ϕW�6i�N����zba6�eF�-�|濓�.����~�;R�-�/�]�d��I�4=���d��&3��}waP�m�L3x/k�m^�z�ڱ1������ݻ�Uy	7Ulݺ��}|� �gS�A�[E\��s�h$�����l�0FFFN>�8���#'LR��޷o���N-U+��n��'?�ɏr�v�Ҋ+Ȅ�������N��� v�nn?����p�%�V!%���rj�'�[ʛ�U�&���d�4�-
X-ܜ?>~pJ�����tD�Mp��|��Z�F&�����1֠0Bg��N��ڵ�G9�|� �>��OM��o�x���w_��J�����8�8K��D4�텹G}�����a�o�ٳ�n��Z���ι>o��Y�ت�]ۉ#w���Tz���.;��[� �/Q�ȑ�lGV����5k>��O�_��`I��=�{���_��{�f�[�8�V�l������4��R���`���� =���L��,�^�B6ٻA�BǕ�i��yt3w���V��4�4A�>��8Ҙ���ñ��g�u�)��23�@c�_�W���|ŕg�y�2_#I�:�zk׮%[�F��ș�j��V��	�ݔ�3C�bט�FpoL�V����ё�@Wnzн��ҠJ�Q�؃��h"��U:�Τ��q��6������?O+�w_�;�*ɬY�f�y�w��wW
`�**���)XG��S��N0���2U�	Cd�hKB��-�ej�q&��S瓳.WR>9c]�==K��h|6yQ���N��5I՘J�kf-�ܑ��+U"
�������D+��� -˼����E�w��b�޽�ѯ�J�L�4�*����:�,Zk��@���a>@��#�qw�d��C���f����3���T]F3���03=axl��R��P$*��ڌ%89v����'hFh�x⩬�W҃W��tf��0��|�V��\�F5��Y�<�]|Y���(�~c����Z6l8~�:��굅��ɖ�;�F����J�0���+BU���h��!S�ӈG��%���M��^#�u�'kF���Ef � ���3���)�U2���0�M`����|�\P�8���+k��tŇJ��^��:���k��a��HC���U6��g�9 �%�G8ld4&Z4M=�%�>���L����Ey�L�3o��=#��2��̣�9��a�B~)�)H\k�[&*uQz GK�ru�3�۶!�SY5�c�( �u�0�����"b>I�9�4b���4L�a�˺��ih�f�-���0�/�;;Z�7���z�nxE�>�q#mG��l�x�׎�!x��_��o��Z������S�?{�;M�Zojł�R-d�^�=d��r�4
��!�"�.9Bwբ׉�-��( }�cR�ل��dvD* �n&mD~˧䅴M�"'��1ȣ<VOe���G~t��H�A��t�DOsW�`�3�G
V&��X\k��QDkI�d�K/}�߹�o?������R�J���m��(�u[q4��0�tZ�YD:%6�B�v�҇�ڝ�_�C6��^�hb�@��OՌы3%��#Q�1=&z����^� ��/Q3�q��*�F�+�,��٤Qˣaj��a��?L�tэێE�od�N?a� 
C�_h&,mlU���W��*�r��O�Mk��p
��V��}�����Z���k4�mR�Q��k�S,��D RpL�|�:�'����@��G�m[&p���H� #�r��7$���~�3,55�:��03=��m�!�Z��CLr@��^I��qa;�K�0������� ��/�,M-J��>/XbkC(�'�����5E��gb ����[O���^B�ѶG�a�4u�Պ����%v�0����+U�"���ܬkt0�w�L ��NJ�pGK�����Ȟ?���&� 0�i�76,
�0��F�,�FWս���)��(3�:*�wH$3�Q�hk��	f�*h&�Sڠ�K��h�J���z� ��X�;��\S�o�u|f���>�=4sd��0hX:�y���46�d!|-Hy�D�E�Ed#�	3���F݋ǧ��-4I6߷�00Ԩ5HyU�"I{�FU��h�Q�	��e�� ��tu�Xec"��c�q�5.�
A��H��C�s��@�W(�\�2�-����� Ee�/2��B�YD�,r�n�Uʃ�!�;�  ��:	j�q�Mr��#욠�-Z��EWQC�N��x���1&{�\E�z)\O(+�TF�9R�Iy�eC���4�5��E:6�R,s}\��I���6��R�(UC���\v�r1�P��J�Pk��f�u�J�Z5����gaf��Ȁ2�X��gP�H˧*($�67+�a�-��ĮF{;�9�z;E͠�9 ǌH���h%��>�A4Ԃ�0�B�B�
3�Gm�gfXd�;
􈥁?�|��N�]����|��A��Ut�r��65��"�IEC�떣&izS�m�[���� �W*A�C�4�l�EC��H��Z���C�4Ƶ�$�a�N1H|G��ʅ�>gd�2P� #�,V��E�@�N' ����$AeI赁$��B=�]���?,�>R�%�u�/E=���-*�yD�5����\�2�uA��_��	��Z�ځ��Q�&��-�4�c����b�" �!5���ȷlG��J<���LQ�f�Gd�����j{���@YV�RM��#��a*�11C�8H��J��3H�**4:���K��EɎ��*z�۽C-V��H ��z7�����]B�����Ҝ��#G���~H^%W$4 �2�0�+��J"��t8�L�?\2`�W�ĉa��y�@�ф�����r?Y|�j�k֝R�4c�dܒe@?gٴ�:�G�����|���Z�8H�Ȍ %����Fn����%�;��q����x�W_}u�0N=�ԛ~��6d]ڶ�v
�i�x��puZ��t�Nx���ɵ��T6�0K#Dq�Df�"��ƨY�q|���Q� ��k&ǜ��A.�M7?�P���]����L�C����,���|@"t�
~�[�z���򓟼�+hc�$��v�i7�|�;I��� �LS�L˗�!L���F��ID���R�U��c���\�d"k�2��H9���(�Dp-�G�j�h��5���ƞ���dE5�n����K*�^,�8;?5;00����bq����$����D��v M[�|��6�'럌�����9d�Ȱ[���ު"�a/,,�q����<� �@0Ͳ\ٽ��eK�Y]nd$�����M�U���x3G71�����/hr;]�|Y�q>e�4j�Z�Yz����7}��:���j�66���� a�B����F�X���� ��y��a�F�.���"l~6c~�/<�������_���;���|�ᇟxp��w�I��\p�."�?���۷ص묳�Z{�&�A�1h����wӿ���&���u�fI>�C����"z*	�c�e�U� �c1zR�X���[�nݰaCن���CѼ�GCCC����̜�?G�;M)3P%�$��:�.�1e�4PT,�yK� Y�[6�wۇ4?4�n)���<�#52a��l�o��ʰp��s8�۶m��{N?����oݱc���]�����}�Qgv��rP�eq�ȹ昭N��LK�C�?1T#�J���<�@�8ʕZ�M �)LXD�9=/����4Y`+W�,�J�4��a�h��O�֭#Y���K�^�v�y�G?��o}����nz]�Ć�;�a�A�?7FW�-�kRu{|`jLx,aH2��j�P�x+��tӦ��:هY,#K�~�ji��l>��i�9r�(!���Ifc�9T���իW��<���wN�p#��J`�B��x���(
$�<������i�Li&��ʤ3�"��1�65�3�
�F��lYA�<��d�E�,�2��4��Z��`�ː+�Hl��H�5[�i�@�*�F�VF�S��0��df�ZcF�!W�!]�q�F��N�5w?����'��ɸv���g�}��Bc׮]sR���B����	�����'�<�o�N��y�5�����U*S��6m��կ~5��Pk iQT��U�"�Jj�����"0��/���Y��i��۔���G�Mlt�"]0$��`��S&������ϲ���)���gF5̠��(�-ŴpH��5$�9�_ɐ��._��}���6�
ȴ�Voԋ��q�"jYU%���g�Yq :9:M��P���\!�Cz� �&��.��p���R�@���(���HV�!�(��m`� �@a#ӲQ���h��BQɘL�X��mr�F�6P�'���|i/K��*(��u7$�XŚJ�%�����n������VoZK6���&�B���[Ȓ���B��LƴF��'���+w�2�n-/�7�{�׾q���~���Å*��� 	��N:irj�����eڶe��*"�
��d2�������e}���l6\x�Oz�1�ڳg�q��C��Jvf9��S=sљ�6,��%�, �񏧸H^'ݛ
�e9�Q�Ћk�:>hѢ��jA�҄R��"�nFע8>m����?��mZ�Ip\�� ׮_�d��w������|��-7����k�F���+��~��1R����6 �2�W�_-��$� ^���t��K���I瘹PѲ�O���>0��d�蠪Dak10��h�<H��d�O��o2m�NE^{ŊQ���B4��=�n�Sӣ4J��-�N��J��E�G��g�''��/��(LK;�o�P.�[�R���	x`4E���t9N�8@p�	rȉ⼖����+��W�F��3��u{��^��
�U�� F)��u���|h	 �2ۅ�b����ەihd�9shrR͆Y�ꈸ#�㸱��v������}N�/�h/�v.[p�O!G��h��l�~�,a��o3?9� �Wr��Z�����˞عSյ�v|��?�ѽ���y��5E�������͆�j��wh��a (�L鞱�{�%&��b�C�A{c�y��R,��p��R�2�X[8��xj:ݪUcT[�ذv`l���	ñ�M�{�_�82q��4��,����l�O� H���a	�u�(��L#5)�8�ڕB?]�]oDAK��>�5�����d�$(<.;&yU��jZ��̉I�p�N�f��!L�"��⨝�^����XB�H.����cy����æ�-����[f������l�G4�j�Y4�aL��PT��T1��tdȐw, j:�jt�a�X����*����,�DBU�Cץ2����s��
�&�f�<�|�����]�*�S����'��:09�g߾GS�����I�1��=l���h�+����j?:�BvHC�1�J�������~7����u�h%kp�xe���w�;}�]+E��{���!�	����n�E��
%��DM�j(�x���+��r�v�%�����&E���)j��D�I02��Nb@A�S��:��Q�p%iL��nբ����� &e�\�Τ���ɠ���\�0��@Ԧ�y�t:����to3�|��%��S,�^�<[Ջ��P��Vo�NL)B#����	���H	�p�J� D�m��}�H�VY�d��@��L�4|��<X��$�pjn� �'��o�ȁ�i���U��S��7\5�?�`�1=9K���<p<"�K�
�䣐��_,���GKr6byY{^� Z��E���'^:f��9�8�KVRO�.�m��ٿ|���+AAbjh�S�O~�z��M	+���җ�t���u��ia9�j�F���F�GH3EY�%���kV,_�m�%���J�G�	BH�+.����_/�P���^��o~���c�u��WJE��/y���ߤ&�����r�%/K���S�	�靡P{��.r�8������<|���rK,����ދ�D.�~M��I�!�$�-c/Y
�g�v�5Sʓ?I
�PP��9���&*�#9�P (�DZ��;XѦpC�u�v���v����ێ%�;I�H���_��;\��<��Ͼ�v�رu�Vi����,���Gk�lAgs��o����{����?�x#�/�$��}�w�����2�g��<�I��L{��/~��^�o߾͛7{vͅ�����9g]�bŠ��Ŝ�z ��Q��t�!� �]LB�:���|jB�h{	�pxonM�RU��L���B�&N�%�5�\s�g������c�b��Mo��g?������s�)��%9��8z���G&ş�ɟ����"c��?}������5���z��z�7���F�;|,�HkIF1%��900033CbI6}m���?��$9���f��MLL���l��2D��&<EO��`�,�ʒ�	����0w��<"��^��z�?GFh��A����̪U�֭[�a�ZzM��R,4��qZ�n�D\�����E����I�LU��j6��'S�V�]�`� 6�k�@��[53�z�:99�tm�����w�_:��ar~�!"]�l�����m�X��G���'n��5p�����/y����W��[S/�J�sN:�x�˅g���F!n����l��2�w�y�5���=u�,B�� r���ӓ��¶Ts��\�Tɒ�y-�+��O?7�����8��۸q#0-�|rzz��{�K&&I<
-��m5M�t*�T�g)9�5���)�Ɛ�f�^�D(���T�Kx)z���~����uW�Rז��(�h́"aF���ٲ'�ֹg�}�������<�ٵk�ݏ�ݳg�`��e@�D��mL��%c��xt�ls� �� �l�"��\�6�s�L3�Xn$l4��J	i�z��#اY�޽��6��_o�,�{�tW۶m�{x��Г9>90�_p`���< K5�y���	(!+H�+|зhE�����I�MV!uf�����qd����x�l�$�2�n�a٥I'�͐ ����Y�4�l��c�R�"SC��&)���Vҏ���.`�8*���%��ڦ$������V�5�RVK�:����29�ȯj*3SE\/ݢۖx6�ѳ�`�6p]��$T�]K�HT��S0eh蕚�{�M�0�}'��I�8����q\CN�g�B������O<AW��lr��W5���+�*'r����|�|8�Iڎޡ����߿w�.��C����<� �;j�M�6բ�����nM��;QA�nݛ�'jO:�U�J�>|�!i��{!$�����ӈ�誫���w�������/�>�w���@e��v˖-���wN{�	R�e�7R[&�gʮ�����W\A7��b��X��[H"���w��_��VkU�F��� �z~zFe�oUQ/��R����v	T#�J�\r�M~C�rs�]v>Y|��4�v�k\�YY|����.�lީ%m�����4sHh	9H��L���~�SW��3n�����LF�9���_���J��{��~�3/{�kI�����D�_z��r��?8��S#�cU]I�y�u�6�����K/�!~
{�����k)�X�Ira�Z�CxLqt������_}ֳ��������_E�t�V�Xy�	[�L_�Ǘ���Vs���+.����O��;�����L ������]��O����+��*ITF�sÖ)|Z�\�*�����y��>�~��Ϧ��R��y�`��_r��j(�$��躝�Yu���By��Os���s/�G�Q�t爻�p�����HЧ	�'\�MBd�T��#h'�ڵ뮼�J���0)��Q��V�zի_s��vt��mw���3Ni�@0�?���k?���^%_+�RYN����NY�!�=��c)h�J`�J��g�Bim��"zM�
+���j\=�ZE����J�L!Ț��i�ޏs]�e�����=�it�%dF�>�[䎆~��A��0�~�c��o{�R*��E.�n����!CO۲1h74�ݼq�c;���5��L�DZlx��xM���0�ߧfe�06�[7?K��F����YaO��]�P�*��z��'�N<y���1�Z��T��D6�d]CD���!�7��I��+�=�K�Þm,�P���������#VT=�%��|]�2���
ϖ+O5$M���`��LѰ��E��i�V����_�;w�����G! �g^x���Q�����9����+W�DT_C�~��޳s���v�v�r��z���m�c��|��dy���԰٤����9���[�秦f'&y��MȊpٟ���e�g!tF9��.Mqh4�4:j*�_S�\�֣�Z�>3�|��䎇{�vˤ�v>�#��w=qB�@���sS���¶fk~�����`���F�=8X�@=�X�-SSCU��p=ڮ�NI��*�v�~Eh�B�rh��-r}�  [�n�X*ͷm�5Cϣ��� Ѣij6�5�>w�Bi�0��Y�u5m���خ�W*��v�3�8������֮]{ܚUd�k�qū.-��w�9������~M�dU��'���i��X��G!�������%��;��u`=W���c�#��k��t��u*2Ӷ�d��._688��SSS�8��3f��f�,W6�Y���.$Kn��2��w�~'YÖiH�y��Vq���$�Ar2��J�$��e�_$/��[ru�0�x�"�6x&��5�2/��4;�}�oʹfZkvN	�V�n�^U.���9��I�����郳���UJ�FcB	�v'G�gTu�K�JBwF#0=9��RU#�O8D�>X���U���i�!m�,Z�^�.Ҍ�1x�k4؜���I�tE�4uq��ܸ���>a@Tk\q����B�����,�j�P��L��V���d��k5&-��a�[M��ț_��[�<�Ja������}��ID�^!�B
ev�����[�n=��3i�'�/޵� -������j�a�;"�+��A�6����ۭ Dѱ-��E�cۣ��#��rJ�uV����N�b�̙ظTrt}��)g��7�C�K'�*կ̔2V*gYUl1��0���L��tG�Y��<j�!xa'Ax�w\x�E�n_t�E_��������s'�|2y����߿�&��K��$��>�KA0S�C������o����#����e��I�m=.�^8��6à���ᕯS4����뮣�/J"[s��ַ~��O�����Mǭ��⋃�E�G�������Bs�|��S�s�?��/��g<�DYKG��y���m��#Si����k��nH�)�f��s%���$���'����<G&������\��);�T]�E�V�* �D�Ț��3i��o���K_sݗ�Hn[�g>�s�{�[����?�Ť�h���I��3���;�{�{�{ꩧi��
eY����_�w�^�*����ް�/٢�e����1���k.�|۶m��O^~�対�
	Dd���g�������U�a�W����ۯ���<�9���K��h��7�@۪�h�$"�~�k_���j0���-Ĝ����K.�������?��7|w���({�u5�^��\r�+�.�?�W���˃ӲV�)R^G=�����0����vX
��#Wt�'�T	�4��XbdD��׹��>��Oτ�}������G>������w�9��?�r}E����x��i4:���Gփ����9|*�'Y'Iؐ�k��ޅ���$��<�i��ɒ���;a�J2��_��l�K�C:\�̴N�fv�%(d1��W����RT��$JfY�:zB4���λ�������������6ߙT����VȘC�4��'���K9Uz�pMl���28_��-�M:gvv�g��2�'&&h����V��T���}��Ԟ=t�S�����l\�9��w��8�f�Nڳ{7]�\�͛7kܗB�Y����1�'8��ơU��O��B.3$��炻te)�/L	u��:(���k8a��y��ќ��Y=]�~���'��������{Ow[#1��}'-0�	2<%0Gр��
�����(�B5����;��F,�������`xA��n]O2��t`H�;�1Hd	K�iZm�,Ќ���"$�ae��Q���!�����N8������4��~��3���'$|U�sk
�BH����{���b2:Z]68D�@޸,𖣍��M�d듍-;�d�!rΌ�D�d�"��>Ea���.6[��ϫ���d��P�}��$u���@�l�f�m�H���$��}||ooRK�b��,
e�L��������4��3��8�.��X
:=�H��?cW�Iǂ��k��%�;%x�A�����s߰���h�����'�X3*��|�O����෬�dע�1Y�t���n�c�}�J��d���a>��5xe������rI��uY� ގ��n-�fffd%H��X�\M�E��e���yR5�O<�D�N��Aҫ�K��j��"�6�����\Ȁ8� _��/);���f�#	��J�I~�.���OQv�b���8�C?W���yE'<�W\qi���_�p��%$�W�%R;/���;３����	Z���-&=OcD�������{����*��Y��5��t?�F/��z�[o���g>�>%3F�4�\s͛��v�x�����V\>R�7��k�J����r�w��^q�eO<��Z�B.��1��Y&5�^΁�s�C�#��dGx�R���ݵ���ssQ�S��H���c�K��I������e��
��3��m:� G��)���駟��w����o���J�<c.�ٽgϻ���ӟ�,2�!�j�Ӆ�U_��o���.�$7K���{���kAԲ#�z�b64�]���>�������N�}�h����t�7_��L��]�)4SD�׾��t��'���h�it�Yg}��� ן���ř�K�A��N- h��c��iŊ\�W��-���u��[����x�{�M_�EnY��� 4��G)9��D�e�4D�~���<�^�;�:���:I�a2~N;D�L0Z�1�elګ�63E"ק**�۲�c�����X��<)8�}����s�>�Q�M��[C�Z��g���L�vs�9�zG�a�Q��r��T�.f2%�F�:���^��$I�8�[����C��O�´X-;�L����MQE��T��r�g�2�}��UF,���^]'�Y�`%����'��'0�"�%tQ,�Qӊ<onf*��2Qߚ�F�n���u
�a�(qD[	.2u�&,�x������i"�R;x*K��N~�ǥ����u77�,��Ftdpp��Ȃ����0�;����_D�e�Y6
���H�J�'���-j�,{���j��aچ�%ӌ�X�7H��&��������I��W�Tcarzvrrv~fvb���زj]���}?�᷾�ػqr܆��s6Y<��#��ٳ'Z@�f+/��bWUo��֙�{�}|��;:�L|�GK���/����IOEJ��=�\��.j�� �8bC�fiF6����W���f%9{_��7��F�������t���'�|2Tԅv�(Z@mi7h�FV���O������E^KF�v4��aS����{�_=���n{�3�U�&�J#J�Z��Ґ�I������r�I���ҫ��!{�T�k���")�SC+(��)f�
��Z ^_��p����鋞󜓞~<  2񆗾����unvʱu��B�C�(tt�#����n8�|t4ZV�&����GyA@��́��sI^�\��9q�i4­Ч��v�,�9J���)�0K�R4��%S���Oֶ#Գ�����dD�y��'~�Њ�+N\�����<x���z��-��^��l"�C�&��$J��6��صQ��;��VK����dȆD�ɖ�ʏ<:Y���&OԸ� a����.��*�4I%�,i"Z�`�JQ%�-�$�k��
 pF��y��S	�ݜd�U䬗�X���"��jt��DDX �)C��/+Q�-P �:���)Ṗ+�����TA�E�.ѡ��_�G
A݄�Y��FL���ǟ�M7�X7��,��!k�u��F����2�]M�m�dLZ�ٰ�PQhJ�<>>��(�Q� T�,�ɧ��g����|̨��Ւ7� t����m��ʃZ�yӺ�ʏ?����&"IFb��Qo�y������v+Q4Z��&y���fZрt�������^��Q�O�k��kӸ��������^}�����Z�].��}�L�s"fIy�;�1>>~��O�Д^�� ��h"�KV��(�7n����i��$Z
�*�bQ�j�"���>w`r����N?=L�d��03Z9���ݵ}�����ԛ��m�]���qh��`�)�9�ߑ��a���	4���=n/?��7,���{DyuF���`6G����l/_��:?7��+ȼ�Ѧ�di�CH�)�ı-��j$#�|�#W]uՍ���i[O���?{�������������~�\Vr�.��E����?t�k;���uM��۟�Et�{�~�FX��e~�� _��-S7uˢ��v�Z��u�qW�eX��(�C�궈C4���(!��=��KH�����{���:�dLڪ`?��5���:���v(rT����?�я��g!��H��j˕��)�5�U�2���s�L�+�$98R^�{���1�`RQQb
�dqX�E�r���>��w~����� X�~;
�������˛-�d��i�� ���g�Z�K�ɝ)�S�\�ߠ�´�_X;ϯ�q��ӛN�3���H0٩�s"�����HM���0�0L\G%L��Y�!\a�i��הQ@�Ւ�p�0k����jD5�e�LI�&�%4Mb7�[C*zY��&]�ad���y-���u��-9�����uF���S<.��O���I5�8i4P�8d�n�꾴Vߵk����׫�h)K�:�B��MQ*�$-Ld�F�q��X�߿l�2������>�`w�tM��<��@������R��Of�������3O?c�ʕt5��[n�ea�6`!f������U#�]w�W�#�27�q�J�Q}y�L�SM�����|���J��W�d�Sʒih�3��ϼ��3��/dFuժUQ�H�)CRt��G��~�M�6����'��>��8`�͵K�B�a�F��Υ'~QDΛL&���|'���(5c���6�D��H4F�+l�٤��ÄF�.888X�&pdb�&��ܣj`]��*��*^��DХ�n���+Vl�B�p�C�oذ��]�}�Q�H#�V�Wz�!��.)<����֮TRۭ���pȞEz���>n�������`vv���l�P�.�0�.�����σ ���[�._���������)�2�6\��9��{챐�0h^v�OCQ����D��Vf��&���$K���u�ꧮ?�Z�U_G�5z��&=��#'0i��A.�4lG���G�f�^�x 2��aQ���+�\u^#�Wq���(�,C���G�Hժ�u�I}uceD2�1�g�]V�n)��h��<� �	�&ur�+c�U��Q߁��t@c��N�h���U�&�λ���hf���:��G�\�w��1<<\dtP�$$9rrc�Y�ӕ&4�3��pY�Z(XP�^T,ڴ ��7tS���@����\y��*�h�}�Ne.R�D��[��y-�,�; �L�޶m�����L ��MҀ9�C�Vh)g=�Y����T	5��#O�}�К���V� I��jJ�!�wJ��s�N��s��\$�L�Ѐ�"�,-��M�y��j���~���t�Zc{�i�$�n�����ӟ�.��l�X\ǍB�7J�)��r��.����#3]�7�-)aq�I�u8�S+L琛���`ܺ
!�=;� q��'a���N��Ku(/(�/i'1u�cΗ����{>Y�]t�_��_�ڵ��?󏧟~*�*!�����_�5Y��|���y睬��e3��������9@�kV�%���X���1��$����N\2l��-�_lh�����)B���Z"1-8]�Ⱥ [r��i�dQF�;�m��v�st��Bs3�jj"?SlK�Ȥ�B������L�4���H�R�I���D�^n�?�@ȍG�<n����ti$�,���6�!*�W����	4
~��.�V�aX��H6��R�Za�;��K�'�NJ��jc���hU�a����zn"�U�h�}-a+E"���R�̳���|8r.�A�)��$�@�n�A��k����7ԗ�Z��&�q@�<e��EY��E!'X����.���"�ܡk��4����ʕJ1TBc1����L�L{�c1lJ"����D��R��NͲ�(�H�\4��h9I̬	��	rJ�
�J�kr���[OKI�"���$�~�˕��&��ܿ��>Kk�M�j�wϽ$�nvO��n�X�\v�Qs�%�Dl BG� U:��I-+W��̐��:�gnZ�z��8���;�߿6q��Y)6�9��o��o�ET��%[��6�kNM��=�ɊR���w�|���i3&Q��7�q���]���{�yxۿ�Y�r����\�nt4����\�j��ā���г0ʂ��d?L�K���1Q{n�%�w�ǳ�ChSЌA�[�m�>��Y�@_�Yg�E�����cc�4"���7,)˰˚���(x|�.XIHV��X����Q�T��w	�T�T�bXŪ����]V-�V��E���ˋI��M/Z��c��d�'��~h9IGOM��!6T-�J��r��.j�H��J�$̶*Nan��v��'v<�p������ߟ[�� �[W�fI���dz��Đ�O�kX��75}�R���Z���=�22d���3>>1:4H^��P4S3����J(Rf
i�0\�niI�H��(N-��7f����_�k�Gj^x�M���X;�z��g���oٍ_�:�d����h��u~����"�ЋG�]׺�?�J^V@�Hy��%�!�����U��S�sb �		iqz<����H>�T^� ��B'��?�Y
fb�V�,cht�f��h�D5�-���6F�o&�V�%#�TTm��i'��8h�����!�NF&8Y�N��Gaƅ�*��'i�����M�L�Tr�$t$Z�P�[�g�`��R�4�����c�ڴ%r5#'+��F�y��Lٌ�-� �b?���%X�_V��w��"�p:��fh���}�$�iNa|�]n1�Qf9�8/��$m'��LM�Luzr����W����LE�K3]K)E�h�h�H����IT���(�8��h�S�O_�'��T��rx�G�
"�)A��w�� �݆H��aY�ض%�Q���A@�H2�,���-�(�������r�_���Tx*�@�j�Q��l��nX6m԰a�� i3uG��%5W�"]u����fLʧP*�?������UWC⤓O���`�C�3�Φ����w�EF9�s��H�0�n��s��Q��k�0�`�"�p3�t����!L�<��5�u�/�� {C�X����d����[������=W�/D$1�[g>�Yo˛>�я��K��n���{�+^}Y�3��'���o�� -"�f͂Iޗf�$���B7
q̸j�������k�h�`�-�.ح� W@XN�GD�>m�v�$B����N�m�$[�H2�R��i�&#��;�y�� 7�Ű�R�E7��b#�8�If@�D��@ ��i���Q��p�L��If*�F�V���n�iI��^K�/��X�S�s�_i�i+�����J��ML��C�����E�|$^��{�G�����2a���\�,�+v\�6��R��i����y�R��,�U�krHC6�o~����C�ge�Գ�A�ό��g�Vo��7m�l��E�pIW�L�����bŊ'''��,	���<$-���;�m�HZ��L�x^jY6�:��F���´�D�#i�b����d�˟Q�ܿț�"I<*���G	b�I['����KƘ(w[t
�.:��9dS�g��c�=�O��d����� F#TZ�]��͛��׬����#���7~�V�֛dg8��#b�K\q�4��F��w�u'��dT�US�8�g�_��-[��{��֭C���ȹ瞻�o����������K�c!�:�%�B���4Ila��7���,
�/[(s�6�֥d9�W����n8��={F���[����RV�ZE�~�����+��GF������i�C���D����Ł�d	ڸ�pS���z-��6���|�j�A�|t�-.ւ 2:}�5Ew2;S,Ә��4b�*���pc��֖tUX�511��ЭҘ���C������Ή�333��#�u��O�9��l��9Z\\ܽ{7]Ƕ�f@/FF�����V*tf���3�x��Z��<Ovsal��p�]+&*Z鮁���$c��������O=���'5[t�~��������:6��9�V�֭'�7E{	X'4��g�*��,��n����2W��{���:R�U�峯tkY�E*o-�A�,I
�-`�ꨉ�g�_�!��R�ѥhgD�X�P������W=�L���>����`8�N�n���#���]"��s��sYS�?�\7h0���r��� @��M��I_&�HNhw�9�lg�����|�v .@��}��48�Ez�9h0�<�H�(|0�![]vp�Lbi2]��s$��邛.k��#��Va�S�u��&�ꍸu�����C=DʇF���68���g/����:Z����%����>'B(vz�W]�j�x#4Ĝ3��}��Wl[j��V���\.�������h���pe��5FT�;����@ш�p�	t���r�m��X�e?�mۆ���Pfx˴�"x�������]ՙ��g���e�rP*�$$� � r��$�n6�t����l�a\�]��A���t� ��aS��i�B�hHI�<�e����̻׷�9��rP�����I��p��^{����[�靣�e��>̒�U��s��D$��V��ԥ%В8&ì�ȝ>C-�|,�߼|���yϯ��7?@=?��9�"m��Y���n���8�����#�t0�Ї>t�-�Ъ����?N��@\=�\%R^�y��*D�˦c���k?�X�3Vs�p���Qk�&U	���q-��I�v�2C�r<'�tl�6`U�`Ij��i�BH0�
:�sPt����¾�GFy���v�[(j&��I2�7qu6V^Z����qQI���`�d���Uj-�v��Yg�0vC�1�s��K@������$J���a��R��<9;��h��4�W$���L˥��N�ϻ�'��FG�,��4��th���h֛4?I�j��$�s��lh�*m򬜪��*��΂�8@Eue��V�.�«�0�Z�ݕ�.�]��Խ��ױ`�U'D��C첎�qt���+(���L*�XyBJ���0�6�����Ldgf���`�#�"%��E4D�V5_�޽d�m(����0�*�Ģ"a��Y�ȴԠD��<?�b�[@s�i�آ�H�zc���C8��'�R�7y:lʖ5�h���VVa��Ud9�rV��$��h�Q4�BD�hY��d�CGN���7�2�v����f�Y���f���n1ӶW��U��.w?���#G� �����c~=�u{��Q XY��ڑ� H�V����X�y(9}饳��E�YX�,;��<�3�X�m�> ө�I���0��E�}���i3���t�ʗ�z��\�k�L�6{;L"�"ฤ�D����ۿ󝋂.T�D�S2G��_8p����k�PG�KBӝ��N߱9�N!��4Ԉ������\��u`��B!^��O-7���dr;2:$��w�f��g�%��ju�{�T��O<�x��/��s�u�%��N�?u�������Au0X�emR����ڣ��������neVWHs����ml��aw�uQ	�4�2�F���}L�:�?�	A�F=$��f{�X�0�5�UEo��f��Ω�X�R6<�)*���jgqo���.A�1��cbff���A�h�����j�C,\trc�3;w�\[�$���Y�\���J� 
-��u�;���Q�u�Uuf�G��c�bd$c���Ed��ɗ�T���{����λ&cJt.�[s[-������� q�ܙ���}/ZK�򬑶�'�; �[���Uo6G�8�϶��Hǲs�aMk`:�HVC(}�+���8>k�`�|J�PA�0DPDb��웂ׂn(���$��9�]gm���	�xf���=���Zg̫5���߰}ǥ^��?N�i7���$���eԯ{�8@B�Ss�z��� |��N l���i\�$Z��Q���5C56_<$�1Ғ�dlb<Fvm8=3e�~-�����4?�喤��K�]P]p��
���)���#�
ia���k������_�ڴx.큽a/�#�ϺC'dR�Dy(7�R�h9O\d$sF�vw_rŽw�W�1@��D���F{z��<>�j�_t����Xm��Xm�,IM?M�Nk�Ż�Z��@�B�6�A������M� 5�������������_��X�G�qק�6S9O����xB�#i�ҙe��h(H]�����"�<-�� 
�fQ�3L(��'QRe���e�����0?	-��[4?����-oyKtۭ� �q̼Ǿ��m7}�#�E#�ɉM��tX��Bx�8IYi4M������ �unx����ڏ?�:Kc�L՜�\�X��{��":"u�N�&�?���b�D�������d����5��0J:P�<�4��d� ��%\�\Ъ�I���\��N��X�Ί�]��aR���5I8冒�-�1�>W����j�\w�$���JZ �,,֖T�:��%Kh�Kx�e�-q��fB�7L��ۧI��D�%Y�@X ��l-f}���f.p��EY(��ە��[o��Mozӫ_�j���ػ��~���������ԍ����2���Ғ�H��_R�髫���F�؁C;v�X]�}��K�=�H���Yk�I�}ѵ�\r�%<�}I�!]�YV��\;e�����K1�g�f� :��Y�5U38�y�Ϲ�]��.sQ��b@
�d�(?O�ݦ�(����`�g8����"`	���n�����ހsBP�uy~�Cʦ~#���'C�V����?t�����F4��<�O}�StBx#k��7�l���￿�D����:�@���z�|��_]Mx�*_�03��Jf����e��J_G�a������_)��m�q�Z�D����c��9~�[n��CVO,"#?���=u�$�a:8����<x��0��	�(��g�8��}{ ?{��y�;�I����?���*����۝�}�{�$�K���n�h�56No^uʻ�������_y�$���i����^��_��-td�M�&Tá����w|�t�+���k�i5�w�q�7��_�W�~�{�=����o�:�_d%y$��$��'Or��-;"���mۆ�k���C��� "�Ϙ�ڋ�]���a��S�A���� U�k�s2��+��h��}���?����v��R:N�O矘@�*W疯R2����R���B��7��W瘞r�ҳ�����Pc�Z�N:����������l��x�2Db����.�VK�I���)�59h�����0J�D����8��F�n̈́	�{"S��Τ%S�9��Ei�$^*�T&����9��(ԃ��c����L�v׍Sü��Ƒp2y��A�[$�$������u8e��K�911q���믿~ۮ���*wUp䓫��	_|��aBk� �Ʊc'����w~~9n��{��AW�m��4�h�Wp�$C��	w@]?���k=�V���i�<��P흙q-�욍�;�����=*B��c'�^�`ĵuׄ;��?}�[�O���[�3D�����gЋ`�hM~�G^��/��ƌ}/F������_��_�~d4�i�c@�,����׾�����H�Ųi�Ypgk⥔���K�h#Iz�j���&UŪ�jQU�2T~.���ݏ�e�5l�������+o��o~ӛ������'?�˿���j�6�{~m04�t�;�����G�Z���}�{ߗ��Rh)bO�2ل+��(@��T�A?{�A~���k+ �ޭ��j�̑��#se�<I� �@e^���0��[mq���D��M:M6x�R����i���z�����:~Xo����������b�~�l{3mX��"��6w�s�Y0F
T1��3�r8���xU�Z��G�ֈ~�p�������x�8���Ta*S�ف�#���VY��T�$�%1'��1[��݀T�سX;ڵ����|�s�Cژ�E�Sm%��jCC"9���^r�}�v]z��_O��iX{��C����<m�>�RԥW^M�����N��[^^u�Ed+v�n�>��J7:zb��s�^z����6������A��� ������A�9�;ﾻ�k�-���}7��1uQ{D�iݫ��c��D��U��XB�N�&�u��;k��ߖ2�1�P3K)�=c�����(��f����m��ZWs�̆sy��� �n^�L��!�����l�N:��FƩ��J��Ɲ��9�[ێ��X����@H�xւh:��<R����a?�#��5ި��C����G�g*}n�V	�?���y��{�^]�
F���g3�mWg���,��%Z�f��p��7e�R��B$~��hl]Ne�,���{�|A���(�4VF�M<�D�׺�mm�j3��	z�4B��F�i���0�k�e��$Ka.vP��'	˘� s���~I�M��ݓ��cV��7�ֻr�'��.�>�u7������f{�9u,K���R��>�����}�֭�	�[��бC�������'��C>���}�Vp��`G��Ϸռo>z�Zo�hG:ӌ��=�.���K��}�_Zx�u/n��~훷6�����A�4�c�Vo�+��P1�Y����,�e�&m��8�|�ޙk�I� k���ԕ��L�TL2�6��&a���I-�5VS��Sk��v��~`ֆmR�,�x{�mgn������ ��\�\�0ZI[���~M�2�A�B��c�ez4ͦ���x��Hb�0�d"��6�jj���^�1<D��c���e�>c]����&`�wZU:��A0t������ӲI��ɐ�$��9�Id�^f�������`.�\ ��]�wK[:1\]��aa9��.�-!�M�����u�*lo:wȰ��q�03�τ��D$"s�Jqڥ�ǫF�h�i¼5�i�4���aMi��3��^m�S�Ӟ$dtjy8�t~��Ė���������N�z�����K�����4|�uWz��زm��֭��>1�6����N g$�njכ��[�\ߵ�9�T��9���y��B�ۻh�ΗOM!�u�ܟ�v�7�I;�Ӣ�uw<EF�k�ya�
�`%�D�0Xa )��4)�CZu�Zl�		C��C�*�UV�r�<^E���Q�֒���oĥXړP60��ʛ��+�c�������u�4d̥�$�dP�3���>����	��������std�`mH}����˧К�r��$Khr\�N�_'���o����կ���������D�Ciq䱞��׾t�7��7O���$�3��X?JS��^���_�z{��,��\ �����!�5b�bGV(�>��2���l��+�%���Y�m��I}�j�.mK�sd���)���p�bͦ1MhIi��t.�ӟ��g/���w��M��ܗ���7 �Βmpkf�����7��֩�u�}�y�k���_�峟�ś~���惚:�9���;l��9̂!!��>��g����O3��{�u���ֈi<�[�l�1O����ת�詄��صjԜP��[a����:.b�B�֍:��Ǐ'�����ݗ��5�	�]��致�/�����޾�~�!!���]M�r'H�����뮻�o�颋.z��^{��ǗQsu�<�޽�#V�?�>N�$ݾ�j�����n^$,|t݉F���a&��18��U�y�#�p�$��5�&Jx�ti�A(偷���`�q���k�Z�Z���Fs������PK��`j#�%;�}+;�Uc�*�b�,�t�`��G�Cl�T����
� "�i\�-�4�Q�Ņ?��ѳ?{φu�|[�0񧣯�"R��u�{�|eqYRQt��}��o߾������;��|���?��yf��!=wii�[������D>A49l�z���	Xm9������b�8�rnH2I%`rr�o��ş���y��^G���J������T2�����$��Ft�2+G�|���b��e��2#o˴�RK�$�Q���^ojf�7U�YQ���h�P83G���+�Wr�j*��M�y��$�"<&G��l�MR���&R�Īl�������;wB �:x����j����VG�rU�
���(m:MC�6dYu����	3R��f��K򤭪��iZY��~��6�`u��K
B��9���5]a&�� ٞ�����^��j���Qk@/b�'u�~E�������}�UW]Uo�WVV\�UL�[���!��Hڧg�/..���;I�i=�g��Ft:�y��s����Ն~E�6�c���ٙ�[�B���[�W�y�`�i���e�����M?�&cGr�^�_��_��?�?����˟���	�3�1��w4� �N��H�b�~0�Z��2�S@�D:���z׻��O������_��׿�e/�\�H�Rt$����O��o��$ν蚫h�����M�>RKU:_���,'�;2l
�<:U
�<ϙ�4_!yJ]H�yIh��%y�8���$o�+�a�yɐ�*�L�#����A�[~��R�z��Sᦆ��Խ	��ӟ��+_�s�\����:3��e ��������@��_���_����7������������Q����a��hȃ`�h�"���Fs�y�?y�k��=}��q���s_��!�kI}(ؠ�ʗKX�m��R�|ױ��4���`@&����\��x��Xg*�CK{��q+���ki���~�'���C��\R�5�Y�Bw��c�]Z����a�-w�څ���[�n۹uv���v���,7�lw�y7���N,0�t���jpjĽ�Ғ�k��s|���[���4"�:>@��5�mG�H�Ճ#yB���_��qXu$.fE�XB����^h��F;���)��A�]�6K�����WdWv#��0�xal��8�'�d�����K�X�`uG�Dgq��88s.f�	��_:��(�bj:��Qg3�T�ذ�U�4�P9��M�&i�Oq1Q��9��s��i���m�r����Nb7KÁ�z>�y�r�X�A��_wi�39���n�7\������^��mO̐9ќ8\�_#U\[��;/�1u�%�������(A9)¥��_]�`��y��z���8�y�c�=�曖�nt���՜С9���S��ݻ�^qɥ�p&Z�J�&�V/��a�� ���M&^Zd� �V��Vڌ�=\�E��m��� ��4ܒ�?77gI̊�%́�Υ1_ �Fr��mh���^a�Hj҂�,F`<�	JZ�i |zʒ8f3(%�s�&�*ܖA�3�dF����^���\���`-͑�PO��T�N�	����%%.�ʚ�@�\�VZ`�f�0%�@VP�".j�1yX��,묢ޙ<��a!��(�]�r۬��R��QPl$FA�gb�,�v/
(6:�Z��~�p�u��)}V�顖����[�>���W��^�ʗ��ؿ��je���n�I�߽{�����j����>r�T�;�(�D!���8<w�]<����\s��+^КY<5�To0�L�n�Q����ɸ��qח~`_w���z3�tj�������s����/�NY��i��W-�8�D��y\��}�+�W���+�����*�.��a�gϞ���0I�.%wٮC�䂾?�)*zhv��H�l���@�����ԧ>��W������>��Ϻn>%>���ٟ���?}3�<��F���n��G�ˇ?����G�&��+_��'����oض}��[��Z�cFj��BN#Н��@��cK��氽�(a��V.)���O$�
�L��%�U	�6�-1fy�=�!���\q��c!��&�X��X.-?)�u�n��x�_|��7��'����q�۟�짿�����7�����(^�����o��/���{�o|�󟧳� >�!ݷ݉� a<�����ԯ{� �U���S����w�P��u���v����Q,�Sl��H�R=���rŴT^��^Ӣ���S��X\#��ѣ��~�ۿ���LO��ʲO�<y�����y:�;H��֢8_\<"Hȓ����Ys�;��O|�v�v���W�jǶ�`�����>�Zw�uׁ�H�&�ִt'W0���W<�J����<����<����P�ז�����ի��.X�͸R\���6� kI��T1��%���)���s>=�%��eVt�},���x'�u E���������~�g�`-��2�^�,�Ҳ�.ʣUG��YZy9�U�k�b"�ODB����l�rN��[0T_���M�{>`T9JW���s�{��23�xo�=��?��?���oz�[��vZ��
Ӧ�� �qB�˃�Ν;���e/�蜤q� i{|��J\��dHG�_��f7]�A4H8o���-�v�����m���<j�]�I�����R�j���؏����gu�K����H^O��[������h���j��B�K|��*Vt����h�M��
d(�ZVw�� ���H�e���R	|�Z����K��C�iQ��M3�L���4"�Fp�99��z��(L'Dy��]\��
�p>I�,�O O�b��ȳ�hf5�d��>e��q:j�$Y,2C�X��5��^�Ih�^%_q�֭`�N7��6d���"{��P��w����~wl�u��
Q�8b�����k�˴��������H@k�;�$�£�.����M?�轷�r˫_��_��_�_������\�>t��]߹�������y�����yţ��ߍ��S%�4E2	M�뮻�_�������C=Dۓ���Vb�ㅰ��������%;&���pɣl[9��e�'��Ͳ�d�b��%/��ۮ����}�k4.t#�R��e��𶷽M0��>���}�s�����'��O�����3���g[#����d����z(|���C����E�9lU0�$q��Vff��r6��beH�����o%��$6$I�Y0R( u;/����v|)�T�=�������@������K_��,N8�{��{�?I (�1���>��/���p�-_��o��WhM���6� �[(��$��F��U�tm��a��x�ML�dm�2���c�~�n��.٭c�lN`��Y8`�E�5��p��)��)�޵��������ݱ�1�e�C	#A�O�!]������Yfܐ����:KM��z�-b���J;_�����h�;~�x8���u�E��>p�-�5��a�5�-�v��ς܉BRg�*3J�p$��$8�_p��VҔ���2�����`�0(eʳ�d�5�{��(;ZȠ�g�wּ��a��L�˪N�\1�#m��� &�ء��]"_�W��=�p!
� ��U�#��gI�m�ƃ��X)���� �A�<��	�t�J	VV��AX�s`� ZJ�(	{OZ*w@YJ_��\��,�y��"EYt��b�CS�xz������n�ǜRg|��)��S��ԩZ���:,�?�轷~��'������0ǃd�ĉ�j�Wv�Q�y��2j��z�m$�4�8�0�N����Y1��'��	��<�����ۣcs��@/��r�=�=p��������q����!�u���p~��3�V�tDi�������;;f�R�nD����T�u.l�cdDA�����^!��O^bz� �\������9Hx���[�ܶ�����,��m�*����(j�D���"x����/���	DIͽ��9�T8��G+���a3�s|oiiɰ�H��2��>�u"i4��C������'��NqIMF�%��Űt�J*�JDQ�~k;"�ea>Ѵ]<8Ix&����bRfL�ҭ�^�(h��gY}�d+Kˉ2���ۓ4zk��`0��ૡ�'&&<�k��آg��tow~��{�k�C�ٳ�U�z��C;v���C�>��G�Ӫ��S[Y��D�Gcsi{�6���S�=��8N���}�T����]�v��Q�^����{����p�=�.Ԓ�ʴ�9���H��6�*�E,���h��맕H�����l):�l��4��������o��_��8B��*���?�{����z;�(��ǳ�q����m2�8��Q�(����8!h��+Ml��k�}Q�����?L��:�%�׾��_��WE��W+�]��Л���[n�;:7��/�������c�A��^�����4)i�2�r�2�X�t��M��z��[�<�H�a�,�J�����UH\^beȊ�H�+j~H���,l�1s�Kv�K+���0g ��	Ou�%X�,v�����?�����o������۵��������SK}�͍�X�u_�qH�t��7��5������_z��4=5����t/tM��0���9�e҈��l�~��f�7l�'���tu���0՜q�qq�}�9�q2�������8�wK[8ȋl��^\R�?��W����ӎN������bW8��-�X�Z�#!��p�3�NE�����+���R�G���<+��-��-+�����OD�+�X�R� �J�9�a�Y(�ϳ�	s{gUf�E��f��7#l�9��3�sӲfǛ��U�}W���Rⓕ����4sr�	�˧^��?���?��[��̙��ة�o$��Bm@T	na�:u�A,������E"V����
�UI�9z�(�f�r!�qȢ��[q��aꈝpQ�L�#il��*���c�I4o:a�5v���Z�O�"��]��B�@�ɤvP&�F����{jˋ���deeE8N���j�`�f����Pvy��/�L`T#1Ƚ����`��&��r�K\����4[E��4�7K��$���[��(7�mfE�8�/ɿ����	Z c��R��$�P^K�B���*+�g�Ye��,�m̅��}��SҼ4%���9҇�K�!	���vt�!7�%ל�պ�+Ƙ�T��|�A�[�l��"�|衇k=��#����3�7/SR9�Uc_�����J��%��~��|��߄@��%L�,�4$���d��\����E]�[�B'���tul��믗T(�O�%����bj5_H�������]�#�1���rM�%����ꤥq�H��K�As�C��G>�A8�0�yZ�"����|��K6�	+k=�zA�$�V�.A�� UȰ�J�f��[	'."\��'���q	����t!o��G������P&k��At٤���5�G �y^0Ro���N�١�Ӣ��j�o|�?��~�+_��'?���-_����淾�-63xE�5�D��n��~��?�������%*�f:��p2+�K���S����Z��ig���'-���L����h $��N���݌��K@��?�ެOMM�zl[���2!"���ٶ"^�t�����xr��o���d��Ê� ��Z\����j���./��=1�j���ж�븝I��8:wh����)������`eq�~������N��8n"��kYX����������E�f\�.�+vM��"��&P��Va��[�:��p�~-O�j��p�/1C+�,|�~3�%�Y��E��	F���x%1'!y���@�R�� � 	�m�3�I;�����Q[<:�ØRS2�,aH㧦�99�i,����J�(�v�QV��g�!j�@���0g��C&GcT�>�Qd��������Q�3��:����A'c�����&A�xn��N&ڬ,,ح���d����U0N��%��<�9�=N
mRi���S
|h�ƱX@_è;�V�I�fC95�k�:FksKw�}w�9;H��͝\+4����lu�0�l/������u�]a�8�</ϫJ�����z�|����x-nI�o6���&&&���ggg�
w�#vS@�!��	�M$�� a�Th��۲3�	v����|�eeT$a����Yfa�Q���UIe,B{<i,���"��;�4mx��x;�Roagi�ڠj�`�(͸*1g���h1�(I�OG��0�Ta�R�藜]#V'Q�����))�΍*Y$�B�)s\\�Ly���ih���9�����.���p���Z3H	Jx���O|��K��Ƕ��A�OY�'���^��p
4BA�n��{�[]]���o����={�ԙA{yi%h��J{Rn<-Yvp\0�J	���M�CXrB�d9$v���-zbK�;���b�5F�3\\��ݩqT�d��<�;t�]h4�պjU��'o��ӳ�Q��|�T��g2EJ�DӮ'�6u,H���~ ����>��e@.�Q����<�wy��r\G۵$͐�x��%�zS�������P�<�4p�����c��(���ϹX�AMT߱CN��K��G�JR�g0����Z/�u�t�^'���H<��BNR��!g;Bb-J�G� B��EYXT�Ip�M�w��o{ǯ�bG��kºH���ā#�����}���9�7r��z+����z��G������8����~� �?�o��ݿA�hB�ΠxV*g3_+o�Xk�=#팘�G`g}�5�����\�a�*vhT�T�$�6m1x����:@�<�.QS�^��/������0���N%K��mc�NQ�����*�j!&�68�#����ؐ&�>F�S@K���Y��Ѹ�	�i�����lէ��V#\' M�4%10eZT%j�|��2�'��=q����*4l�dSa�{۹ɞ����Y'O�]V[#5��2rSR������|f��↷�fk��#*-=���1%j��r�^��c'���ĩ�3��f@^�9���q�Xaߕk��@�p�Lbiyg��r�\�X�=�KKKiN,s�`�Vf�	ן�X[�y"���X�����B�r������UCXeVf��Nf�ŵ��Rn߾�&)i�!71~g:+ϼ�j� �"ZT(���˄)��۠V�aW�mxB�m����6;/�N�/
%Q2O��)�xD>������	�.{��~#��?�<�b9�Fɨ����bJ9�2V�� p)��go�cc�s\�0K��D�Ht����1ZC�U�����[$Aq~pZ�k`<�B��e������H ��drI"x��#Ip@A��Ҋ�b��*ڙB��'�:O#[Vq|ψ�L�t����%D1B�&�,�ߎ�
E�xJ�C�R��?�W���\>��<%�I�����.>�+�?3+�����Τ��pGz�~-��0
؋�T2�d�J�r]l�"Z���V	�~-��^�~��� [ʝZ�d���P$0�1�A�o�XS��͝B�E�Pm>�dd�������ߥDI�h,��9B,�Ɋ�F$q�F8"N���S o.��R��4��&�à�n�B���>��Q�5i\o��I�50�������ٵ���6ۏ��8N3q��*6T%�xW�l"aafK�ua�f�����cC�D� �H�I�j���m�D��Z��*c��O�!-Ď䈫B������Rt������S4ž�����X��2I��zT/���y�p�p ��Uf�h��K�Ӯ���z��%T8D'�!!�0I�BI�5J�aO�2�\L�/�r=R�-ck�����{��3�wF1���:c��+�ҩ��Ų-I��Z*�e�h���@Fx\P�۬�Hn��aU����c>h�t+c������l�Cq4#�~P��q5pN�O$?��/�FN����f�@C,(-�9��+c�:4�4� ��k�Q�`^�FɠiS$^����Ͷ8؏5�8DDS�=���'��u�o:��ɰf��V�w�T4X�ݶ�fJ�l�vc���j4�4_H{o��/8��?:��b�ކ��%K
Ԑb��Y��fsj�������M�f/.���K{��=��I���N��c��|�Ͻ�;v�Y!�q�_\\<y��=���,۪�@���~?�����h�w���A�lY,<Uͦ .��ViS��Ѯ���q	0*��`�x�]Vh]�����<�Ġ��K{L�\G�QhC�;�(p�B����f�K�=!c.|>-e�R�Q<E:J<��i"N�g�<9K��f����,4��u;Gwy�a��;���t!P,���	O	x\ݎA�%b��V�/L*qȪń�SCIq��{t:A�%�*�k$*U���HT�6B�\�8r���S(�f�57޸�w�y���`m~�Ә �#Dn��JS�pj4��y�f=��W��َ@����J%?pxm��#�����5Z~L�X��Xl��W?�J�z�I�=�fgg���cǎ=��>x-<�T[�!A�#��a�
%�3�
��D6k@�����$aR>Vn��u\;8���L4[�]�{LXɜxJH�9�͌` <�Vޱ%m:�poQ�#��9���Y�X��t�R�4��X�����N�U�L��˙�˼%�OI�{n�8<�pB��,�\E+��r�p����l��Y2�J��8fA����OJ��4�X:3�����`8�5�Ɂ���7�~�����<,+�r�,�=˜�
ӧ:��$���u=1F�r*FB��2�QFOzY��D�-+�h���>���l.+�������/���b8�Ԓ��$���.���i��?�mkm���[u���%Ѕ�Cb�S-Q�v���#eC3ɣ���5��C �jM�|��_���T��Z��OC�ZBFĭ"��p�B\�X�����h1]h��U1@���N�t��-����xF�F��T��T�K ��؜r[���A6�4՞��4�-�Y&NF:.��c	����4e�T��z����Q��S�9krܓ*g�0&��m�%�b�OR��@�D��,�GT�<��'²�*���Ů�D�V�,���H���Q�K)�ަ)��"V_HM!���p�ĉ0$Ce��J������������y�.q3$$�5ccc��E73>�X�Mk׮]{��i8޶m۴]C����{ｊ��Q�uG-Ɋ,*����,I#��`M'AZU��J��g/�L�ˋ�z]jQg��/>��3�����4LU�R&�z�(U(�M2fqy�a?����y�~��f
���ʞ	���k��I�<B�bb��Ɩ�Bf�h��K�K V����)�(ʺϩ�D^Q�.�=iQ+���	`4֜�b�v�q��o��@SSS�V�������ە�����1iy�|p����䨜� �2[���
ɛ�Y����'N��҇�$��T"V����Ɇw
#�W��_IT3�E�%\��%Y��v�gZ�OLf�(S֫�-�:�#5]Hr���+�|���]uׅ��ѯT^��.� d,�b�ʡ�D�U�ʆ�)~R��(��)�<�(&Q�(��̳�]���UGVy��OJ�����0ՆS�ޙ��9n	�c�-�#u�W�v\�w�(�ޜv-V te���"y�mh�Xk�m�h�~1����7$u`��X�Q��l�����u@Z�I-�%�?�� ��>�y.�`EJU��� 1���m�.�~�T�./K�.���U�M\�6&!�ہ�Gy�]3*�� 6��qZ�����y�!<2 P�%+��8����[l^Y�f�4��e�,�����J�Y/�>�f�1����:w.�{ �Q��JsĆ��^�,�8�B��(��$0���c��m��r�:���R�*�[�7��s����Em�=,�B��f����r����G�#"m�q}�o�H=X[����S�ҩn�UE[0@	DAd�`ϭ_\�V+��V%�xO3�82	I$��Iv�+��	��1骄r�z���l�[���S�9h�!u� �P�����Z�pP�5�{�#�Oе:����jCO5�=5�TY}llb���?�5j��������_��W����i�(m���u�N�:���2Q�{4�.���f����3\<e�N���#>�3*7�J�z*p�e�6W]����*���A/R���1���S���]`CLOe1�;�GKۊȧ�"q3�ad���M��6�<)����xb�g��%5��B���i�g�Py���U:'��t�>ʔ��^Jp-q�@8���&�pmm��X�#���-%9�۠�n@w�"+u�b�{�����_hTLG�;��MO��F������{��~��i��^����� ?x�8�l�ѧ�����ZJQ*�$�XC�	�H(Ȁ�jI���a��U�3����4�=c͎O����`�s�Y^���u>#.WP����
� ��d�1҉R���	��8"�UJ�L��A�SQVs=� MȖ�J�!߽F��s�T���W�(-��c+�}յ��\A~��U����ɰ�>s��Q̄D_c��	ɱVNU����F�<�)E���.r�����aP�k����L͊�[-ϭ�-?[;>U^��1�T%r���A���VyX��u%a�m7e�<&���-����%�nA�ņ̽���|��*mkm��v��X�	@V��jX�H�|��qf�I��s �I��o4ZRC�Pr-	�ѹ� �y	�˲�:^j�J���N�U�Q�����.U���mU8�kd<�qK{|yYNh�K7�A��b���hKkcc�X�R�W�}qcoo�V+��<�q���h�p�*<��+]ƾ�i?�i+��3��*�T"X�>K��ىmᡒ��ПrL��N���Z���d��4��u_��$=����9Ũja͘kY�IR��=�-1i-d��]N���;-�X����+�A��ѣ�a��үZ�촹.)���#���i��ɓ4#�g�HyP0�'F�{������e�����"����oԳ�_�җ��яҷ3[����;aJ�mz�����$���9�ZƤ�tr:��gbbbll���P��^�QD�y�mi��EB�.\9g`Q�MiY��N�xnf�?��L8+�\7ކ(U��QLOY6��m��Yh��$.D;qt�	]�M�/��az����V�D����rW`٩VY�-�^�7 ��,,�*��rD6xS˿���.�r��`-�#3	��[[�?�z0�?�������&�&�=51�k׮c�N��5N���1�,9$��"�1��Yn�Q�#E�`���x���Z���'������%Y���'H�`ŔxB]0�[���/��1�^��� �0	Pz�� ��_�z�F�(�]�5\�ݔ�Ȝ��#H���C��Ov=�T�|Vqi�+]�����r/V�<�6�V��+-U�qѨ�j~N'�����l�g@J&œ������s�D�!���l��`�n��q� ��Iu���/��z��|���6��f�lO�αށ���8���^��46��S�^�:��,p�Yb��_wm�Y�3M������ jE��x���z�^a�N�[�\�N�D���q<I����u��,ac�Y8�8K����:��^lW싺���R�1娼D[HB�<p,و�Ʉ�H�'�$UV@d�[���M��U0�B��Øuz�㊶�r�#�L�lK�pG���غ�C�ITJ����{�%e�c#�z����Z����E����0V�����{���j���M��C*p��a���a4ԙkS�!T��c��jn^st�j���)�ܲ���[��e+�	p���(�	(������xp4"~G;��GX&B���
u�R���8�
���kx�`�ֺ��$�U���+��jo�ޢ�&���m���n�)�r���H:}�_��lߋ<k��r٥�����Zv�(M#eB7�O�V�ݚ��G��f�A}�Y^\����κ�znŅG�ŵI���b������;�ҢR:��ߊ�U���䍄�����(�C�tޤ�I�h*�!�u,�0|�<OR���j,�2����$�`��7���%��<�RA�F�ت�3jUg[ S��(��{��`���T���Z�k��i�b�{L�Dz�%�$����,,������̯2>S�BXX��L"󪒲6���9�T��]��%�u�\��Y�h!�nzz���"����hd�'i�9T~ `��wf8S������cVP�p�*���*�q��z��:>=rw��%f����㥤�F�
�ˊѾge�����e���f�!���THߵR�l�It6�a�z�,FԦI�Wq�D�R���P�.�^9�c�JV�)B�t�H#}["	�����<�'�ȷ�C�<'�%��k
eF���Fn(|�ޟoU�J���X�+�&yn��d>	-4����}m8����yA�-_����[�d�ڕ|`	a��D5�<N���Xbc�X��	�9ϯ#��V�V��mӯ��mb�Ͷ�ί���]���<�N���)�â~�8��l��M&�AH��������9T6�u��0W�Q�ɼ��:����^6؀��s�]A���i�M�j`F@c��\>�`?ֿ�C��ܺ_�Ē�V�C�RSU��N�1���64I��RP��{�ɐ)��xҠ��S� +����7�J�P���xc�{�?Z�VST�A����د��v��n��0do�&��ը��= y�:H)�C��9V�:gP�:LUt���.�Lq]��̠b%���_���ŝNg�Y�dameii�r��.�Zk��+)+)8p��no��ڷo���]�~��_;@�owb>�aH��r�������۶m[��JO���HWA�S:\[ieeՓ��-[�t��D�;Oy8co��`0�ZT�'�z�G���Pq��d��74���>w!y&�Q�Y�d�)5��u��:��%@~�Scb>�qL��]�Arِ\JS�נ�p؎=>>Ns��	8���P�g�|�p�E�vtk�J+/�+�2^�$�0�
5�Z�	y	��t��=N�����\�����v��Z�`̑�$��̄}��5g���x-)�.0^'�Í1S?]�mã�@�^�ȑ#�f�x��ֱ(xm,�b#L�M��P�]��H�"��3N����δx��[z::L8�[S�P��$���mX�G_=�yq��9O�חl�D�s��T�v�K����IQP��%�R=�SS��;�JZri�6��ҧδU���t�ٚ6�4���(��\�e�ٸ���P��mb�Ͷ����se�p{�`^Ҙ�v�X�,ꄃ��
�(IH��%]%I��D�D\ױ��ȤJ�$�%��Z�����e+�`���Lj�ҒW����6��OS����D�I�D0W��=��O/�J��
��t�iqa"{�b�����鉤���v("Y�$1��kk��gb�u��E�x��r6{�Zf!� �$:��ьV�L�m�HU�����v�j�enBko�AdUFY6�j^\·es�l�v����9�7j�-��a�D�]���NZ������$2�Oc;{�3�,�|�$K����p�\OH#����d���Bו"T9)%���Jc;�m$�D��	�H]�3p]d�DQo��$<�F}fvK��@��k~c�<�s��+��{��<J��4V��$�*�A�Mgj��j.�,�WWfg�/��E�����\��1M��f�Ls6�8����ĝq5�{�����dff���~@s��K���؍gy�����c�\U�O��8��X86�D���EvV��\6x8���Ǹ|��SN�ri�U��{�'Q��wY���c�r..#���T#Le:�S�s�Lм�8���:m�Ǧ''�}��R(	A��6��>,�(T�k��/��`"1�+�z��N��7�N'8�r����[�g����ܹ������|�Y��$����{�Vo�a&��i� p�	�i�9��ä�F���Z�0��ݻ/��Btkkk��i�c�&�3�0Z�gՏ�j�`��>Ty&��__�)�;i�PiDi< 4�����|ZH���!�?������>e�0�36ʿʀfEؠ���rN�֓��7S�F6��	�0�V+��B���Fs�@��_s�e����<C�
�j�D!J���!��L�/"�:s�U��ϳ=duzs�
�*@r��.`��c�!|ʃ�䂕p���%�8F&���6l4����]y�+���Ρ6[�6��f�lO����Uۙm"�8P{rتd3K�A�]�p�
悟��غu�eR�N=�����1�ifuG�$�������1/�)Hعm4s��eL���۪��?��h@7�
��t�u�z����MZD@�^.z�=0k\�멣�����k���ol9���Ա�q�D�CH;I�f8#Bl�pg49֒\8yR�Ѩ��U/�V6�*��X��e��$�[��o�85�-���Jڕ��
s6�Jb��{��%U�*ǡ�!8�j���I���"i��$kv8
%�|z	���)i�L�J�������b�ߟc���6az����K��S��m�{=d3jT�����Z.����8"�m�ԍ755����
>|x΁��s����W_���?~���8�Gh����*|;QB�в���1BA�fO#8\8s��ޥ�%z��	�~?1�����c`
>z+�/yI�Boff���["�*��\�U�C�N*V�!H�Ho*����G3+Ϝ�y$�'>�,@_9f�n#�M�T�C����Eb�|�IM�k�����d`��|��u�.�)�qqLY�+���B����@J� I_I!g+S%��b���Y�I�!�aBؾ}�E/zю�]Ir�q�Ko~љ��:t(M`D��T��$3J�	�2�dU�"�������"�_	���nӔs��-���Vszzڀ3VÈ$����t|��r��Ojr�$�QN���"xPl�9�2e�Mֳe
�&
Ǒ��B��C\���w���8�7?)͉e�Q����w�*���]ȕ.�cH
h���ƈ1t��:�����CoYQ�y�l�AAB^=F�1�H|G�f�j�(��g�4�ԶM��$m��r6NK=�U�lU��yVy��^��Z�����=��ֳ���ٞRg�I����,I9U�J-΄V{zR�醤�*���v�}ŽHѦ����;�Q"�?���P':S�jv[��O���Ñkp���(eG0�EQR�\�����&N\ѱ$���2)��3Ư�F<[�9� i��HU%���MĎ���Wc1��sh.b�t#T��LF�=�#%<�����NƩ���,�`�܀�sS�cD*vm��>p�{�bG�w��c�QW2s<"��k�d�3�&�v�x�_���W���=F��p�s|6�F|<pl�}4s�BW�F�p-U�,���L�f����4`�5r�����嘢�]�*�øX���S5B��\o߾}�>�Щ���-�I�pY{cw��B��B����(H�9��r�.�W�ڦ�H�ȑ���]����;�=1��.���]M?셮뗉���P�%VJdT�1�1c�Ą��P�	*�s�&$��˧��������|�D�fJ�kf;�E��ю��i�Ư���۷�D�c���HW���c_o�����$�{��ܽs�}��❻v=������|t�{%!]�10�fghV�Vzcg˖-���@[��������|��)4{��=v�	�G�\R��񐰜Ժq,�,e�ǈ��U��f5?�	h^�X{ѕqAb��R!�)7����Jk}����"ᆿ�:�	��L�g�LUb����p�hf�=t�,yp��0��[�0�j����ք��uC`� � 5��L4{�R�Ϝ,��:9]��1�h^&HVCy�L��La1��{+�^v�sF�L��(�����'�x¬e�Q��xϥ��)����a�/�F"�b@����ڜp�ճl��x�p��:��������T1�pOc�H���0{�o����l��hϞ�����&�����ٱsw%sss�Fu��b�)�N��2�wdȚJ5��s(v�3nWS�ka���H�(�ju�Ա�N��w�s����ujM��23[��}�����E|�p�|O��QޑŁ)˖ĉ�S ���B-g�����We:2���2�C ���ba$B�yb�Gʩپm��j�:��9\�P�4U)�Tg��q���sjU���?�*+�����(�;�*?�6܃."Z�Gp�Y^��Wo��x��:�K�4Ugz����je$*�������_|#(̵2��	y_���oգ�?]b����M��m�Xk���6����������355�sf��.�~�K���J�.-�geI����߿���m�6RC	�ONt:� �:f׮����J���ٶ+A�kkk�kOLL�AD����o-//�CI�9�؃ܪ��l��`{5�ϵ���P�7L�SKL���'�&��Z�*�s{�ȉ�$�X��[���\3�g�KX�I�}Q�!HQ�O&������<{��5I�����wl��!?���!�ˤ�V� G��DNE@�&���ʭђm�@�$�{�=R�|h��0���s]N�Y΅ģ�|͂o�ծ�U�ؑ6L0ft�����L�(ќ͎sf!<�W��VEޔ��0`,L95�ĝ2Ed�	%���ƚuO�p����<?�f��c�iT	����G=ztq�CS�G��lA���i���D>Lo��i��=��R�Ç���/<�hxH�a� :xvv�u�{a����?���zb�G����)��=y4��KR#M�T������鴒��E�"�kL(S"�	�g��=�>��C��I���+l���6b���j,.�ch����q�lt6�����̖H��s?�h�_6<�lpu�s	��y���;.68�p�Q�pH���63AG?~��E�a@�5�\�~$�G6�a(~�:��z�����iL���K��1�k��EK�1v�5P�m~�G��LN҈9r䮻�Z�_�3o�2C�C�K�I/�;rFr���y�9�#�3�2���l�=�*ߏ�T���H�}K8������P"�i���J	R�Q<{�yܢj����r$E&Y�<��|T���H�L����Z*NŲ�"����<� �sɛ]7�yᦆ���L)78��i��[��m�X��[EP�W��jf�:o��Y����t������A0�Q�b[N��U�ML�gMn��ܱmϥ{/���BK���Z�4ű1Ķ�������Hx�aؾ��#R�?��������Q���'qL� mä&z�K
����}�رz��t����Yh5�n�@ZU����6/�c��}I�![��H�_)]�j��b��=t�X�n�%���m�6rnP��>�wდ�1��8�A���'�|�H)�%���cDc��}��C7�C;?4vfP��͘��F�o5�c}�{���o��u����F�3�3����D��m/ �W-���f�ő���<E����u�d�\�`|_��8)8\��x _N�!��X
�q�j�����o���U?Y�����H�ST�Bw���HG���Z�⟥U�����{�T
�H*鸒�UqI~�U��e#ߏ�I����|:�%@�Bo՛��.J���y�� XC0�}����X��}���=�����w;1j��?q�K;	G]q�%ti�z�4�Z}i8���i��[g��3�c[|����M�޽��s�h�������o~��&�[nY��'O��dV6�}���j�Qa�fë���N�#�5����F�&ݎ;����'q�_�o�&�Fk��"����8��a�3�)����gc{�@���L��������1QK[�ùp�%
7�s��ޒ�����5vl/�3��4���B�&x���t%Sg4�6_�V�4�i�*�^U@u�(C�\��$�N�۵k���/C�V�#������aI���j�U/~!͸��V����d �^�� �ƫ=:þ�����i�K��A���+g�g_4���8��5�9�%xs�ϼpff���t���ضm�V�ע4 ���F�.�&��c%Q(��H�8O��$���fL����i��I�]�֛���6�,�?H3�Gh��d�]�5�Vc;�l��Tb�D"�Mc,p��6����K'���כ�"��F�BVԕ� �-U5�Z%M]5$�`�����Z��g%�ћ���6�֓��g�l?S�'��6��ȰԮ6���D�'�A�)�}����~�z*�DÀ��p��N*L���4=5C�=|�0W�lshS���Jǈi1!|͕���J�+�UR2��%�^����t U}��0u���ٕaU�2il��Jk�%���ϭ
\'P��V�,s0��E�a���c��	��ɶ�	9}��rI�1�/J������f0[��:6����&��r�-�HOBw�f��:��+�9}s-,�L'[��8)2�=�ߏ�5�O��V8[/H��P��1�q	ȑ����L��������krN�|�� +�Y�G�]�8�χz(J����٩qaQg����H�I�`P�b�,cIDR���4�_z�`�Y��x]t�Et�V{�F�ךƥ�j-]B��}q�+�D�S�.}��tdg�8a?H���tї���K�B\%i��K�_!�XZX�ҟ�E���C?�f������o%x��z@�ʚ��e��8�.˼iA�(�x��k�|NI��h���`�z�,F&��Gy��
�H�B�y�V­��3>>g��Q��8��b��yǅ��Ա.V<��J�ks,.Mjd��!�i�J�XQ��������m`�x9�o?���?e�3�<H�%k��������7���D�\�nO{�=�v�C�@A�$@T�+ ������+�B�+A,�φ�,}�J�B���*@F��+D��$$
!$77������V�֬��:�ޛ���ʙ���>����\�s�����C�5�� ��Ŕ�4J������׫S��=�MK�`b��-\%��ncK)��;��5�9r�vA�}��R�G�z�5'�|��|+�w���}���&��8+O��4�	�n7Q�1�Qk�d�3U���4	���Q���Yv.���P;���O̜���h:�i߻����c��\��z��W~����Mg\T�y�1�i�r�y�}{t_����8�=����iar��m��+�G�sHQ�F�����J���p@�z4
����<$ Xs�:qj��z4:��� �I���9٤�B����� �v�^X[[�Z]G�0�I���h�k�����Ven�>�UU�O����0���8���/D(��e�8�%E�~Y8�r��"UQU�ϜV�S;gxf���3��:'m&�{)k)�(.���=d�d�ӕ���+_�R�<t�w���W&����w
��|8�T{ڙsl'p�YL�VĀg��f�U�Ut�E	��ͺ��L
RRvHS����6Ԧ(��v��Ʃ(�cv�A�I-�k�C|QF������KM�8m;ff�N�IW��mݪ�r�!c�D�8����=k���=�ҔP
�^�A锱=^��!������vTR��ސ&��hdRSFq�vfh��zZ���8��o����K���GOt��5=7�ĉ���g��%e�i5�ן�/h:�h����3����fo���C��G߾��}�fg�����h8�"<6X	������\v���.�)�:�v.�d-	�8�
u����3�!��zz�AޣY�FJ6��`�X.��.������omї���z�zj�>��L	����k���RD��SjW�٪�W�����+G��YD��H�)GFg�]h��d���-Qe�}쥩�.
���58��9��Z��Z��R�E�i+o�{h����~�q�0�
��83j<c�+?F�Ngi7�
#Q��Bs�aG��n�_\ZB��G �=���L��h��:n[-�X{}���Đ��7��
oz�ja�<��3�I�cn�U�t�4�@%�^���{�O~�/��,..�Y\"�|��)Z�߾�n�vF�4���V>*�ii.�'��#`�1*�@���l�Ÿ<[ � ٞs�#�{V����$� ��u��l�(6�z9-�"��Y�"�XE����m�c��HҪ�Y�'y�� �Y�B�eɓL���x\O�}bc�+�+����bˏ)4j<?9�;s������v��?�������v�Ԧ�RBA'��4[s��(ZfRw�˖%�M:��V[��,l�=q�i{CNY!��ߝ�R���	��u��fR�����m��n��Pg���k���b�U>��	Ȕ<(��P�_K3�r�vH\9����m��Ј����i���I��)�� �^�H'��K��s�����S�qޗ�����ٔ�d!�t������覭4�U���?�93k4�ͮ����
��zDzrb�����Ns�|��<.Ҥ3�2pdQo3�����cÿ��h߅Z��5��(�hņV$�l"]QA��]�X瞻D����\S+Z�E�<7�.l�`��ݳӳq|�b7�F֊��Z���B�L��+�l�Ȥj��� �kVWi�e�ųAˌp����H`��<�����������{�=���+�P��S�"�f�sf�������}{�� DL�){⣃ǘ �p~�<�%��CG�4Nn��tQ�KDX!3�!��B�6;�e��p�P�c-�X���N��)�F��Z��۬���r�����aX�A{C����A�v2��S�#��R&��r�@���V�l(�����$Ć����{i�h*!y.�����Z�xjf_x�2��b�A���j��Ǐ�6�G���U�9hb�����)�W�骸�Upr�ã�37�5�8�k��G�&��H�1�Xɼ&�(�'B�<�9� �TYM֤%�+)T7��8<�Zb�=���$Ɲ3TX;����?m�N��VKu=N	��� AmR(��A(�N{�mk�����;��h�2[|L��i؃��uf)�ʭA+�gcŁ��]�cZ�ӵ�2��?��diii~f��˵�5���.�_}� wh+㔃��Q�::A�f��H�Jz2_��s���$5痹�񍂿�K��
���+=+�۵45������g���-�� m�%Š���.=�_�̃��1�#�jDQ)͌g���0e�Ŵ�%f���#�WI��h�`�'C����m���w��?������x�"�h���Ƭ�f���,םjv}�[�t�3�}�N<��ۍ��Z�&h��3��_F�������2E�b��=�#?�.��}0Q�\��=���.�g\ǦH���W�,��I賋�����[<x�g:�f����e�E �
�	�@W*U�!g��wj>�ŹU��8�I+�7z(Z\� TiR�F����ƕv�X��O�"����F���W*��z����ztó�}э7Z���|f���{�#B`A&���l鶛3�E�8�$'�}C�o5���l%�d�"��==Mpkqa�����5�8�{ӭvӛI��5X��7Lu�����v���������766��I���ZM���*.��
�6����џ<IH*�®9Bw�gX�{�e��,ؿ0��զ(J�0����xVY�;$;Z�,'fGb�L�O�dG�<��x�UM��8����ao[J.U�hRdbL�~_�Ϫ&X�@j�+읅gg��4(�mI���1���tgM6�(�\glI���!�솧.!�d�k���6W{t�9{�_��'�ӳ�M`�J�� ��K�܌����"�`�bj8�0)-����<�a	��2!��T���݊�V��tըV�+��,�77�u��,���O^�"h� ig4J)	 ����無��2�c$�́�3~dX��	ZM�$�Z��۰��)��8��é�N>�zZ�q"*R[�v[�`k˘�"�G�v��+������L�۠'�<y*�*�Y�2���-m��鹒����^i�w�K�HU�J�XK��w�xhۆ���O��`����C�����M��-��*� ʜ�p�mn���fsW�\��fWxo4x�K��G�R��8��q�yr�(
l�!{�p�a��yS��IBU�0��@U�o�ˢ�x�F�c�-P#�B�4�3�O�Q�����`3f�\.���(9͵����y��Cd�CT�"���Z��ø<��޽�Wz�<7�q%Acl	�U�vt��"T�m�>��L�������--�{�}]I�МC׏���V�C�#�~K,���<k�۔>+IJ�'�s����#fST��=Pqd����ۍcH���H(i�`/(��2���WDst�rd�BJ�����n�;^xa>�@h��bYG������F~�&�8�k����cr�G4�`��Y��.���ǧ���$��	��6��p��&4��1A�>�oc�Rd�S�D�����q�5.��.���Q^Z��PY� w�z���H?�����`m�.�0�O�v��c<�j��9�`:� ��Zx?�kwI��d�4��2�Zx�Wס��C)!�������,&C��h�ν���#n���!)`�"l(z.D�j�I��6��n���JTZ3���1[#}�փ-m�0�!IX��tvn�&t�����f���I �fM,h�4`1)���0kE����&G��-p}VJ���aį%XK�+"r.���Y.�������i�	<�ն��Hςq���Qv����K�|�w�1A�.��Pf>�8���6�ˌv���T���1{���>��oˢ��GR�v��j�]��총����k���͈�*G�b�$�V�Vu���I�m?f#��Pu��o�)b��=��rޗ㺖eN��.˼�$��V>���<T-(��!�"��#�9jS�</�Y(E�3?̞$z�C�>�G&��`���ط8ӡ��:-R=�g��ֳfƤ��~��7�-YQ�M�O\~�d���Ei�	���i|��T�\��jR���HUwlD��m��n�8�2/�,Ƿ�h��a�ҕ�Ek�Tت��@�� ��H��q�<����JY�V'���9YBS7���%k�_���*Z�m�xT�.Q�xDJ�S&h%�����&%�[.G���GY�g�wA�29.���RC&O2��^8�c�	�9.Qj�i�l;3����vkv����Ϩ�/3#"��رc��g� td��
۔�&߷�O����XmBG�H��X���I�
L%e�͓�OA��ձ�yR��O�3�l���D����(�G7BU�+�߁Iv7|�����=�g�v����]lA��x��6��a�ޮ�TOV-�����i�O�U����7��K�;TU�V,��l�*�F�P���X_V�(ۦp��r�LD�����n�S͌��:{����3��W��{�w��J�<׏�݅i��"�n�e�P��B�s�Nkzf��U�Fd]�Ф�-D{�qѱMC�u<2�f�1���O�gw��K��aw�e�Gc�p�W�!飃�@1�}6�q%(Q=۱<�l��v-�4��ٳ���9.�p2��l�ok����(L��>h��(� p�4�(\M"�nðм�煓US�_��.Kr��:t��r�Pa�G9���]V ��V�~>$�:b�G����!���&�7Ƌ���2��j{M�ٓ��]*�����~8���$��D��̨͈�"�5��a�M��QZF���iqHv%(�������g��������IRS�}/s����]�7��i���"#(�f?Ώ���T@>.����I�i�Aɏ�c8qP85!d%9 V)iO�#j���kP��(Ui�];58X�Q����Q��J��,�$<�$��<Դ�u>ó8	��vD+�uD����J�s{�Ϧס�L�o	r_]'��N�A�K�Q/�3Z1� g�DA�X��������︉�t��:��ip5mR9�ǝ��ϮM
������i��=S{!��HF�x�֋�Yb��lQ�+�-��6=�aR4E��?[��\gC�`�5�0������E՛`�Uc��i�Xc���4�mo+�W!?�����5�-\�ũ�g�E�|&� DO��flm?38�T�SU���#g#88π�c,g�L ��w��!��ԛ�� Uz	w^}/[9Q�f��RW,[���_+�Q���E���SX[����e���h��x�`�n�	�"��⧓�@��R�e���BԖ�4&��GY�3�>�j��=Τ�d�ʮ&L�����b,(B�����cI-�~����ů%�a� ��+�+�ߘ}Yy���.���q�P��Yu���ɓ'��{8p΁sss3^ާ9���>���s�d���I�;��zYz��w֣��a8�mkjj��W<�. u:7X�n��Cǯ�{�]C9�����s����Fx0XkϞ=^0��iS+�ͫM9�Bg�~l���M��|�y�5�I��i�����LM�Ȃ��r�
��e��k;���'�H�ꪫn���Ct�������_ZZ*����~���q����qz�����b�;��4�Q"�DW�PR�KR���:��.�[� Kg�����!���,v���3����BvPij�ur}}��f���wZ`��%�~�ܖ����4_W�4���(Aĩ���K���d&��#�Z�������#5=���'�NM-s
mj?LU���*m��2���8�0fZN�c���P8wLo���B�#&���F0�,E�?UwK3���*.ll�Hn�C�ї��F�GJ�>�<pW�	XLN�d �cь�8v^��<���D1�hDw#aG�x��Q�����u+J��&�R�>�Ͳ�Q��*���!�!�
�����o��D	�;}6c����|�.���I��Q��t��%���	{�ݚ�	��l��۳[�*�f}Y���ifCmu��Y�D%FcH�ur�^{��n��V��I�҈�_�z��u'OF̧ڔ5�.��`��$��U��Ff�keC�Jڡ��	��v����q��$ר���TƂ};�p��d!$� 7:���ׁCL��A��d�}F�Cw�M�q&�uʹUg\e=I$c�pؕ�Һ�[$�I��J����8�G�q��h�q�<��!.6w�.��x�Pވ�Z�O0ͥJ��9q<���p�)}c��"}��`��Ǒp��Sी�*D��.�8�\F�� �����U��5�BWQA�X����9	��9��!,̬`�m�S�V���p�)Zy���t�G�g;t�k���P��*ATe�Lg)�VA�72�Hɣ�r��yH$�I����k�i��N��y���*���EH�G�+�u��2����KS3�r\kG��K
L������Pq���x��skG��K�I���Q��*���рPB4O�-��I�KXu�b�3�4��J8��4�+���4�ke�����hu�Y�����ſ6�"�����gH�Qyʵ�24�S������w��p�+c��_�b�,��`:
:�y;J��5��n::�v��ān����ӿ�`�>h_����~�Z��(���=�]fM�R�'eZ����6��Z�K;�v�=Z�[�e���brG��>���L�U�	���`F����*L�����C(� �*Fi�}�/�Ea�4��@���bh����U���|��m�����}�h+��	�Q�\�͊ܣnٲ�uQ<&-r��B6�bn������q��W�XǴ佖��J�UNn��LBr`�i5I&�{��ۤ+���WY!��m9��^�9�ƈ�۞r�u�/]���R��*���~n��3���NMӃ`e*�d��<��ʅ�s7�-]�j*&��a6��E:n�@t\Qt� ��������U�#NaŠHP�=x���%�vA���;<�:ؚ�?��ѥI)�H
l�Ad^X⚯�q�����֤��l�ev� �B�b:���Y���̔[�`��I�|��n�ws����I��i�'	L�V�/��O�IL�H��)�T�q�0���"���;4݅�ꕰ��H~�$\s�x*��� ��� aH%5r��+;QX��E$!a��MErW0Iά�d���{���e�ض����[��F��3�>�L�(�5,�[a�a'�c��ʑ��{���i�Dy��������[FB��i�$Or��̀�(MIr6i+ ��n�õa�F`��v]ߤqn4}:h�y2d*�y�)v�1%G�$>X�m��R���K{b-U�kjۿ��5��&�?+K��o�1ѓ�����@,�7�M�7zL8V�p�ժ>�P�1~@}�D�Jq�zF��`t�zU����C�	�U���όD*a��\���J-��Zq�
dB|EYT��*�䭤{rl��u>&���`'�J�1��d1�㈔7�C=�lǤ��W#��w�O(ۧ��ge��� �(Em��q�ݔROF 1���d.��W�\���`zו�����4�Y���V��>�QI�d2�Tz�G�����9�V��7ʑ��>��B��@q���`n��矿6L�d�x�t�g�)'XȔ��U�N@�.�顿Z�S���r˰����8�����/|Y��C���m��q#�>��{Q�w��V7p8/�O�:u<�O���j:Z���h3������.,,�^z�]��-O�尿���6��F���~�[�'O���{�5j����k��΋�}�ɧdK��U~?�z�l� �w��L��_�1׏�����W�������I:~��!΂�mIC���9菣0��׾쟦��h����vs}&�96<� ��-��W>����T �X��A�~�7��ޙ�=s���;;K�����v�}���������<~���il����<��W����c�<}i�Ւ\YY���={��<~��|H���9a���?���6�����_�M�������X{ΐ�c;�L$;����(� ���n��� �W`ʵq��,^�%3� l~҂9!H԰c�L!���D�����n�jj{[�X��:�U�EFЅ&�� �yzz1�12T�Y�C}���!mD_8 �%�tZQ��6a-�u&���Ւ�����l,��=T��b��r���1C aL_*��6��&U�fؖ�܏ �$I%����L!b���Z��>l;��5μ�-N.�����R�qQ�\�c8�%�qzFZ�j|��IJ�_��[[[]涍c��\��kH�]�K����?������K^�ZS��G�>D�j��K�S�`�s���=�V�WYKU}@�;�Z;m�=��x�Z��W�[D�Uc@b��WRK���<+��f��t,R��qy&VS���C���j�DmDb�W�YGlb/s�.��Jb%ڪ��pN$���=p߱�*�B��)N��ۊb'1~�):k}�M9C����0l��h⓯'��f�,�;K�fGa�� ��j�是����|g���R��nGJVQ*����r�2'McFY9���$�*.{�h
������ZX��3��4�� ��2��Q5��㶭�rV�L]��2����"�B	 ;�G�`����O8
x
�g!?�V��i�"�Ep�@J&!�+*Zb�5�_�!k<���t�g�!�,Ƽ �<̈́"C�u���3�uk<�T�W�bH���+����p�sx�v���3�BZ��!-��NWe�� !q�0x�
�i!lԖMJ���\O�x�jԄ7hH�[|Z-�Gxdŧ�����t��Y��le��ND�Uj:����^Z!k'����]��ZEm��BGy۱�����:X�U+��L��8����a��HeS���2yhV^e��T��t<]V/.�z9�is 0��ꅡ��^z�Vk�$�����A��#׊=;v��:p�{.縳�̭�6��X����N��g�Ώh�ԃ�*�B�H�p��/��ùF�r9?K��ea�K
�ɳh8\]9q��*W-����[̌7LJg��5k�+�Fx�eg:sJ�4���oY�|xZr�0:Jhf����l�333�t�s�����9x�Mp�U����Iė�mD��jϾ]�v֎��pY���ea�K�,5�	�u�@.i���Ei�4�@D!5 	B��rS�v�b[����b�?��Bc��3�xH�9�;�y��25IW�a4�k�z;��VZ����D\���0�І��W���s���6�+eq(8��fau��m��$c��-EU�}�N�gm���h=V�>�&�C�I��D����t��%�7|T�s����4�b��+}Ǜ'��ܡ ��J7IJ�7V����|�����k�s�;^׳ E}p�k~�7qR�~�1L��:S��|cym���K&S��6HtbC#�I8�P��^���,���z`��ca��f�~��W9ڢ�1���#�d=d
z�����=!UB�V S�Uꅅ]Q�p��i3L��Kr��3��y�\�=�����]gjz�15e�AI�^[��|�a+��JV!0V��	��v!�ƪ��7�N�i��=�VU
�,I�	����=Ϊ�"���)Q!��`�"Q�Y��!_�O3F��`� S�b������d�L%畄&����%:��������������	pLI��n�]���N`	(�@���f#�QLq�K9#-l����t�ͫ��:|�	�L�כ��;�����d�"��e��)$�ju�M�^��e����Gk��~�S���Xa�}��"�>�[x�����8�5��@��w�j���y�>�~�/D�*vP�tLJQ�y2��;g�j����̄��L��\V�&�C�?|��.ݿ�f�@P˳':��+Se��1��E��#@
�p��(X</�'��]��lbXZZ���Ͻ�
�i���F%�v����y�[o�U6���*�Σ�x��+����E9{�7vM�Υ=�I��3~��A�ᦘY��T�9�7J���J�@w��f��Y@��I�R�����@���.V晫�Q|��ʜ�8���2Sc0�:k�k����fg����'��"E��+��t��&�(Isd���Cګ�
��%΢�L��={̈�Vӷ�~�B��P~�~����i]���׿��'��+�z��ݻWO�z����3��t��!	9�sN����I�u�9� �ly�O����j���\�w�^`0��I��07���#���Qf�(���Ű�☆���h	�xG�\�Ky���wYQ�k�#�Yd�"�1Me�YF32�y4���V��X�c�CzM�?�=�"S�)�p��}��ѯȍ�  Yj�R����U)>FLY�#q�f`��E	�o_\v���W\q�מ:���8~���4E��Ũ�CV�2�)�{���jo�.�m�T��e��2���J�q���YUT�Z���IU��O.۪�[^�X�٣��Լf*��b��2�vv�`I���>���ѣI���]�vi>J����4��n�IOz����'?��hD�Q0$-i/�ɟ�	�Ï���_u�U-ۣ������5�,�G!���q��bբ 9����-g���!�i;�m�C�U�a �8A��Ҕ��?�ο�7���?���8���f�F&�B1�������7�x�>d+��L���.;z����o����_|��m&��'8f|�ABI��$���/���/����w�����?���~�h�	�|�/x�>��OGC:��,y�����W�B�ӋЧk�V���gn��k��~�w7�� ��8A�2��5����-�ܲ��k�g��M�?�E?��7�D��0���֔:/�F3 �_(�۾v��������_�#jB+�JU�8t��N��|�^���A�T�n�k���8r��ӟ�tҽ�٥#�����QS/��ַ����|�m��F'
ʞp&�w�u������<�9��-q����v=�o[ja|�%C�R
MF䕜Y��tz������p�zN��ĄD� �������Ȕq������)���\V*L�Q<bgnf�cc4��V�t����Κ`t�'�M��5?5��ģŏ����ɒ����J�Y��FiF�0+�x4��l�r��-��J!�ђ��4��`U��iK`�S@�$��g��I�"�i��**qGE^x����=Kt�Q���:~���-�.l�<d���ڳ�_�N敩�3?vM<�����M���+U3Q�N�s5%��>�uo4��Bɢ:BXÿU:�Љ^l���i_EE2���;�i��i;�c{Aa��gt��q�ڞ7:�C���_P�ź9�*3�I��H�w�؊��BcƎ�G֞ES�8o����T�!��U�
__��w5'��*S����e�'a#@Dhq�q��3v�ͭ�a�	U�����EX�IK7h�:�U#��"5�#I��Y�]�S�b/����rLb�_��=7,$ʪ��[�lc��N���-��ڻZss������7�8C���,���<�'�gv��k۴�8i�ɀ�͆X���F>8�T'��b������UQ��I�/�ULˎ�L+D.a7c���YQ�s�>�.��LhXy��N��ܳ�T{aotC�[�����)6Dц�S7'F�3�Ð� ��r"�����X�ؤ!OZb��R�t{����+Ƿ�C��JV�k6��$̀�������U�>�5mő8��ěY����jA�Ѯ=��M?�i4S�X��o��9ܢ�	�4�}�<@8'}� C����$���.Vp-`Z-����}���|kI���
G<#̓��q�ҵpl���3e��&r��l��J;��t�dϳĢ��Zݹ�N�G��	s��|[[ �/hƜ h��"ȓ(��� I�$��%7���{['WW��=��m�%q���p-��u������v	6튉Ym���">v�N�i��=�������*I
��!�Z����L�}���?����@�D]�r����oll�,g��W���s�=�����O��]��:h���}�k^�7�i׮]y�	�J3��"�	W9�#�χ?��뮽�'�'����Mu�BzN}#���}����.��ry�q�@��J��|8�.yA33S0�۔�g4�����Þ�#�y�kk8 A��i��uH���nC8�]ԟ/~�����o�3�!V|�S���[��xG����t�.--����[���H�g��0�3g��GA\u0!{��(��қ>��a&�g�T�q����ur��[ߪN+��t����Xk0�g�&t�{�흛�����1&Q�����f�������G�?>���q
\�mt�:m�'�[�_� H����(������fffj�7��"�����7��RU�k�?p��8N2�}J2>�9�V�����B�۬ӕ��:Bź)M���U�0i��6ܪ���M�h�2��*���ŵ�b����q�F\���*�]l=��j�+��V�Ԋ�������q=4yqF�����Ȍ�~��(���(�C�͊Q�[|���[��့^��e��;� ���T{k�?;�k�i{h4Ĥ�s:�D�b����f��Ji��6J1z�$EU1B}ۆ��X+�?$`���SSS��I2�v�m�]f��Kþ@_��o~sks��\�n�}^��S����x�3��9��@����<u����ŸHF�}w���.K�!�%����슻⑇���=�1{j�u�H��v0=�RU�!R!W�.\��4u�q]��͞@�%���:{����3��<d+'����.�]��^*u�����g^r�%ᗾ p��9yѿx헛�����j~�#���*8����r	���MT��9r�ȗ���~8;;K�>�	O0lsI��Sr�<�h��3��f��lܥ�t���WG�k����ˊ0�~_�f�blw����0�¶�?tZa4*���� KUi�3m]y��m�xt,f��1M�ݳgO�W�k����i���n�-6Y����`L�E�uu�my�?��y��5�/��|�=3�$�{�}�wuj�cA��k�(b������N�i;��ֲs$=��z��l/MR��o�����0 y����������?�:��7�q�#\��M��7�����[��o��_�}�ʗ���O��M?�S��f�&)H棖H��c�����}���ޟ��_�����L������W����,�8r%�S��(5۳�z���������?����QkK��Z˛��˟��������o���2D�Lm:�f���_�%�#9HT��D���-yP�i��J����F�ȱ�������|%΃�� �9.�:n��Q&r��i��%��	4�u�H}��[f����>�ן;��>?�jʹL�Z���_��;�]�n|�ֿ~�S�dt�X�_������7�v�s���k�T�Vd�)�]p-TǎI}NJ��.�m�c�LQ���J��������ڀ�MW�e�Ŝ�����%��؅���Oq؇�*)c7LL����AKˡJ��/'1�wV��9���}tn�$F3��Rm�]LA<�%�����򣿇*J��i��a��
��8L�t:β�|?��h�G�x}�ɬ�8��ܷ���f�uŮݻsc���Wl�ScU�r���U�������ar�VW������N#̆��teB}�o�����0�w�]C�8w�h�R���m��9�K�L��c�0\�&`~p�Za.R�aC`h�q�i6�2$�eĦ������������4H륵A�Y���^1�-�a]����v#4����C�߾����w=CdZ+ '�U��=���	�.d���x�Ӑ���x�i|�rP�7$5�Q��AѸpi��n���=����rv	�`�:iH�>u	�W��cG�Y<kO99\e���� Ip�����XeYK�uO��l)׵�a[c=Ês�*<��*�}��b����ͭ��V��Co�w$9c	,a5P�����w���j"26Ni�����`�����H�:��r����~����'in#� {ڈ�J��i6Fz�9��y��Ȏ�:��h6!���j"u�IF�f2�u�����u䶃w�Z��#��	�3�.G]��E�T''���J�#���ۏ|%�4���m-��5�p��t�;�T��Z�� L�'N	 +�T�Uѿn�3F�����P� 2_Ȗ��|���9A#8r�]�=���x���r�sw�Z/%������P�ʓ<1�B����^�́�N�§��TtܦŠ2��E�x��V�1�U֖�g�ǱS��P��ǡ�-���e	�N�F���"a$"���}��zn�Qy��Q�8�O�ҿl�b����Ջ��O=|����[o�����&���xޣ���d��i�c5[]ۦ�ۭ�3��̃���g�?��^~��{w/�h��	����4�Wf�,@�����	Q�
�|'C�B#�Ȕ�V��!d� �`<��g�v�r2+4x`�d�*���Y�����,u82_s8��e���p�p�;bp�W\$�-�����k�'��X9e9��sZ��(p��uph���Rv���O����!���뮥��_^]]���U����}�F��H.僘��F-�%tP^g�kÏ�h(J�A��Vn�y�p<fN�pP>W+�Q\�VU,T����j�;���]T�Yл��U�9߉$���+_���p]��g>�����F�)!�U4�o���'=�Ioy�[���Xz����W�_�/}��X�m�Y��Â�۔'���?�����rz�UƔp
�*����t@���]���>W��˿��?��Gn��e7��%/y���뮻������陙�{`R΍�R�V����~FzCI�b˜�	��fP�`��S�r(�))���!��\���F��i���)�׾�������{�+~8J"R�WE$�@=|����UObbr+ɒ�<���~���_�4]���J���K��/)�;��wfVP)i�W=;'�s8ԶrC�!(ґ��h�E*ċ���VƵ���6�2�ܮ�<���mr�w��ٵe�qL��]1��q�P�i�l:!qA\SNe�9x��ѣG%
e�3�{��$����������=M�&7�5i���J�g`�d)��`�j�`����Y�n���h�:V�,;q����K1J ���H�Q+����׫�v�6�>���c�j�� ��(��0���;anMћ+k[�~�t��UZ��cH*/�D��c�͍��ٙ�����������AD[{�������K#9��[R8��b�*1\a�;>7�Ϝ�L��ɝݴ%iw,--�w�y��x�����	�[2��S���69���w��u8� ��M�%�P��5 �b�dW��k��=�l�Esn&�E$	3p�8(����4�:�ϲR�yYQ*�*1�ˌ4�)Ҳ�m��Vz��Ɇ_�T�	�[(Z$�i^���Lz��;S 
v�LQ$ʦi��R.~�A֓���FC�tӼ�oir�"���*1���V�s���	Ƙ<O��z�E��U�YX�\A��bz9K��-�;�\�2g�\�1��81t���+5�|?C���������~GU��{���a��^z��3VI���+���d�W��ezar�R+�84����<@�]����믧�Gt��������-��(�LO����y�Sh�Y*[��6}��>E�p⨺��8�����
y�k�A�l��*W��\V���x��G8�cq�w[���qH�N��Wi�l3����fL��:8K6�0�ґ���9�e�O��J;b�3��#�E��§\Hr�:	�5����)Q#N��E̊o�`+��oz\nT�PdBa�U�"�xj������k���b��A.o8���PX^��s���w����������n��w�p6��.U�5u�}���Vc�y��]���^��L�[�c��Wf[����;�$y��Wgi�i��Z�[�e��g��_8��`�s�0-<U^3�ֻ�������x�;��o���?��G6V����{�3�����j� 0��=ӊ]�g��##�Ga4�WLn+j+J����X�bY��4 E�A]2���Ŵ���F��¶t#��:����W��5�x���K���q�~���m]�r����C�����/Y��(����Go�	��3��L�ЙvLV2�#2|�B�����{mx���fu5�0A���9G������*��b۰2�m;UĖ��=��&��<Z.��{=q�$�	��)f�`��a\.r�}��]������kV�r��i�h�D�Za������(V���{�o����mVpGyJ���WŞ9gecji��Z<ylzÿ�+׆[��syl�U�b=�bY?��?���U^ky�ǜ�}Dm�1��m�tP�-�����}��8�Nq�mH6����g������ךU��5C�!�
��(]^�@)��t�&E즯���s�l9>��.<*6h��{677���h��r9�=�ģ�V�Z��N��P�x���3/�\XX �jcy��7��ԉ���,;)��:�cc�iIf�]�l��l��Ѳ��z�O5�#zk���y{�3>�5���� �
��n��$Iʛ�J)S�){L%"��ie=�yxV�� ��_�÷1<��YՆ*O�.�^cV?�9+�=G��.X%� q�����4͙6 7\��sH>�nLwӦ;�k�.k�Z\\Z�]��	=�)3� �F�+CU3+&(�e�B�^x���^����ѣ�h��nx�(;V��.�՟�����f�LƩ�S��ȯ���0N��T6���ΆB��{��aok��k��Z<�p�g���R���S1/�vA���z�M�.֕%�G�U�K$��ߎ�J|�m[e/��0:t���� .��G@̷v3-�T8��(ˇ�c3$tf�-BŰ7�lNuI'L5�m�L�@@�eq�r�!`�U�#E���Ta0%�����u^�h|®U%�
���c�,�;�+:�|�K��Vy�w�}�	�*�p����s�M���V�n�<���w*�3����0�m�'�a|�O������g�Ƿ�ٽ���~n�,xc�^S�kN�,߆�lL�M^[v�Sr�^�y����R��<�����T9Q�2�N�rIIul�]�b����/e?\۪����V�\K�� ���uuerb�{�\��q\x>sp5;���	W~�=�yO����/��Y?����Z~���S��}���[ǎ]t�Enj�|���!��*�g\�Gm�v�,���|�dHyN:ʎ�j����wX�"5��������)�I��qj��T���c�I_�P&�ɉ"ȇU��h(R��|0d�7$෾��n�����X*�*��%�5�o���`ii	�Y�
p������`L�UQB��7q���M�9�~���������z�������_����׼�5a�t���I��4�N�CP���	�V�ŐH@�
g��`SԖ����^�	!CLz�]p�����?�s?י��e/{���}�=�\y�����O���K7yի^��?��K_��4V��A�!�멨�2���7|�y!�M�a�3�sT�y�m^\�X��e���_�{I�c��0�&�+��!��~�ΛN�͂�ᇅ�),�������&*8�D�[�a����Ndt8�υ�8���H�3��9.��I,��vٷd�����l�-����V�ɺ��g?�~9r�����+E���D�-n��E_^Y*��W�Y�5�`#����
v��l�-�@L�L��$E箻�b�JO�e�ǌKܪyK�T���!|�j-젴�0�	�G�4%�z�ERz��ϣw������Ǿ�w�w/~�766��� ��+#���l����� `Q�m�E��~����"�tkk�������o�N<;���=�f�2�܆�hDK��pIA��@��!X�h�A7�R��>���I]�2��m�5.g���3�<������4�y������nL�h�����.h�c�o���=�Ϡ�y�UO���2βCn�a,ʊkY�9�qd��@�ƀv:��&��<˲�`Y��$����5���P(t�U�j��+�84�ˮQ�����z=(�rO��V��c��c"/+�\jm�qP4��dˀ,��w�Y�n)�ĲH��Pq�x�T�dm4��O;Qj.�\�i,؎��K�L��Wj�!T!���u����zH��#���v�����<��0LpsH�=�K&1�冤m�#`oS�Jr�zL��w'\���}�w����~}�AZ�帢c�e��Wv̌|��0�y���(P��I�� ք�q����g�yN�8�R��z®�8�mL��S[xV<��<�2�٥Ou�^��O�ݕ�`-��ؓ���X�1���SX���{��DBI�u���2�)n#.�YU[��z\MQ���.��luM0ck��v�N{l�q��
Ji��P�D0	Gc�:�	K�"ODf�e�0G%gI�ƅ�r��^Ȅy�	�f�����C��ʯ�jӅ���6	qVcK.G����;~r��W\�����tLA�,���^���ZQ��I���|�K_��'��m�������?�󫷩������)\߇ˠ0�q�T����)p��cB�;t��^Ǚ\���C�~�M?�t� [@i�����O~��QHQ���%NI�3�pX)�ETJ�s�ȑۿ�������q?���;��>�ɫ������@�-z�u׼���ɷ��]����3T(ڤ���[����3��)?HHI��=�yυհ�j��r�=盱|���r\��G�(�;~H�z읱�U��
��#��H�1b�4�c@�����-�=�o�dT���i�l�s��Tb��)�\U���3�nsDJ���Xn>��B�zjqDY�ѕ��T*Oe^�z�58��p���V!�9��3���'s0�D�q�3v�W��W�_V�a�%/��.�KhFる�˱����*��Z1�l��7@���<n������ۨq��D[%s2R �.<�s�aIu��	��7��g?�ԩ#ǎ\s�5��y���g��a�Ð������e���ڊ�(�V�K
D�+��H�=~�A�Q\�s�;�ib�rܑW�g�Sټs	l䦈��'�8Q6=���t��{�7Si�vJ߇f�2�#���h6`g1��+���D����1�y� �q��i8�Q�?�Vq��o�n��Jb�t�u�kU��-X۪53��SYՎ��%g�yA"�Gf�\�Y���mfl�^�\��>�k�.]4J�o;�N� IF�ӥ;C*�/}bVd���8`�;�`�,,�x>���(��BtQZ��Q�L����"�d�*C= U�"�!�(>�����@���Ӎf��8([�=�8+�-���<Xf�{+r�Y����Np�]���Q��<��Ĭ�Pqםn3�K�)���*^.k؜L�U�H-���Ѩ���f� [���<�$	��1nS��m'NY����f�2���|_M�KP�^��x �ܭɧ�����0K���-�
���w������-�q���Q �Y '��-��(��z1al�1�����j��~o��w�w�ϻ������>7�+��N�<�5X'�i3Z�Hq��\"�M^E�KF�?p�f%0X�fLR�̗t��x�ަ�R�,��U�@ܖ1�eWf�ڒ¶D�\�]��%pQs�X+ mZ[�Ǟ��/��\��D*lF\���=N|�7��R����V�ӥ��r�������Ç[_��̚K��}�P������y����][�&�v�	|(2�[�H33�8���?\�@��\,�L*㝶�v�#��֒�P�ׂ��ӎ�Q�\��F(>JpU�/��;~I'��|��_���~�/������*K)�l1Y��@6:t�^^~�問�@�
I������Zr�7��b�>foc�5	�]c:���|�+���w�T�FS��y��n�"�r�Ғ����*^b�#5��4�*�⼁����k���Y9�O�'.�����YYYy��_..�����������x��^ך*^�QE�~�7��y�S�5����뮻����_��_��7�2|3LK8UI�K���I��k)�y��\�z�
ZI��A8�L��O�uoX?��m���	q���ĵ3M�ޫ��WyG�Ҥ�X�b5��Ƭ7����� ,l�K���M4�s����*�Reׂ�Q��$�E��T��RF��a���/��Y�o�#c%�mI�`ߣ�e�l[��K]�6�B��F̷�+�@���#ǷE�+k�\OO�d�ٔ��կ~u}}��/{ֳ��Zo{��>��\z�W_}��>�)(F�����(���q��Fﯭo�E�gj�>�!�����!�bd�5�
6T�\�kX���V�d��B�z����>�����z�� p�D�)roR�Aߒr�Q�� ����Ϙ�4˱y�U�.�a�$KǄ�B���DT�yQ%U���/Qu�!X��5;;{�E]x��Mד>)�qs~~��sRW7�Hw\���={.��xi�%������~ ܅������z�e��=����DpL�s��� ����mrp�;�3E���i>�G9�zL����k�sAe������ڿibG���t�OȀ���.�*X���o���Y���hyyٍ�T�2mT_xR˪W�[���Wd<����R��@��3V�䯕��m����)x~� a���j��m�'��Ș��BA�D�<x�6�+Z0�*hp�M�����OY�� �}L*ic�Ml3�S�0��T���9�s��U~��@@A3l>Dlfv  ��IDAT@����(I��c-9F%�S3��k߃��1\�/�}l-��<S�� s�:�ٳO/�Y���t�S�N!� 5�k.X܃ukt�ף�������Q��ݱk)4��덯�S+��9��C��v�ck�;��jK^f,1];�M����O���|�#Ӳ��`얩O���6)�&�]+��y�?|����7���/���+I'�J���UX�Z���k�����y��V�]�"En�P�����y9���Y^ �e 1���^��D(�N���[�����=�أ��7��g>�'!9�#ʂ���6��E�t��6-��UE�-Lkt��k���}��}�{_��W�X����۱�������ʘ����#+�	8�;M���_��̾�E/1HQtڭ׼ꕿ����ӟ��+~�E�[�l��]�i�9�	���t���֏��~��?O���o��Ҋ~�o����(����w<��W:�tE�k$K>�u�W�R]��'�Eg p4`�ãv�W���e[�?�y:�z�9�M.�\%�k�m�@�N<���?�����4�Ă�G4��Ðc`">�6����c>�X��d�q��&�D��>K���4G�|q_p��9+d'֖��zw�޽���(��7ng�a]b�/�5l�Uu6�d.{���>t�ń�4m{!�%��fIK���1�t˟��J�u�|���l#��#T��%4EI�~������iK���]��j��b�S�c�>0X�0�<иK�����w�~���v���{m���S�k��u��H[n9��<uu� 8- �����O��.������L�	�שsT�Iy��-����L�̎Cz��N`����Sȩf�*�yd�v4�v���U�B�:��(1Iac�3�&�Q�sdճ �c�٦�H��ļ��3��+ǎ��J(�$
pg����YP)��4^iV�Y�����B�M��k&Y����8|�����.���k�9|�(I�;��_�d@����0\��6	��Q����E��a
��:I��nB��4͘�Ғ��[U�?Ť�h�X�b��mU%.�[����`��bԁ ÷b@lx�*2	��O������Y�����f���Ѵjs]"��e�a���Iz��2M�iY���#Uw+��Q�� <���]�I �l$�`u+��խ,1>�Ȑ�[$�
���2�0��M�4�A���R�I����&��r_8�U�<�����k!�����n�m9CK� T�u�$6I:e�X�I{C����<��r�j��ă��n�N	x������,8z��׾����;��W?�@�����ʉ��ep�Q����2H�\�i�P����]΅'=�lU�Y2wt��p;x�B�'u.���q�vU�;��r���7і2�lo�{�����y]�fFJe8v��E�FV0g���%ߌ���&H�<y�V�۹��v���zG�5�c.-f����F���:ut+��#Ж�jgQ.���'"'OT����f��aK�1;��;m�=����Z�hE����~X��RcMBۢ�q�(��`p����?��?x��~��~����7�F�����j�mD���c�,+W 	0)!�XiF_��Z���Qq#0ƣ�ˋ_�bRSn������>��O~�o~��^�e������M��m����dEM"+��A�P�k;C�c�M��G����9�:R�i���Ε���v���<�&�A.�̻�����n*�3)R[ )���G���q��z�?���R|F��T��XaeL�%�:�ʪ���N��B��0�@�E�p��U�|�8�1�ɓ'%Te�9�=�����z��d�nI�)�� e�U)1|��Q�D���$�E��k��i%������⋛���֖�n�z�w�q��4�]�veIz��I9��.8S��:��^�䳌QYm���_u��Y̎�Xc��a�jӱ��@�7����޿�u͕d�a�[>Asqjqz���U9�:?D"��=����9r���eZ]7\������^�;x��׿����/�H0�*�_�	�eeu.��o�g����'F�@@@cr1�s0�5q�F���F���I~���^���7rՠqF�2HC7M7M5g����w��w���F�͟�<�6my��>�����]�Z�Z^��\�,�3���3@��fI0vEwcNmw�1h4�p����8\1�l,iį&``��q|||yy����9*�r�M�~LcΙ	�>!IÎ��c=�����济�P0���bN�=��Z��U�
,{�i憙PL�/MMM��? z�U�977�gϞ�h�MD.�;��Gڛgff��o��ܳ�IOz�(�ѕitFKcB�OCSqʎͩ�EYxM�Z�=��J
���<U���L��"&#tYGT�upJ��Zˈ} ��^�.����u�Q÷0���3�47m�d���>H��e׶�ԡ���Ͱ��l�G��J2�ٰ�[g�v]�c#e@�����X]�iZ�3E��d�By�O�����,�FE~{d�w:���@=���ݮ����QL(�e!\z�lz�pVj]Ԏ�T�{��뮣[m�^x�oC;�}zqO2�ѳ��OחXk�l<�[U�<�� �	ǉ�U%~.?,rX�b"Kȟ-�$aE�2�Q�+Wf�kM}�`1�tIi��Q����⻤J!���iԕR�6G��8�ӄV�plqt�����\0?;KW����6���E���6�w��5?:�*s��>�,s�]U��U��[�r�2��hRe��]�!\?֏p<谖m�|��O|�������폯�l'�}'�$��<��8¾bRO�V��x�F��$4��,e������}�#����|�������j��axQ���VP���# Z�Ɍ����?�ClO\���:K˰Q-�ɠ�N��d�����Îy�����b�����'l�擟��q���x�S~5�4�[���C�)r���9�(|G'T䬣;��;�����+.:˦I�q7կ�(� �hƀ��� Β����.K��at��k>o1�-'��|k�z��K;w���[o~�c�w
����Nn��w��r� �^p�9����~����ԡE��;�%t�ZJs�'�0�z�݁�Y�>j�v�l�<*��%	�8�TWk �jN@�����tC㳂-se��tn5��\�ŮJ�0�Ǵ[`��:��%���k���	ԋG ;u�Y���R��
n%a[�`��H�������U:�I�7k��u������᏶N��L�o��w��?~�9yk/^,p>�D��e��I_sD���K��6&�C�S�1�e�3,0f|~��&����Ţg{:*7r<�@f��灪&S�h�X���`�'k�������F�2�
6>[�nC'R���3�[�d/��L5��v�9w�os��s����$��;o��֛n���A�������3�ȋ½�
�x��"u���՜tc�Ka�&J����K��k��$s
y}⯉��	�wH��zf̸��ta%�>�y����r������{�Qv�.G��$�I��,r��6�[r.zEb���w��鲆�?���6"�f~�GY��Hs5�(��i�.����|�[ͯ,�碸�gxlM��̊ܳ	O��F82>2�at���c�1'��mmZ�B�^�{K��46Odٱ�L:��,E=Ϸ�Q��r=q��t�����,H6���Em��X�"E��S� ����U��2y�R����`=��i0��y��fa$ �����׶�p����H�rV\rh.�.�K9���I�����w�nNM��OM�2+�xa�GI�jT3���<�l�z�:���,Ob�2��0X��3$���m��L(.�	SF�GX��q$�1K-4�e+����s�s%�N�ĻA0����mTvT��E��MK'��D,�̚F�H���c�/��Ĥ��F�B{ZJ+��#�����[޸q�	'�2nsg�`��-%�Ԑ[!W��mǎ�A�r����\x�VZ�I�ƥ�wꡘ��<�b��"Bvn����5-d����h�TX�D�$�Ƃ���9�0��Z,*c��%GN4��v ��WJ�����w�*r�_�h���B�����!�3�����B��IJ�!�p���
�n�O�rRZ�2ܰA#�w��)�4��2h96j�\ =�h�֏�c���ǃkY��ђ�s�N.���}�d��f ����ܳ�:c��L3	�L��������g?��g>�����������2��E j:����y晃At��Xfp�º��ق�p���T^$�dQ�0M�f��������~�+�v����N+ݹ����~�'>񉗿���ڗ��Y!j{���%A4L�\�"dU&T�A$'�λ���� �@y�Up�N��"RO��V�%&������ܱ{�֭�#��� ?�����W��뮻����/���k���v��u�cN�%-�F�ln����۷oڴI~�M�,���9�E�zz���H�����uJ��}�UTۚ�W}t�&VU9g*��nY��+UU��"�)g4�U��4�f���R�Ӥ��O�8�߸q�e��Ȇ1��&���{����n���}�^���q��	�P(�K��^ѥTU�
�2�Z���I+��#�/+Pq9�ĺ#ԏJ7Tc'���tk�g�\�ը2�t,]��d�c�lB
=����A��{c���n��F����X�(ݱc��[w4� �ypi�쉱��0D��m۶���v�ڊ�?H�u��$�`k�����|�8���	�[.�\���u��������ǵ�d��e��:b�
�g\�Kv:22B�-i?Կ2-V�K[������֚a����S��k46����k��'G��i�ZՎ����^3�js\����S'�g� ]�:%�Ъ����GG�O�v㍻���O}j�_���\Ȗfgg7�Cu}n~��H�JL��ztԳ`3Z�Ç399W�kɴ�yXy\c~I�Պߓ�7S��:�����!}�,�n�˙�t{H6,7�l���:��hѠV�Je�7�h�0�Kע&�Hg�ӜZ��!u렏2�Ʃ0�9�����y�a�Β"�3�xM���J��L�ؚCz�O�8�C�6"�#���JCU@Qh�h�B��ѐB�ز�0v���>+��X���M<@���x�^F������e�ܹ@@1#-7�RZ|���<��l�����dRQS�7c%��uei�7t�Q?�;��'��`�oV[#��a�/5`sK��x^��~&#O*����ꋔyqA��,+���J�k��J�!a-S�Y��OdZ�꓊fA�j�
��5z��!�Ɨ�s]�aÆ����i"�ۥֻ��Q�a����0���~���x�a-S�=���s��/���{�w�}�k^o7ڛ�?� � {��ڻI<�ȀL��� �m{� �ꗾ�����/|�O}�I�yv���k�h��C�y!%�lZW5T���O����Ɵ���/�6�˷2�����?@	yZN��d_)��vv������E7���G��i۲���W}��\����S�����|Q�z���Z�dN��<%�c#< Y��%���BDO��D��Yf@w�~�51	�Ȁ$qȱbt;tzz���fY�� h%ly:�or᏿s��{^u�;''7�&�:�`V#��K.�`b»��w���/o�]��O�ڗ�p��g���p�f�v�O;�1��^��WЖGF����[-5�i� �O '���eȤ@B��A�hS% ������[�0���jZ�fQ����]lGT'-�O���̱&e/��������d���;Ƿ�2KD��9e2���{=�|nnn��-�۾?��D�3�q���KQ�Ѷ����E��^��z���;w�|֙g>�W.�=77���.;���!A�3���b�;�����-0f�X��+3�
� ��-B?�2M�y��h4�et�d(�$��� ��F#�$Ȕ"��r
��M��ɾ !;���c{��Lw����fiѧQ�]"��z$̔ݍ��ت� �omv��Ⱥ���o�N��˚�ye�k%����c#���@DƂ��p4l��a�98N�|Y���s����r\srd�{��d�E6��EWm.,����m�/�����W�X���kk>��B�o,M�����`�����t��޺uk�usx&��԰����xV�+:�Cf(�Y�d����b�,��@m;�'0'�0h�c�i���	/�_��-�_�����e{&�'�\�(�ޛ_:����9�92���wv��ܽ�@�2N@d{H̏���|���RE�/<փ�:�������M�+��K#��x��̢�@ЅlV�vHa�k&�_����*?aVa]&֐���Ǥ����p�q|u�`�lg0��S3*6�5�,X�4�W"H�P�e+��@{n)F@��ƴ��ZB�eR������h���QD�L},)�+�� h� e{0y#|^��`�B�6ƌ=�h(��Ω�+ɘA*�Mp1�J�8�4�#*��a��5k��U��JIo�B�C�G �ߋa�^�߰Y�5����md�YIA�#�&EǕ�4ǒ�(��ښ��q�%�V�5���A�K�m��T��H�ĢʃPz�-���`$�2J�W aNIb6F�b��v�L!�Ť�də�f �;��O[I�fQ���?��ж�5{b��FD�*c~��"ÀVH0�9���?�/��j����?4�y�X?�s:�E+Y/��?��_t�E(�"E�\����{L�f9�b�u�,I�T��d��c��ɛ��&Z�x�&�0���2k���q����\Ҏf�6'��x�9��c����2��J�N~啯x��M3Т����4o�q����[��֙����暍6���鹨������O|�^��K.�$��XehE�4�:��X:���g��u�#522�/���,
/��H�g!+�I�$��un�xN���hDgAq;���e/{�+�s�ǵ�P>���G>H7F��S��Tq	]�����������?{��_���_����/���=���җ��}�@M��~�#񶷽��-���0q�JD�ʱ�;(>?j~��u��?JY�J}�h�Ys>g!c3}T۵��Z��2�V2�����W�}��h�`t!�A�.�|��"�t�E����݋!ΰ�8���[\�)�ݻ�ص�Xʇd���P�5|��^}�������x<�d�ީ*�ND�I(7e|Z^���S�j_���r���mp�%�<�r54��cqq5��,/�v�m����;3���nٲ%n�2&�Ds�
}v��mt���.��8^w�8�
��ȍ�*���N�~	3ҁ�n
a-�Kp�L U�R�k�&8k�\=��m�Ν3�#�YZ�ṫ��Ag֐1u7��0Ԥ�יּNu��|<m��N�avꩧ6CdC�}X�cc�bѵ�l�+����b�K�V��SFF�5"F�}��t�w�;�$�8w�馛��L ����MKt��B����;��9餓�s�l�����{�)�@��jW����R+�y,�y$;=<��	�We��X#�jy����-I2	'�0�Y��������Uʬ WF1�9��.���Ұ� �J�{i5wsFt�tgB6q��Ĺɳ�4��YN[I��ψk���Jo*w��_�TF����J�es,"T={=�E�ӏN����D���+S��Z��a`��I{Y���2��ݤm��;�p}��'\m��{J#����29#̥DJ~�*J&�T�\yV�l�1��l�AYuf����J�R�jV�#K�%o"��_�L�ʗs�7fZ��vbn�;��R�|e�q��6�	,�z%�D.�կ�r�0f�\��ޜ���z%ͯ�41��z!��Q�/S�g�����@��*,再?�մ����@K0Ϯz�;��{oVE��'
����ȴ�ю5Hr���E��:���2=3��&Zͬ2a�N�Xf(��h^Z�\ <'}ί_~�_����G7mE �N�Bđ�;�4�5�c*K3�gƱ�q���>�ٯ|�+/z��s٥RJ�-�^p�o�����G����_�ܗsiq\e��������Q���#7{a�t�*��>m�Q�ůṷxkTa���ӆ_@��62��N�z���-<�i��������''=�!�<�ъ+��79H`3���{�3_�gy����?�����w��o����0����4O>�����$+2����W�����Cv7mG�~�llQJw��.:��-G�HRJ[�	#>� ���F^!A��q(��+�a��х`'j\).^�:��?δA�34�qYiJd�-T�bl�8{�Չ���h�hcc�Dﺞ���vza2HZAC[da �3=�<w���� 7�|�w 9T��?7��_ȝ�jx ۢCh��2�V��2;�_�����n�ȊU^lޡ5�kjV��%��=���t�P�4��Y4[��UA@S�={�v��U��	yR��8�N��(�B���Q4�&����n���d1��t�q�Ӎ����{�67lDlp�G��q�R2��_�!�&�i��F���%�BrB~-���cD:e\T�f8�
9f�E�L�[?�eُ��3��[<���b�7s8(#\܏z��l����m��Y=9K>�������L��_���J����R�%>!s� @JiA����=w�� ���,���P�`�Wp�'�������5��QN���w<c#��.F��c���������2�(qwv��ZY�ZX����q����AuW�ݞ�}�c�>����{�Y�ڦ�i�ĸv���
�
#Q�ˈ�(���Е�XA�m���u���dϢ$��/��K��4�uU]�y�"2#�e%&E�^�.��㔑;Jx�	���8��0:&�����p�f.VpqN����]%@�����i�!���"��]�!��� !�A��֗�f��Mi�EG̷�,����*R���K���ZVt0�B�����~�1� "��{��R�����5�*��Y\�*c�A�ԡ�
t̰1��W�F�:ADqF��劶m�H���[�kvFh�)vpDq�fQ7b�w�F�� �STJ�%t�Jǅ�V��I!o�S��]���^c)�����l�D�Q�5�JO����E�~
�*����L*������@z�9�����������n�)��aڼ<���Ca�D�T'��^��P�8t�v���PH�C@9��
̕L9�UHi�p�����~<��A��W��5�=�y���=͆��L˷����Â���z�s�����t1�m�� ��.��v�̸0�DC�
v�	Ӳ�*=�X�-�AJd��կ~��>�����W	/�����/~��w����AB{/��Hq�/~�|��iэh�(�y�~�B0K������/>���ʗ��dQ�|p�޹sg����{�)��I��m��F������r�/X��ѿ�����W�B�IA
�&]D!,]e����� 휢��$iࡘr/��oԊS��ؠ�`��9�����}l/�"�+�Η$������,�>.��E/C��a��w����}/�	� p��I�랶�����\q�vFF���7�#7�vK��YGH>�������T
�'&&�l�6==-nf���!.RɎXZZB���"v/��{~~Y+��{U��jT�����ժ��w��v�C=��IbaY'Q��J*By�Y[��0L�ԍ#�a4!��cN�QI�r�)�K�g]��A�~~��: Q�٠d��CǦf$��@AO0$#c��WH{�)��#̜��5�����܍NDB�0M`	uS������ꑆ4��R�
�[���\�Xڊ9��mx�C��]�5ÿsCͫ�~�mA�`8f�,gp�K�$��}��W�1*(M�#X5���Ds>^�\������=p�SSS�G��,``���iz�ѢE�3�B�oڴIq�]��ݻ1�e���ss}��!����3�L�����C(��2kꙢ��H�C!��,К��$�`���L&�p��ł�Si�N���P�Z���W��WE�2��n�(�t��x����h�Rx��5Y�_"	��Yi��Md�T����3\�a�D�uԌ���Zg	_!�jf���s�5���"x(>/FI���Y�Ƙ����EE�ԄR��B�� C/���텁4/sA\��n�]��m��6�*��"NI�-Y~���k��f�t�D�V�,Xġ"{�3H�Y+^͸kIr�����l�Y<�I�^&`*�Za�����.B�S�2�E�_[�$�TE��b�k�X?���Z�{sC+�l�o+d������&평�>I��dʣ��\��Y�	hI�T8i�V�96]3��bEx�׏�����4K��C�����;�㮼�ʯ~��oz��B�V��w'���p!��Ү�l$m/B���fd�p�'�kR��R<606�ad2�g�{K���6ZEVh!|X�ڸ�r6pWF�؃<�\ߏXNu��1�L�A��>t'���*L����,u��T�{�����v,O�Qrj�M9����I��������������-'/T��������[HuJݢ+�vX@b��E='lGȕ���j�q��[[9qN���r%��(U*
:���)<׈R-�G� #n\n��I�%��@|�?��rnC|�B���gv��6+�q'�ĊU���/$��c6���j҅�<�]嶚g=��G�s��`qnvv�,N2'��^��pF��B��X�T&FB|W��L�Զ�x�,�ZW�$��x��ZT��]�9Y�����Ʃ��D|�������D��5�	R�<`M�6,r�E$u
ԑ�]q�PY#������&�_�g�=����r���]������f4��z�s��FFl�vbGq�p�p����;јe� mo��$�~��A���ſa0����*��M�f�*穇wbi�phXK��s�Z*[^���hf��ws�Z�i-	sd��=bEi����Y���̵��M�ϱ
կ�G=S�e��*��u|té��C�j!Sn���!l*��~��A-���T����tZK�Mغ������G�-,-��.�Q	]p�Ӟ��"CX��=���w��LNN^�GSo��8j��\}5ac7Kӹ�q�sf0�Tƴ6XP�%؅C΃af��+V���Z�B�$���Q�e �����8J�hT��V�[��2�@�X��ܶ��
��[�aa�����yW��*�����L�h�A^?e�c�]�LP� ��m	�o�S��uxA���q���RA�L���V��!*����2!S�lذa~n���J�YV��m�qB������Ǵ)@������5!�9V\4�ȕA�#WL���
�� ��~(�s[u)lS�c�iIW+��i#thԅ�Fga#\XZ><5w�C2�����O7�:��ȩ]�Υµ)%(��+�SQ�ҀI��}+�+��`��~�J��jОKmb������e��q��ލ$DA���dF:g�	������37��F]?ad�\+�R/�Gř;y/P�M�ў�^�Pt����,��*Q.�+nF��:|G���J���[�Jk�X?֏|<����!E@+Z8E��r���s�Ti��UȆ�'�(�b�Q����h��Qc�\���i4�R�p�B��XK|������}�3�y�������.2v��%k����_�Y��w<�
2�<��m��� ��ig�C����6���������g��Y����  eWY7����*u���<�LW 4�Bp\�ȍ�xh���;G���~�[�M��͐\P����hb��!Fh��VE��a���9PA��2�m�SJ�e���d��E�&�,u�&�+d6��I�~��O�ڎ���K�dMw�V�Zk��ڮ��5�����5�١�t�UYv�6f�Z�t7���V�E-Ɓ��򂌤�2�)�b��ґ�b%_�~?��9�X�T��G��儼�8�+�r���2]��c�{�ʎ�
�����i�y�zdd�3�g�(�c���s�cX��e�C��[Jh7�$ %2��4�"jV]��/�ؔqC5Qy�51B-�h���*��P�(�S#�:~�4��,ˢ��񳦵h���*�C����B��e7��<
2������_�|�B�
�8����}��x<NlZXX(X2ά�U�F��Ȝ���n�x����n��>NS�:w�=��~ff�*�9�C�X�n��e`];L��a\I��v-Y�i�՜�N����u��h�"�e0(��R}([Ѳ�?�-5�R3�Ъ��$+�Is�(KI	�R��>�%d����I�Xجe���(�! m�4�V�?+)�(�� 4o%�8/hx7'}�����c���w@i�F:�Uv��f�A�V�Z�h��nO��j���u/ׯ��8a݀V��g��$�8tW�7o����KN]4L�YI��-c��������W�bR�Ck&����ܕf�XUy_5�oU\�A�<E	�U����3B��Y��ZP�O�\X�?�Q�m쏪���%��Z���K���&⎍�֢s�4#�+z�����]�	t���c�X?���O���5���Ӆ���{�J�� tPأE�r��4��o׽�hq���	��Y��4�6�*�劖~�Ю�b����[�V\�"0�h	FX"!2�ݦ��ç>���r�+^��&7���_n���8��Ɩ�����p�'g��v5��Ei��3+�(�t��:v�-94�"��hqΐѠ��B�0$͖�-ªP�M�|�B��N�I�]r�h�#�A�B�E
�F(dyʲ���i��+�	n�)�zȰ�DaB����T@�}{aS#a*�m�w�>�����v[�䲜�:����M�+j�dr�,��*�wu'ӓ8.g�L�r-����F'�q�]���SbR�C+����M�uQW����u$�5�8Ɩ�]�p̌��ڙ\��`�0�!�4NcO�aK�I�O�g�����}��l�9\ўc{��";�D&�L+O:N`g*����J}�u}]'������!���֑X���)Y7�T�n �N�Y`�6�fq;r��le�s����Zn�V4����X�4[���i�2���ǩߞ@����aK?�t��������K)U^�s�E�����젻o߾}�z�R�.��R'p���{x������FZ'n�~�#�!;�{��htvV5��۷�o�������}��^�ɬ����э3���l���G�5::5�O|��:�������CI9������g�i�l��կ~u����!�^qP!�q�}ظ����"J�n^^�����D�ck-��*X.g�J���D-�O^bŉ)t4�������hfnayq��NԆ��ލ��F�,�آ�e�̀��2��q��w�l6��8���
�	��Z���n�d���2�p?���O�|����/������Pk�x�C��h�;;5������3�|�igܺ����y�O7J-�z�؈`�hU�PfZ@4/e9�ҳ�ܲUFhr�e9Vr��X���m����b̖3y�2G��=.Mf��xnz�	��Ѥf�́���YW���c���ݖk�&�㚊�V;gG��IK�!��[�^�8H���+Wl�;�=�F�M
TSdXEN��ГpE��l'Q��`��!��/~J	�b�!j;=?��0hJ������i����"���<�˶?8���~gQ��ɀ�!�{�b�$(b\�g�fA$�Ѭ�ћ��L�q�cc��5�z(E�E���D�z��cj<�|��;�`.�����6m�v�)'<��aza���l�0Ō��k2ZU�0tI�q"�CN��ҢڊL5��*F�s�EIFɒ�����NW�0+��sP��[U�K=�AX���B�T�ߜ�\9���c�����갩�����?���kHZ>�o߆�h�h~�����9��g*;�gҝ��ٲeK�C:Y%�����e'��˜*�\*-� ���E�|_��R�O��O!s�V�F����~��?��c��@A��G؍�B
����!p-���ns,�.�����o<Nn��C��'�lI�t~��I������E��MK|;m$^x���,��w�_��A0��P��B��%B��'�a?�%��,@��~��k�C��GzQ/��0 @��8ʋi���6?]5[����	�C�b�n�bKg��
���Z�n�ūye��(�:V��АAa%O��R��g���4|��T~���D"�5�/��X/G�٘�iKo4Zd�d(@������C��7k�*�^�Z�h�*j0�D�L�G�]�d��������2�jo�D�S57"�b�3�DR\�7?�v���ϧv�WN��&�%�nk���Pk8���o�i1*3sl������b�	��z����O�ѵs�4MZ㧜rJЂ�f�l���^���<䬳΢3���}���XgӦM[�;���ג�~r��j���w胄���G�g�M��qD���m'N�pSSS;��O?��V�\���N�\�e�$$=��(�Ky�#RЏݢ�y5lPCT���<*�"���S�)v<��?��ZNPW]�H6�1�)~tx���n^B�1��F��R(�g���@���klY�zt�]�v|�����PD��Q�]Q�I0B�T�JN�����p͋�>��V�:�b���͒CI�L~I
�TGZ��ŕs�yy��MUgI�#c�^��;rfȷ���x;�Ye�U����w�LdBā�GZlp���	s �М����8�"r7n����/--I^%��XgP���UBrR�@ᐫ?�zH�<iqk�s��^�w�]�h�!cO�����J�U�U��gq��⒀t�x�YAx��2l�e�K1��g��`��3"m4+Qm���V%�2�x���j&]c�H��H�׽z^�輠h*	y�|(jdI(eB�l�wrrr۶m�;�,;yU�7�WP�ͻ��2h�q�X?֏��:�E�J�к2��i$p����Đ��O{��F��������(�Zif�[ǁ���E��톍N���J�r��Dy�b,��Ts����1=�ba ��q-��������^���2M7����6�����d|�d�M�˰���6���n����9��G�e!�n>����5M�'�yg�|eף�;�"��1j��k ���͒�(^�U�A��a�[3�ܓ�B�H���2U��4�l1
��,���9<�6~H�Tx��~�����=�f�����Tmiώn��;ÖD�AHj��Y$�f�=V^.`f�����=�&f樹��Ba���5-eP(TA�[�P��Fu]C��2?�D�dI�E�mh�9�+�DZ���������)g��6W�a��5j+�-!�$=oغ�FrfV40�kTj]G�u�R��oPe`*s5��߁0�����<�ޑOsD:#��϶�ȉ��}xv����C���Ǎ=��U�����o����9�3�?�g��+�u��k�髇���W�yƩ?�����'n����=m������w����bh	�$,{��D�������?~�ʾp�7�pb{��QD������믟��z��qOt�&���x)"�-�t�0t��r�č�F��K	�h�-a��A����~,��®�Y14�4I�������jw4B��A�dc5h������p&L` k�#��rPcY;����6oێi��Ǌ�$��D}��fHX`)K	mh���DE�v�9:m���[7n�z��{ﵲllÆ,O�':�ԃ�>����;�;v�{�J�P��cP��]��L�C�{?QV}��we�?>�J��W�B�7���v��
9�>a�>���� �Qa�
�+Hj�8ʲQ�:aM�^܇!"4:�Hc�	VO+zyi�,�!��7�$�� 
f��ŞT��3ץ��o].Z��]�dN��eK��hYC��|�G�'d��������V*��2�����K��B�����\IK @�w�!�mhXsOWэ�wk�2���ʹ���U��t�F���GA#��,,,4c'Y�o9cl��'�8����[������,b���>@`�k�o�/l�$m4�.�b_:��QDW��0!�d�-���83�ȴ2U���V����^��֌RUɾ� ��{š�\��-��8A�%�Q��6!�^�>;�K��ϊ����o?ett������o�ؿ+h��M0븡e�W��t'\��Z	}��g�X?֏p<���huR�N����r(;*��r�H���$r��TZ@#�q���q��(�C�5�s�4I����9'���8(+��Y��n�oӚ�"�ت�f8]9�9���R J�7��F�x?]�xC�B��TY��M��5m�yb���O���Qኌ�.������ ��o�ɦ[%���'aH{����=/p�G���d�^�r���r�P��&J�T�z��¯��] =B
���,�\�M����i���P���݇����,4'>Z��%0��_\n�E
YV�:�e���a�����g�O�8��N��5��>Uz4y�'''���eT���j!�( b6�:̾��޾}�\1ͪ|�����8[ͱ�j��w�v���j;F�YG��z���}�?�b�j�D���vJG>'i@H�t8ɐ�~����dg�(ٻwowj��N�69��iS�y����&섐��;!X���śo����?{�sN�@r���1V�tnn�B)y$�y���3h�s�#Hq���M2�h`[�s�]v�fYӌ��a�9ǂ�0�87�
����Z�p��P���b嬿B�(:rE5��I�.Ǉ�����R��G3 4E�v��ֆ&!X� �t���Bxޖ-[��޳z�t����D9��*�0|���bjZk�v�ʭm���C�9�u��46e���3����k���j���,p����q�j��i$��e�������18k')Y^l*ۼє���e�u��	��m�f_�ͅ	t��Y������'���B��!���R�P�%�^�e�V-�aU��>�GT'�_��7(����acUL�L@����t��ޖ��i��8P�귃����݊8�J\�QVlɑ����M]�=r�Y������]uS�]X�IJ�p���h���Ь�^�S�J|g4�d�	�%�C]&[�Rs-����E��VE����̻uvk�X?���Z��g�z��
đ�I�I���4��ˡM4�Ȇh��!�Z9���X
UF���J�b�r��	8���N+b_��+�Ѳ.6�tx����~�m�f���4-mfi�A�Hh�I~��,Ѷ2KcF���F����C[�&ΐ����6��G���d�*��4BJ����$a=�hO��8���"k���;IF�h9*��di������
�a��i�
I��L��f'�91�lV��}�����E������@s 	��X��q�5DtMT�2��*S �xe�ж��w�2�C�{�k%�H�_��pf����R(َ�����K�=?�Wm޼��q��/��؄n�kj �r�q�=���et��(EI�8��|�=(;[ }yܒ&�
cvib(�]�Fx,��)-6N�*�qmX�*�%���ЬF>b0j���Z�+�Te�u%�GU�m��U�t�3}��Nq�)�y�Ī��Ә�?������^���߶��M�[O9�t���sw�<��������gPQ�������[��ؽ��M��4��phz��@g���C:J'&&Z�M��`�dr�FV0�����M�_��K�;4����g�O�~��^�z��~��<*,���u�����`~�A��2G�c\f�w�9����p��$+�-�$ٗ5�J�Kx0�
���.�
��=�$Z�2��|Ϋ��N�;ȗ+\�F��g��h�{����A��&�E���9��h(�xZEE�B�G����F<�&s|n�91q���BT�>�-4�ܹ�5�)�6m���}�Ç[Hm��ӳ-�CJ݋�:>�>��?�22}X�@r��̘�I�9��Ѵn6��d�B�iVDqJ3��n�t�H���H�:N��
��&VD��[����j�o/kى��D����  �U%���s�J�t���	��Y���	د����]TMW��7��Y�a��D��RyVXIݘ�˗!&��豔-́?�������Y[O�0�d���T�������Y JY�.Y�)�4c�-�4�tڴ��r
]�|m�!�)�g��A�]�LOOG��C��1�I���G��^s�I��=�cۃQ�����,-�}�H/k��Ǽ����5C�2]%�U���@�|T�b�oN�RY�b�XN�����A(�)?C�geԷ4����B�kwF�,u�
�Ґ�c|��v�w���o��5f�w��A�Zo��$��ʬ-�JV�e��0�d>��Yf=_k�X?�u<��W����O}��+_�8JB7�}γ�!~��o�ꪫ��G�#��.�H��g=�Y_���������/���?/k?��>�8��ʵ,���+��ů;�j�!���O���G�pp��^�����ө|0�5;,9����O{�?���i��;g�a(��!Pw��=g_|���,x����ݻ�[FY/���>������MR��6��k�]/���/|��I�x�?����ǟ�Ѻ�{n�*�sT�6=�������+^�#q��4���!���W�~��>�Y��H��4�����#��<JА)��G<�|��j�����~����@�ᑕe�Q�^�F��.��/}���ȇ?��O~��tl(��O}GT
�n��*�����l����W��������[Ysd",..�^bX�Xd4l�M7��z=�kwjzff��$���P�&�TT�L��u�v�t6��y�|R��V^K#�����������g�gL!T�5���(��N�C�sii�����A�g��׹������0���M"kcrrRR�ԩc������A��)����>��l߾��s�y���Q�ʩ�Y��u�VBq��s��!�������%:u	�;��Da���?K������-C�rK�d4�!���/E��6�E�mH�����J�<��#�1I��s6o�@BL{@�o$���P��5U-���Og"M.Ə;���~��ǝB�v�iE�۝Ea۶m### �x����Y\D<'g(I��^	m���X3b���[�3�Z -_���T��	�G/D3��~�K:�XqiH����Mi��/I���*�+X���20��>1�KH!�?Wd
�J�N*h����{eH�*d~�.	Egz�Ȳ��ҧe���d�;eU_����ș%��9Z�iE�#ֲ���P1+�Ío��J�s}���߿��t�]4�}�"!H'�FL��c�x؆���!Ϙ\,�&��U�P�(����w�#H9U���W��͖ٶ�YD�"�h7X32��c\�?�$�,��������I'����M�븓N��\\&S�c�eG�i�5x݉V��X����~<��A��ʬ�G֚�ђ�eWg���EQ���;w�������1]Z3� �؇?�_�����a����rw��_�-go{�#lFK2��h�T�_���y��]B3��{���k��������m����QYn6�t�S�=;K#)�� V�5G�a�p�e�bq��];��w^�G���(1v��Fq|�	'�ޟ��[���I�I� |���st
E
�e-"Nq��%������2��Ԇ�,j�8L+���'q�{�F���N��N{Q�[���O��w�`�e}s�/~>�y�׿���{Q��'��n���E���9nD���8�#�����/~���~���w�	��k�K���Vd���~>H���jI���� �R���]��HQN80Z�A��jWq��O�����~(ze]�����\0��o�8.����n�;d�P)6]��f�wXW���(Tl���V�[��^�Ui���{m����֧Y�~ə��WrQ������K�����`�[ �"��Mh;��{ <@�4m{�F�'[�'�׊�;���m���i��6z�$�޶4��h����;ф�n���b��o�.i���4ӾZ�ٜ�12�B�X��Ғ�"7m|b2!���y���7�|����'\��G=���n9|�>�Ӯ]��ݱ{zn��)s�3��#M���<k�-Gۄ�}��&Z>٪���b�ܪ�i�TjaI�7�P��dtK�����5�(�x�2GJ�I�k6�h����2K������<&���h�u�Z-2�Sm���Ic���n��'����X��G.PeA�0�hy#��}d����m�i;���'�_p����b!���i���\;_Z�Ҹ�v荁Αy�B����7�9y��K�D#yT��'��ɇN�G@���"�i���<�I��"
�H�bfi�pa[+���r�^��`(��O �X�>g���z�����+ ����`��g{�nXH̉��z���aq"�P�}o%��º�2u��(%��Q:+���a�8k�qQO�f����Pߟ��.�.�'ZU��v��[��I�m^��g�
��l�U]��v;B@�q}�W�qo<3��}�,/w�Em��e����L�EA����ަw�V@�[�z�>ݤ�B�4�r<K!̪�+�N�P�vum�#��AUU3CU�Q����J���jk�5��Ď�̥���hw�\��3����ƴG:s�(��\\^j6�˃>��- z��f� z����uFX�Ci˴4k�X?֏p<��Vy��H;��>����y��"M� ��Գ.���x�s����<v�}�[�zӛ�D[��W<�s�|%N�P!*�w���������<��}��_�k��������Yf]v�%_��?E�Aބ��-o}��>��w��'�t�s^�"�p��wЯ�:,�i���7o��7���ؠ^�C�۠j���7�p�_��_����\w�y�9���t���w��]�\r�c�<U������g����\�(��b�o�*M�bqE�~DA�A�1�溰��,�����|�3�|�宝@z�8�vs\������5�(z��_�����	�}��M4'ޘ�o����}�}�3��{�����?��?}�{�kxoKbs�gLNn����M�e�zp�S�<�)O��מq����.ST{LeH�߉X�'�&t�q�ӱ�:�	�%/@.J�������"�k8goddd~~~yv�l�1�\<�|��8�\�5׃�͐���n�ZxD�C}��������Yk��qߔ�*C�
\H��`R`Ά�D�.-�J���v!w�e��	7nL���4h�>��OO�4�Z�&EWw:�'�|2A&j����33�VK����z�Q� Dې���s/zu�/���[o�t����M�6�;7�xc�vN8ᄅ���Ҡ޺u�3^B��k�Zi�?H�Կ����kڭfxj'����O���Jn��pO��.�!fϞ=����I'���R�=Up�5o��[˿����̵�^K���m'P?�;��_��_N�t� �j�rF��u�8ר��j����k�f}����W&��؜�S��(�:6S[&}|arD�3��Jͅ��,�.ޕ,]2c^ȹpG`-�o,e9�fd*Cj��=�s���o�-�sQ�,�$9���h��E�P�W�ײV̰.1%(K�L��$K-#�*΄�u��Y����k&�Ъƹh�R�o������#��w��{���\\�F�@Nh8�K�&��f:󌇟µ� �%Sk�@��C�p%�yE	����~g����a����u"c�W�	�Vݣڣ �8�6O�f�����!�6w��J����5MU�nǦm��;�ߵ�&�����������o[�׏���|<��VeO`u���NC�R��!����ϑ�u��n���)��--��$��_����$-hw�&Z����?}�^���\�����Ӟ�d�7���w�K^F�Ʒ����/���O?p@-����/~�5�}�#/zū~�§^�iӘC�������-��Oeq�[qYui9�mmvN��'>q��gc�C
�����o��%�~�W����6� JXt1��L}ɡR����w�4�!��ͦ�ı����Z"MΚ�k%�2a6\���3��I���ih�N��qs������c��G>������t�6������?�L���|�C�뫮��,�8�7�l�~�� ��8֘*@�{��O|�������_�2 D:)�+R���m.��Pp����6P%��2�HO�:Ml����Pq?�����8�۾�0�|���7��/gi����/����l�Y�P�V�H�5�Q���*��Z�l���`�U�e���� ��#&�)��Ђ��X�e�Zm.���*8��;��l��RSPu��6���Q,`�)�e��
��bP�\��
�&M��*_9g$ƅJ�fSO��ۭ`|���ǜy������ן��z����ȕϺ"DP`�.ݶ{ܺ۷��\N���'6jZص{������gn��,�j7�,��,����F�������u6�	�e����ѱ�;ow���ɍ���[7>��,��^�ρ�N:�x��<��r�K_�R�_���0�V�`���en�\�����Y�uq���4֕�b-f��4���ϴP�6��O+���hd�oJ�� (|���Ұec���w�}�����.��5e��ک̸ږ�Sm4-n2HQ�)���ą�[�����}�z�E���7�aö⸿�mذ�N.�|�gX�ή6*���]>l�Zp$���1U:���%Y���ӂ�]M���PTHl�'iN�sD Ƭ��� �{y�B4DMGÎ7�+x����s�0�U��&�L*�h4,A�����eUŌ}�v�߄�(��<�pڨ�h;�y��%�(yn	�DVI�	?�Jk0|�b"��_ZV��"_X�Y]2�W�&�pP߹@�-�\�\��VM�X��5�)�*r֪y�#r��_�[*ˠ�Fz*|��\���� 	�d�ҍ����������A>ݟ̩��͒������X�sK��;��~��a�i۟_��q���Wc����y�b��)yQ���ylH�sA���?<J�) $�y+U���eL��uėj�ս��*�N
Q-T]�R(�������7��Bפ�t��'?���	d�ݻw~~~���cccs�hjjj�o@��^���Qׯ�Ž����LcV6k�X?֏c"�U�؉�K4�����2)zC�j��xZ�?���<x�o}+�ADp%�	�d����l�r��W���/��>�w�7ˤ�\s���������>��qJ�+�#�yic�L�m�6:�U�z��?��w���|�8�5��X�\�k� 2e1�D˥(��*����=��Ͼ�e�q���>������˂#6u�)�å���" ������
*�k��o�b��%ZFi�!��(�Wd���e�V���S��׾������8�ڦu��$N�2��;�e]D8��D'�xֳ��[�{�Oo������F[��,��+��0����5��>U�îz��`��'����KKKg8@r����y�N}4]V�=(Ro��^��U)�!�-�"�&��:Ʀ�h���	��IkXF�+�y��8&�P�_^C�]?�ѳL����!��Ӌ�����'�"8~3���{�w^�����?��.���n�瞽�S��.���j}�����N�2::J0�֟�����y1�ns��\�;��om޼y��-������+|�l�(G���M�w�uW���k�O���e��C������с��(��,q64xP�n0��G�6�o���/��P7Uܩ��c�(�=Y�7:�J���g�M ֡��e���s��B.�uᐭ��5Z�}�\e�:�fD��>}�9���V�ٳ'�5Ǥe���7����ɑҬ���lk5C�D���k�
���I�5�<�%��uu[�z%��9\7ס��J�c1ԃ��r��:x��ђG�]�U�C#�̖M�"�+����ϚV���u���d�*r5��ᴮ�Og~��ȧ�E&��G}m��?#�,!v0���-ff��h(��[���N9e���o8p`��8t��$���Y˗�d�yUm=|3��YT��rg�V���P�vK�r2�"�j�\�23�$������S�}�Q)5<EO��X�����BT*ǜ��G�U�`};�Wg�uα�j:���w�AZ��y7�[�k�qi����cF���~<��ֲ|Sd�Jm��/���Հv���i�{�K�]X�'>�B�,y�s�^Zq.���%T=�(5h��P(V�l�/�������*eَ;��>�gv���l�A�׉*XA�q���,����%Y�e/L�]���X��%QH�_���)��d#�j��׼�j��y�s���F�AˋT1H�0�~<H���,*T5y�i�� ��n)�q[d.��.JgizdD.�� �PI]+�t�,o�6aO�@h˸���'w�����Bې���t��¼�6�M�(�ms����	³�����ɯ>�I�g�k_>�HMc�b��v����? ���rrNxPCR������Y�g�h��/���@�	�Dցߤ�{y���;��QKQ��V�Ar�j�~�Ӧ���u?a�c˶��Vbf�1<��C��%4�U������[��J���/���T�h��sV���\i%5$�lV�iO�'��(aΠ�ǚl�� 2�6�F7�%�Q� ���S�ў�;Mv���F�L���󅅅޿�n���=?��<����A�ݷ��ݿ���~�����?�ajj�	�"�f��]���LL���\D�����;����P�����ۄ�E�%u�o��G33s�_��2u�.��xh���^>fK'���)�Uз:)M(�"ie�����f[�gu��j�#�V���uJAy�{����UA�8��=���˞u�y��q�1��܂�T�0I��.F�{��q�V�۽�j%4��р�%�i!U��Z�{�e�U��}�=7V��[-	�j�%�J���	��%�l^����4���Ͳg���`c{l���$ˀ �I-�:�\u릓���9�
-Z�AϨ��j�:��v������A��1e�UK�;�$�
۲)%Fo����� #-��D;���H���L�/S��4�I�$qQ�dBb� �� ���=�7u��*O+��߂fꯘ}E�9�	{�2�*.��XDo��>2dt(���b��%8���VL�~�-��Xލ��I&t�����:��C��;�U7��m[<?��9!�?fp%8��bLk��h��x. uI�5&kWڼȣ�iZR��bL��Jʇ�.���%Q�-HM�x����-�����2�U�*��Z9 	)��f\o=a�z�m�f��V�����޵��1����3j��8z�_3�j���&���C�c"\X�r�=�E�}���Ǳ�l���Ƣ2
Dw�Ze^�H���s�Df�BDJ�S �����1 �cehX�^G9�.�(�"=�7,�9;W�|��m{�]���	��\.�[������(+�g��9�����b�-���<�e���\����MTI�6�dP�}���O]v�vR_�޽{A��Y��c����*��QTlgxx�סC��vO�Z\oժU�R9&�r8�$ي�N仇�?~|��;����I�ӿ���K/����}��>�����=���w�(������.�(��c9q�b�4���[o��樠�/K���!*���on߾]�����b{-��Bn�1@��~���r���/�a#�eL�q߿\q��h=���W��۩mj�°���������^β;N��^(�D.�щ�Г�_������?�P�X�
'�	R/E�iBsf,g��-������TD]�\x���Z�i.5أ��� &oS�M� �9k%�w���U~���Q��&�`ꉪ��΂���U��!W�ˡ:ݷ�N�2�L/Pڲ�Y�{|��ɐ3�[��p~����{�%�)���)h�Sl҆N�i�ߋ��5�ׯw�h'�D��k8�1|v� �0==��tJ�b��g��:^g��yA�Ӂsp>{&��p```��|��'%�C+(tcᚹ�v�)�(j�D��d����2�ʘ�ά-�l��VV].���7@��� 0nQ7���Fn������U����<��H�r�+�g�y���Q�g�7�*F�aA�Ť5fhh��l|�;O�w��R����X���.�X��Q�Uyl��u��_�Kv���BI�~fA�>d^��V*�щq�b��I%��`x�nU��t⟴L��k���,>���bT!�ً�Dj��?d�7����'��h��%�����dA/������UJ����u#<%�� �;�8}��p24�2�6݅�Κ���#&��q�#IC �Ӿ�ng�L=�*$.l����E�"σ3e��"z�z}w��"�!�'�a�a���B�B3AB�RNfI�$9�0�&8S�&'&&���\sͦM`vu��T�nY����`ZT2��k�i= ~�}�­K�*�IX�'�F�e�
����F�_S|���ɫ�ܖ�xb-�[>&/	�2ZQR��b�h@�W�������g*_{���l9�X��Y��Q\*Z*�@PB���n;���CA��>���=#���z��3F�%��Z�ٳ��������J�ҒudK�]`�3�b�$S�ɮ�_7���˿|�o���k.�$\(jv:�v]����?���;-�	@�!�iDXl�k���I�,R�R�h�����t��:dH���&i�h��ܩ�� /��O�R1��i]�[�jt:E���B�LgaMLd�}+2ǚaN�IhX	̄�D�7��_����T
���u�.�ܨ>�n��[N{�,Tv�MQWV*�T���<[����eީTF�� ��&���.^��{�ާv��N��L#��1�,��hv���cN�\���65�9XD@2���,��N�)҈����0:��M��B�S�l���8�7 R�����K�O�ŗiUV6W�E�R�M���Fj���	{1Y郞�T?f��+�D��T;Dr�*#,X��zEaǃߕc��ik��:'�⃧���-8,���Ԉ����A�X�CVaZa��T�vf�BD�Ǩc���n��xR�&�2Xn[�pV���a�
�g1&n�a)�U���6bA���mφY���o�Ó37��UJK4�n�д�U.x2ן�5���ippp�����ɓ�jקg:���
�G҆���:���#::�"W#��Q�n�E?�b	o�_C�P����r�iA��a�:��ʕ+��߿��h����f���� �M-����QT�0-P{�@�T��&k���d����'_1��RJ��?s(K&����8֎f�-4bc�u�����V�0�z�U{�9x���z��r�,�*SSS���4�%��E��\(��·j� X|�lvA�0����v��u�L���f��E=�X3�2���x�PEc�Ғߚ���c�����F$�4#t	�|�9	��qZ���S�@�%WeJ�NT5�o/3S�ȾF^��2�ٽTj��S�{C�b����D���d�=NQ�6��d���a�K;�h�6KJk5�#ь;{�9�c%Yp��%�K(v(�>ZP
��";$���e�_�穧��r�<��\s�ڵ���p`�����eP�z�j��GX���ф=�����Y�zdd�رc�S���=}��/�p��S)�.,ڗV�����\ᚡ����mnn��c1��IMԧ�!��r�D�͹�F���K=�#�$})ʷ����<��<V_n�m��I{�a-A�,�h�����7��$Q��PD��y�]w����|�?��2��l�2Qǚ�E�����v'���6ɂ;f�.��/�plt�uUj �LK�}i�N��eڠ��}��ȧ�yvG�b%�n��d��l۶mfr�������_�����ȇ?�������a�٧�����7�����u�`��We�,y��hRE3�eb��"63���������_��6 � n�6��ㅩc��J#f'R�w��1W�ef|�Ĵͫ�J�h̾b-#?��AO�o�166���CT��_���kn���zir�;g��
�FbRD8�$�x��:t��Q�OS�'�'������3 �'�A�2m�?�b��Ň�U�'��df���uK!�p��Z�̔C�{w^_�޵�'��P�K�$�S�Q�������.]����O�1���bK�0k9�_4@�C�gs4��6�b�x�)�Ӟ��sucٜ�π
MRF�,��B`��(�ꩠQ�2J��P���dJ�����?OS��l��w�� Y����������jpFEq6:3�S�$�?�(F�p	Hd�WWg� ,v&��3>�.�(��h�Z�E�+k��̰���o|��$3`-��$.�Y��Ӽ��"�鋧�3�*�}UL�� �r�6��pTi����@m�m�^�;��y�'l���
<�Z$��,����2E������9��hJ�~v�i�im�+��/.���A�-_�ϖ�΂���킱��������"˓�+���^�e ~ lV��aD��{_���u��Փ�hY�p&^��,�* �$c<��8 G�ȮX1�y��U�VMOO?��O }]|��}}};w�d?0<��w߽g����\s<�}��w���'N�p'"]�0o����Ͼ�0�6n�p�9� �"K(&Iv��6I�p�A�M���+3�"�:���_���@^�=.B�V%�P��f���d�-�%p���r[n��^~XK��v#�z���X�Bv"�펄.��O����v�����[��[*��?�Ԟg��w�vPm�+�
BtZ�MŨN�<y��n�|~���i��ɞg~����w\iF���r�f'h:&�|�>>����r���c�B��F̥%��w�]���\���L|7H�#C@
?���EJ�����W���|'��S��%b�!d	ǰ}[G%�U�q�-WƊ4�K(���[����h���xT.ç����Q�, ��6m�𭇾��i�в��dQxI��i0���P���.��O�d_�tM77�(!��)�B�� ��@��I-�3~��8L�`c8�{��2V"�n*H���ܘI�8�]0*Pi�f�0A�tmnnV��d�P�����Z���N�%���J텠�a�?\5"�T��&��E��x2��"Pȱvx;E؀|���%1Bz��;o�Tr!�R9͉��UD�Xd~����T��.�J�?v�j��ؠ��.�\҃*C ?#��!������a�ZO��!��\�[�j���Z��HQ�u3jXgNnar�c�����N��δ�	���g�H<-�<,���L�1'N"�.��܊���XKA�B��X�� B�!�vpA	?�Ѳ4�	q���}��O[�����(�GQ&!+���1��0FG�}_��	x$ ��V� 0��)�����p��#�n�ޡȶ;~��:f�	7A��v�v���NY�C�sb<���f�\tT�Jc3��?���M ��M�&:�A)�ѿ"�猢:Tp��XL�-Ӽ�8��4M���l/����"����,0!&�^��r�& ���)x����^z���֭[�: Q�ɏ}����)x���}�> ����LD� �@�����?;�5�][Ȉ���&��`��'y6�]Z	��T��)��S5o1��kڅ�LL��d�͚�UƼyH��=ln P�O{'(�ӓ��?N�˼�*{p����ED*@0"���:J0��K& B�"��5�)-(Vq�+��d�4ln�t�y���yPa1��ǟܿ0ϡ��
s¯֪��Ѭ�l�4��6���_�k�60�P� Zs�v�9r���}���y���O�(;�K.���[n&)��ht���`�#�<r��0��~��l�
(%zvzz��U0� q?u������Ԫ+f�����f�lI��=Y4�`�	�DAVh�R���$�z_�##�+�F�^�������`����"��r1�^FU�m������Z
��X�h���g����m۶�?�#8�֯�ʯ|�߾��o~�.vݸR.x~H���� ��-oyEى�n��_�Ʒ���K.�����v���*�L�>� ���z��t�"�O��� ,�"�@����~���A�IU�-Z�e����/���7���* {	0�d��r@��6\�󰄱}8��؜���9̩�L����/��-ȡ��g�
�x��r�c�����~��{�y�[~s�"� d���r���l�رc����֯d�'w/���(��;[����+qf����߅��"]d���Fh�}�C4�KK�H�>��ۏf/�n�T����4bQ��X�' _XDx�[5�:�m,�K[f�)ʈ]=��PJ����TK�N��O7�I>�MwMڋ{�.�W��P�"b����KeY2uܱG��Si��#��w�?5�8==�h#���� 0P[0��`2��I�W�#�I,犨8� q��7�����ѝŒ�&�(�g�R2���01�qZ]��[U ~�����87r&#O�Zh�]���8 �����2Er�*��l��@s�1�v�rM�U��F���#ŋbtˊ|̶oLM���4�r�SX��`(cV����g��E@bă�>�����^6�����B[Z�[t�'ۛrs�3�g�O����8�.!Quy�y��ܹ�V,cT��@_{��ǎI���Y����3mn�4塡!t���j5��=�R*g+4[ًfv�����e�Q_�R��4ї����I��B\���>��/�<�|�V'<��z�D�1� ���ţ��|ӦMk6nL.��6����p`���I�-G��B�Ej��ÔEP���|�ȑ'�x�\.���ty��^�c�=�e��#<t�ܽR���Y�f|~��p�WrX2�(�B���L�-[�����&''�mظnժUXZ�:�1�+�:�i�#�:~�)<6���C£G��m���m\�~;�� <{�l��Ƙ74��lԖ��r[n/���c-�c��g'�ۆ�vhi�[B+y��z�4<=2ڬO�^+6�o������?}��w]���/�\D���:�%��G����݂c��}����Ϳ���?���߯y�uW]uU� ��*���挏���?|�V+���#]�,h�����+u?�ځtuU B�q�[r6y*�w�e�}�k_ۻ��^����G.�X��}����
%,pe�;oE����X�J�T�	7'�����%�b`}&=��;�Q4�X�X+W�@�Ġ�(,#�@jA8���`o2����}�����ɿ����7���'�B%�2��85��ɇ��Z߀�Ȅ�0s�pP��yMa���~�X6�j�$Uqd�O 2A4P��J��2�r���(�ic.�U�G�6�2��	�p̬f��,����*���s�t$-Kf[����b`s���������(4$�6b���x�\���	?D��O� ƺE\�f�)��`���e�"�YB�]�J�t rw:�N�Q-��l�L�,������{���>#�����F���r�(��Qϥ_1���qvE��auW��c��
��ASA<)#���\WĎ�س�mDu{Ѕ$�� V	����"��P���0n Մ,��q
3n�UC�M�"W��0j��#��-	S�k�H����
�Xײ@��a���>�|\�����5�\,�B<.Q�ɔ��[+�i.(��d���C�Q�E�L���zP��2��Mf]��#�h�h�.�e��%�y2y����t=��$���I>�n ��=$%s]P�~��`� 8�E�Lz��rۘ�bC/���?пr��W�t#�I�����aLkvc&U������
\γ�"X��l��V�e��S��.�U���o���H�$ʓ_鬱�IՄ"d��JP|��ɘ\�}U��x럲�3om�>ʜg&��0����Z�l��l�j��t���fͶ�3��}�_8 Z��l����ݰ��O}ዧ�|t�Z��!'�+b���?x��y�Vmݺu��ߒzӋ4;6t�`��걡��3����u1L���.��@��'�G�y�@�qe?�}LZ�䀖�!h\����K}�|�y��
yJ`I�"�VF+"�{�ɝI�ID�;]R�3#�3�������5��*3:��nX�]��(M�*�a�(�m�oJח�,�}��N�G7�7��ؿo���� �l�^j��&��N��G�Ay��=�JC�<�KvG��@�Ġ9�/�6��}�굻�ڽ�ٽ�}�|@D^x�������Żz�/}�K�v�x`^p׻���cǎQ��8^�V�SSS����aݧN�����mo{\���W��CO�f`�J����!���t��C������b��k_�Z��ɓ'ї%@��=��֭�?���@ϻsMʦ��a(LL(y@L����k���nD�Q2��Ƶ% �r[n�-�~����AQ�R��s��X�������?�ko�q���A������u���]o}�?���Ϥ2��;���'>��t>����j5��@�~�3��u��k��榛n��/��{�e[�">��~��5������b��baf���[1Fi0��>��F>�����{��+^��������vv��jx饗�����=��v,���n6���5,���H
��p��Cԭm�A
�U��E��ÀA���#�s�i���̶T�v�������իW�߼����I �?��>v�]N�t�m������I�-������Թ#�d>t�W��6 ��I�4��n0��ϻ岵�υ�REj�~�/+vIR%�Ŕ;�C�=c�o`v�/����v��H#*�Z	��l@�d���oi�^0�h����i50j�Q��� 4���,�s/`?h�3.�[�ƣ���$�)����4K�9�oa�v~�����dR^��l�~�RC���e1�fO�sjJп*!v\�{� �%?r>�<;j��'��u}����3�#�Q4أKV�繁f��]4�1���n��`'�H���u���`��Ζӝ��ۂ+��3 `i�|FK��,Uv��,jyh�F%�}Dnp���@��s�*��������+�:��i��C�ã��\�&$�G�M�
|�#��h"�v���.�S/xiB��,��%������Ok�40����a�u��z�O?��7���Z��������?����2�m�f�{A�-�U�̍7»��]�b��g�䶕�"F8�b���n/��W�ͯ��Ix��Y��в���o����q7�PK+����噟����K+��EW�\%��X�Jcȝ�����U�
����'?�3�3��OK�N)�2������|���78p��nٲe�ڵCCC���0+6o޼c��K~P��wLOO0�Y/����u���5�\Ӽ�R��pdp��B�����	��,����e�1�<�ONU���X�����Z�-8X��:�t��8߲)!��r[n?[{�a-�Xn4�T������[��N�$Bq�>��>����k�l��^{�#�~��˯��߾Z.WI�N�+`�����3��6U�r�F���ڵ㡇�}�W��=_B�*f&zl�f����7��(3���v�er���5=��6����?�����?y�w��)*1��;vl����=�|eb����V����$>&K��U��KiH�X���[��oh'ӈ.ևn��/~�C�@������$�P2��%�R��ٳ��R�C�?��?����{�eWH����S����}Պ,��-
5�D�a�B�+Tǔ�}M"��YP�N�����L��zkBH@��ꥈ!�$�J�¨GT���QÀA��B+�1Kb?(XX�X��	З��S�
Z��{{߯��'u �
�M� �h���10�f%����A��ٳ�%Z #�f\Ԍ��`�2d��㇏`��v:�o��+j� �bS�1�Ԥ�P�?ʱ���n� F-.Z&*�1��W�@3�o[[Fm����E�*�\L�i�
Ka)P�a��ȱ�t1�r��e��}��4��/:e�`8���GW��)Y^Q�����~3bL�*����HVH�{��%���� 1��k�����GE��$�kQ�@@۽��1�2^�L[���%0Re��ra ���V�?a_�d�4�L����A,�&4��2��0�'O����w�4;����@��G��	�>�@xa�0њ�u��ڔ~9jhN�E٧bB=N�щ��u�멉�Y.��g0�."���Iۄ���j`1�ے�Q��8C�Y�u�(-�XO<��]]I��=�6��Ij:b}�.�86�^4����%͠폏Mᴍ�ϙ�I��&{ʥ�0֎�(��AbZXZ�j)W� ���b�0�Ȓ�V�^�d���F[��'��Y8W�Eh��ertk�2j�'r�I���!.�"N��,�>��R=按>�8U(B"���UB)"C��"��ƌ� df��
��æ,�u����h�p��m��q'������R���aBȃ�
;Z�L��qFe�#���&�� �^�r%�C�#N��@Zo��R�4�p��{ ����$�U#�6���n��|�I@� �A��'�%�J��S���X�sBQ���£I����虇��z� M2�b��(n�Ҷ�ɺ;�L�E��ss^��9A��(�ZA��<�{�e�O��wA�2�Zn�텴�֊��@&�q�v�q�Ng���~�;���ă^R��;�|�+A#����_��ߓ�,.:�W���_��ݠ�p�]�B��3��o�X0�]w}�6m���n�����M�
���$�mV'hq��N��!�Ru�]w����b�UAP��g�O}�S�x��Qgғb�`kTg�D.Wr�	�V0����&��h����<���l�%o�����E18��wA�j0��w����|���}]�apz�U���=_�mx_�;�-����s�qu)�4��X��m�ݽt�����׽����2���a�+���nE�4_%��-�5��.s�m�Z�bO��Gƨ��s�������R��Kqb�nkff�C�sB�c�w&�#^��s��ӻR)c��]����	8�s%�x9�ܾ�Ǐyn/rXG�I��$'��l3�k!���9#�<�O�ӘEV@/� n顅U�Hц&�rf<sde�wb�����eZA������~˼�i2:��Ό�٥����eċ�y1&���{i���̧�>AQ�A����b�[r>��h�,�y�fm���� Y>[������w!�?���i�_1�φ~Q=�MυZTu��$z������Ў;�䧞zj�ߵk���fo�3a������ ����8��H(�e�@�M?l~��Fޛ���i����8���������d��f4�M���/�|��-��CT###���c���P��:�c�=63݄^�y�� �NP{�'0R �g��VXR�|�P��-�E�g��S��*�9�Ŷ��6����|N����,�EƔ+85� qN$	E��m����H�D�|*�Nø� O���0l���(U��A����Љ'f��u��m��28�:DJ����"���D�dF1�&|^�fM�p1�[0��W��ꪫ�'�����Ӏ�`�GGG_�ݻ�{��ޅ^���:v�����+kjj
��ַ��iӦZ_�����߲�{�[X���쨔��`~T�b�f�k���+�s�=U�h�Wm��(�K����DE��\�������r[n��^&X+W�Q�RS���q뭒#�I�D��/URDR��D��䗼��룟`tj-&�G�~�c�����ZZ��t|d-S�я��G?��S�F�˘�t;@w��HVx�}�t��Ar3L��O�&��`?�l=wll�<Z	-5!���
v������w�ᬙX�+D�Ty�r�� 
@T_s�u�� �"�C#�dLUnn�o�Bp�#�S�JR�ԦD-6: ��\s-�h��ȷ���TJJ��w*R0fp��>�] 1
="E�*D��h���������r Xз��zI��(_�r�i|T$�>w|��BK-�i).��qjE�|Tfc�n���"%>�▇z�0�rot쑞.\D�Xw�:0P\��247���dujj�A�s�03X���jr�M~���s�Qko�������c����[���q��/�Do�L5�1�+�
�4-��%�@����Mݒh��4P�5����B1����V~��w:z��Y�o�
X�UK��#�������r�T��D�5A^b��A����D�G:�L��!�*B�6�=��w �� �q�*M*�h�S�*�dD"/z<u��]�RԱ<�&���ѷG�4rd���-S&���]���Q�ǅ�{����hi�s�4Љ�<�m��aڨ���.#C�Z��Jy2�PAjc�&°6:��]$&wדa<�b�t�^�32�W�Vk==�J �_rJ
e���v$$o-�ґ�EN#�@���C$R�SH�d��-��S|�凌 �j|�<�#_'����|� U�#��{T�0@����ɓ�N� ��ޏc�<3�����n������np���ٺ
��������7:8��9FB,��gz��N������<Y�ϟ��k�s!dy<�B��*Ef�ܩD
�aa:�,�A:&
�]Mq-/r��h0��+�!��Q���u����6"4_bL`0�����XY�KH�>����Gg�:��4��0Xݲn�\VT�  �'#@։�|���5�G��ø�6�����K.~�3{�}�l\�a���+�Gz���iL�:Im���\e>��M����lvč8�c��<�,,/�U �:t�k���Vr��A 1f��a1�5�TK2�m!Mr7,�7w┆&hŋ�6����bRf(�c�c�I&��̰������r[n/��L�V�a�shh���ߠb����@�T��%5���*��ɘT�]K��֍Ql�$��p�y�U��Jb�
;�Ȳ�XX�X�t�_O�U}i��O:nǶ0��ml u�fL�?Td�
B/�;�0J�aF*Z7���Ec������q����$i6�gZ�<�H��P�j�2�u� ��h��b���A��	�:�t�0!�0�{X�?K�Rcl�y�k_��}��6y=
���Rs�,Rβ�k>��|A����s\��A��
wV��FK����`*�s�9�{n�\���;55��C��,�I�k����OlT��*9�H�4b�-l�pe�[�k�j����2��ݱMP�����s�����o��v�;q����c�N<��c�Ԫ�j;�3���qr��^K��� �J�f͚���fL�&rE���j{���}���?r�ԩSBKJ		��it��奨\[ܽ��\�~�1/.���\�.Y��$P
�*�~ǂ���w�M��G�z�ѦJSlA��쎋�g��dɯ�v��|^�k�*̫5�>�ET�z���^l�� �hR�4�<0�N��O�r�����l@�E��a�lݺ��o��ux|F0��Ν;���P��|��P�Q#t^�UE�u&jcY&9r�h�m�^,x�x���,���gW�3;	e�0T�_��S�җ�T��÷�v��߾{��=�ç�~��������X6]h����H*�u��n��_{�^�n��
;81��$g/������f��k-hY�.�V��`�g3y�yG�%&^P"ǍS2W��k����3��fɜ� l�&��ƍ���t}߾}���i6�vV�m߾}ǖuX�{�*��kv�ȭ��b�-���gffa��ر�ޘ������G���_92R��6l؀R�݆u��bF�׾�� ί���͛7?�� r�:w�q�O<���~�y���W\q�e�]6�r�L=՜m�zoo/Ǿ0��!�%ܫ`c�c�(�`�7R��~��n�y�Dv�H[���_�Z�C�~!+q�-�_����Z�gL'} �"�5p5]S1R�%�=����t:��#*���������5-�aC���6��#���M*u j��\l���M4�׌�K	�ۮC��[z�#'>�F'�^�)�I�Ldo�,�SX������"�x=M	!����
�{��U9Ha�uA����<۲	e1����K���>�,M�C[�Ί3 ��8�x������]�����<W(4����݅B������Ν���>�B
�bPϣ�,��N�	�̨�O�%�%�J21��g� ����ۑ���T����f�Z��Z��7�	�����m�g���B�ɉ�D�7�oC�BC�p�.D�9���S�fk.鸶�dƦ���l�k�Z�q�Z��V__�n�'m�+.0�|����˥�l�@iZ ��CU�LP%A��Q0�M��`u���Z�:1T*����D&�H}],0��L�#����,J����E�F�H�����&��ĕ��Y>�F�$ȩi i�F+���r�t��}�"�LSX�6�����8*Q)��*4� em�����ߺq_��b�!ѷ"��P"�)�8u����vZRƍM�hJ	i���zE�0�ŎO�XF/}�.pe�ܶ@Ś}a��:F��IZ���l�^OG&@o�;u���[V�{��N�:��~o|&�m������!Ӑ"� 5%od��2��kGʤd�����"M��.��Z|�!���0�#�7�431��'�!��i5�7nZ�n������̩#�Ƨ'����W��u�H���{�V{���֚U+O8[��h�.�^�`�2��@2������dK���F[���ϳQ-��Ð���T̗bH��"EEH-J��%�A�d���pA���QrDL�S��E��Jʴ��a�ii�������fd�M��r��sݑ��[���m��i��dA�q��>6�H�:�2h
6}�!D�*�[��?x����,<���ď�cG�R5u3�Ñ��r�<�7 �� ���ɕ#+� ;5���صk���ēO>	h�`9^�ﴽޞ~����n��aS1,�y<5p�-&N�	ۑ�|�DnD�n�� axC
���+˵ΰ̙��IB&	J��it��P�:�30�<H�e�8�Y���&�m��{i/;����1g�и�� ),}S��8$�B�"p���@\���2�T/3a�<W�|�(���V.�!!���
��ֶʄѩ°Nv2$|���+N���Ȋ]Xĕ�QXNbx�\�T@A�{J]e�]c�i��m�qI;*��^����xMh!�uj8���F��Pb�0�9� (\ʹ��|/ �0�ע�"XH}�:/�^Ml�b�F������ݻw?��#П8(!��3� �la-o�<�_Iʃ�7g�a8}��fff`�m�vޖ-[J�کS� \}��߯��ccc��ʎ�6�R	�ER!��B�ja��� ʞ��͙�=����4����H�m�9'��j��5+W�Y�f�Ν�]w��cǿ���c&�i)C�V�M���&�H�m��}Y�g~�O�?'��&������U���NǙ�f׬W�V䮼x �����W��3_A�)7	��<7�	��&b���������������<�pB,�,%������o�+dp+sU���bb$��[q�+�|��B�2Ә��		I"1���j��;`r �O**��'O��OK��e�<r�H���~�֭[��eVpn��WqZ�H�D�E�r ���-�.Z�i��w����$�ĔNy}Ѣ�J[��&(ǕJ��o���o�S�&�N����ߺ�w~�w�Rm�ςz=^o��_=4�\�r%�8�[� H(:EBr%椗�����l՜Ea��R<ϙ:�k!��c=�k��*�5��VdnA%bf�,mB ����g��W�˛6m�\'4��w���5]��s�ZY\K��R_��[
8n�\OOe߾}�g�r��W���O?��'?�INo���SSS��� O8�߸q#�Y�9===�>���׷cǎ͛7���
� �a)=���''ư$�ƵD��Q4�{W�E���X�Kߌ�f�5��JV�ؐm�Z��D��ꂚ��&���K�<�Z�뽄�q�-���e��ҍ�8�wR�LK7�d�'q#�y��j�4�H���|b܁����q�	�=#a��z��x��NI
���`�7_j�'�E��kM����v�\�I9J�o:=��~�
 ��x�I�T��[ 4�
���`���H
�}pb�::�(GKq.9N,ܡ!���u90=�s-8'GXD�pN�>���w��w��y���"ͬ���5v����m�a��:�̓�ʞ�F�XH�_��{<
�)�o�ѹ��*J����Bo_yp�����=:9���C�����0��cˬ�j�
m��Ue�o�3\	�
���4��P��g���+v�X�ˠ�\�]-?m���=�1�a��Q�l1{;�.z������f�9�4\C�&lݡ"ȇ�
#�2ю`je@�(939U,��j��(���6��`��(9H�z,�y/�J������!S7s��tàV���]8��T�+��WFgY�Tހ�L̩�s#?�l��6�iv���#Ta�~D������)�Ɓ��%���2D�������[Krq�04bd<����~N�,<4E�k��g�"���MC[C�@�`
�X��<{���&��3Οmvʺ��<�hYe��
;/���/�n^]��C���� q�d���e�qȱǠ>��A�� Od��8�Q輵,�"���d?�i�'�0q�D��-���ٔ�1������z>��VN�:�)�b�*��:<<7�7+V�(t�=Ã�x�>55�FA�� >3,Tg�d���aq��N̆ �S��R�E�N�}Ο�z����,A\���-�N�(2�Ja�{�ca';�$E���'�}#
`
ۦَ#�p\,@�"J7g��8b��Ȗi�^hH�E�|�)@NH���Ɯ���T���`5���w�V�E���@��2�)
V��&w����& ~1$Wq�p��X� (z˖-۶�{��(��;��p��L:?11q��	����c�F�CCCH�T��c �����=t����`? �������\�Q��>����N�>1�}�C`pj"shE�����
�F��6�:r��2ˌ�,�!ԅԳ��������ܖ����k�m�gn�[,L�-D�.��/��Tze9��ӿ϶X�{��⟼4V��t] �w��z��

:��5�NNN��z�jP�`�^���k��t�G?������G-���Dj�+/��=66fք�Ė�ñA�]�H�=W\e� o�H��l�\�Af ���0��Бi�k5mێ�`�޽'�9z��������u�p�����:�f�R�$��D�8#s�B��������� �T%���^!�ctu�{��������ᓞ1�ݱ�W�����67(IIV��m�2C�]C B_�Z���:"��[#�P@L	2qшTC��t�{qzE6{�'���7����`�m벛��G �r��b���z��L��e�a������j`ǔV���\<XwU/�sk�/�NW��bOI�By v�������<\�R.#=Lȶ��M�?6����.���9C�X�E�}�M��Y� �ٔa�l6a!Ⱦ������k6l������ �NCo\y��ny��ggg�{�9@� �d�o�a�9��C�yJ2�����eZ0�l����b�!θ.$�0��Jݞ�y���	TF4���uR�����,S2�/F׷196�?<��S0(
�o}�Ũ΁
�Xӕ �o��?@{�cR�`B�C�Ee~��`�7f�p�l�� J��
�oݺ��믇K�޽n�Մ�رc�O`	>|xϞ=�V�دV�	�!�6y>�{\r�?��v��
'
0��
��*"�i�����������*C�QH�C������RN�,�,��=��u/7��9ߗ�r{a�e���|�Eȷs:����S��2�s�X�4���LH��Hr	->�LNYnigpdq˙��>Yd	N����䇨��4@z�<�;2���PiٿZ�u�9zv\� �>�@I-a:@������ѭB�ع��kKmB�5�h����G��oPq�P��;fep�Sj���u�k�==�'���'O*���k�G�]85;Pf�֍�����N*�k��A��ʬ;��<��~��Q����X:����E�msF;�Gry�c�e�
&y��m�Q��M5:�mԃ����x��r�����|l�@�?�փ�R��u<�~A��d��PXP�4'O�~�o�V�n�BA�.aN$��uv�	��*LS�2����!�q�S��Ĝ-&��L`Q)�pc�-����5:�=�,R��i�d��"��5���0@� 4�8
�(�v��&�WK�m�K8��v�L,�i-b��5V\�=���L�Y��ĩ���$Z~w�1�Zl.Jr�(������x�;ut&�!X��U�s6>gx�3@8��2���x�J�R��.z��p�(�
6������#s�����t�a���<E!��rq���XšX4��M�d,p��#˄�%$C�f�"���Z�����]�xA��M֏���"�[��#)4��Ls͚5�kV���W�
Xw.�����Q�X���>��/�.������m���+6��:q��cu��琋�m5��8�b',�W��/E�	
ymXx��W�f����1�P6����GI�
"����R�&�~1�ڊi�$���3�9?ƒ'��G����'<xd�ĺu�`8 ��M����vz~��x�\�T��XM+4��²G��ec��#O�?D[ٛ�����Yq�9�p�p8������ u÷pG�{����_�)�j��p�l��v��?��#��df����۹�*��z���,�Q�GZ� �:nL40)m�1L.S�2�5�j
t�Ǒ�	W
=I-�r>7�R-�T���r[n/�����v�EG�OۄN�u-�}!�x����6�3y����^�g���G����[�?�O碦8Z���F�y�U��<~���&d��4S�P�N���-`���e�2��ٳw�ީz���V.W�@�0�vH8!�4̙!vx7$E�F�40�z��	㔍@R�v��1!��(�z{���b*k66vJP�#�!{��$l0ʟ��+z����;v���O?��`m��P���h#�U���5��ݻw�߿v�`A��+8��>'X�.�!+!��U`�?��0�(��{)�T)�0N]���AV���9�%�5�Zb���#���sD>�kٓ��uϜ���'ts�R������n"�s���`�Z���f�(����/��f�tP��`�`a��ru``�\�D�V�4v���"���	#��aq<�Fk@>�2mJ,g���~V��0[�,F�Ֆ���!YT�D���6��[*�� ������^$�Դ�~��z�x�e���G�=�� h��^��5��������n����N����܁��o�]�
>�D~��<%�����8K�Zg����Z6.�L���`z�,�l�5*���a`�I���Ȕ�p�bao��0{.c�a��nҺ�Y��K.����ah���o�1���;��g8~�8z�1y,���f��`�E�	�������������r��3�=��W��<��C=�ⷯ& �G^/���[�bů������8`a�(���b?��M����Q�B������ܙ<�yE�m
���H& �L�]xnc�Y:�ή�c��vr���W,���^H�%�Zy˙�|��U�X���M9(������(�V��^�2g
"!����l�9�����^�-]�+�;�W�3}�~�=a��y60ޙz�T�e��!-�m!������K���y�������l��#�	e�0>�c��D��6Z�҂8츪�����ܚi�O<�x;��ru�V�Mq��F���A���у��4�`��,���1�ɖ)�)�O����|��1͢�,/\h��s) ݮ�����Ixp@\��] w�����j�-��R������щJ�3燓�c��9�6��p�-��<y��/~��yՊ��q�D�4��X�V4k��=y�w��]�^��>��3����+_�ʚ�����ܾ}�? 54ꄠYr�#3ǹ@2E��~T�2�bW�+H� ���,�SB��@��C$��N0T\Yu}�̻�S��8Wb*�zX|	
�x�s�R�Ũ���X�Jݬ�j�������O�N�(���`̡G(^<Kb0y�6��9K�s��ML%�����DUHX��&X������l{'?��k0�NE����}Gs���O�i؀%�}=ox�L��_ի%ϔӝvQ�!�r,��i�~��ډ㧂K��*XJhjb������z����J�iD��|�ߺ=�h$����Cx�!�#�BZ����{�70 :��'����܏���v{��g��vL�c���e@V^tn�����%�/�ˍz�رc�\�d\t���������!6vpC\�J�Y�fe2��k��I�ϋ!��5f��u)E����z���C��.�`��i׭���B@`Fr�RE!
�$�PK�7P�/rm�͸��s�Y���!�l�lӚi5��t[����.��]wL��Wn>���������������l�|X�Dv՘���1�B&9c&����f[��l}f��]w�9��+�JW]u�>���/��<�qx�;������߿�KP@�����+���Z�b!�b��������}�s����[ �z�ǎ�:�}�����Pl7뀯
&��-˞��3P�8Z�C�$#��l�-Dh�|ad^�m4�ڈ�}��{X]i�D\ً��`]+�|��R���.���K�~	��ϥ�4�O�!bg�å6��1�@g婤\���*���^�IT.��C�b3��<���Pr�Ѣ��	��4�*�+U2ev8 Zk׮-U��Ѷ:��N#�bfm!��� ͘�	2�FQR[	�q,����s����ƶ4�9 fffLʔ`g(ݔ�R��.Ո�Ak�]1p�С�sAyՎ�V����ƃO=	O[-������x��U�U�^�y�k֬Y������W_s��6n�;
�G?�wV���W`�t�<�U6}d�e�
�z����ݞ�Q�.͞�n���nebC��B(�,�!F4QDX�K�AL�\��T�K���<�K��,�ꌧ��ₐiy@��<��<�aK�if0d��.��`��3��h�[ ��h1VP=>=��~v����&`fn��ߵk��f�TƠ���4{�bY��<9u�j܉8p��e���e,�gq�g3$[�������p�%s�d_
1��L���ǐSn���J�2]o\�ő�������[�nzr
�掔�Z�3����NOo�UW]��y�}�������~�?$�C�q�N������2��K���I�q���Q��@�Pcr�0�R����J\�E,��A���զcC�9`��xi�kF�b��x/y#��a�?~�wp 5���X����[@k��+K��
I�H8�J�9,"8����}�e;}}}���گ��mx��������8���꧟~z�޽p�Z��u�V�Z����@����v���_p���{?�;8��g���O~2ݘ���+�Ś�a���Yx��[ЛE)e�B��JښLB!�V�3�
�\wV��Y�ܖ�r{!mk-�d5O���oQб�A,:?��1��R����t��e7b�z�3��$Y����Y|d���ˉ�]�9/��Kf�G���n6W>�L�x��K5�yt��=`qX���ҳ2n��%5L�bL�P�lI-B��PG��a�I)h���)�ill"�R�:;[/˫W���k ן���;��WR�i\Պ�7H������5�wɣ�ۆm$���k6=OZ&<��\]�+�*6��,'��~�p��[m�A�j���^���]�'&�&G�P#���)XZ�t�m?�mǮ}C�W��L}�?�ժo��&�!�������~I��J��W���nw_�%�����M�`�B|����1�,Z3�H��ܐ@O"�A
f ���!r�����tBd
�P��)�Ņ�$��U�4%� �d�ڏXM�`���hLa' ��q�(Ec�̫#2]��s�f�g�:M���D_�0����.��D2�aE.P����f��J��Z�IFx%#P��U�qz�z�)��,ۺb�%�����0(���0���Ss�%)A#Ԧ����>�F����QB
Sբ�AK�(�0�]���[s��CD���<���z��K�<��7r�xޣ��y�A/����ޣ>j� �|��*
��6(v�H�����V��~��/޽�'��
��~���MГ�����O�MF�JuljV�Њ��/���{���s��ɵk�n>w���xk����m�  ����٠~f�d0"�\�UI���쯖�/rL��p�V[c���Hi�h���1�D�
Ϊ𑿥{����6ɬ �h�5⎯����<��z@��]�������}p5@\����׽u��z��FG�H**��EA��N��hH�أ����n�˵2 o��O<��SO�:Xi�睿m۶Gz��ɓ�=�#x�6���p�*̫�o�yӦM;w������۷��xŮ]�tA\�����859�q���P)����MM����0+U$��D&B�4�A���ĭ�܎4>���c-B�H(1��k����4�B�����Y���m��r�e�u�&ψ0�{��֍-��h��~���O�#)^�>Z<���V¸�Tn��B@���9�cb���Ǚq�X���QOO�S*QFVÜ��%r(L |�}.���X�x���j58�5�K_������k��thvv��CGGl��Oδ��i����4�1�(�x*��e� ��s�=711���w�^���+����ӻ���HF'���9uj�ƍ�0p�+F@ɀ����w? k�%��%2�b�6y�4���j��UwP��N����0Kue�x��%���2��H�lTQ��Ȼ�D�y����v�0�	M���`xl�1PM��r,�?�c��<�-Lp'd9Cg�ad�d���i#a;�OG�u���-I]j�t�M=k���&f&��:@�;�쳠�:�U���x�!#��iF���thhTI8>16��x�����,�.�xhdJ��s�$`LS{��D2�
�5�T@v��V.�B�������$(�������۷�>�|�X��g>7���;9>s���dǊ+�L�7XS�� ���r۸�ӳ��c"'d�)j\��l4^��D��Z�/Q�\��bdc;���<qU�K�f&�Xf���[�v	]]�P(Z��Y�m��#����|���CÁm���Y���5��k��f�2�-��9=U�L`��,�4�Z������G��i�{��CG���7�p�%�\���.����.��!��c�=��0%�\�ԩSp����������7��wh ��0�@V��-�1e�J�*ؔy���{Q��D��g��d�Ƅ\�{ڢI���d�L��ܖۙ�_��B��:q!��Kܫ+������w��/�+��]^T$����wd����4_/�.y_V��E���Z8����!�(�)��u�#����I�I�
��e�mj����
n���1�OaI�ؗf,�T��.ֽ� -�b�$��l��L"���fZQ(;J�VAٖY){n  J<�%�(�l���20 �|��fgbz.<.g��.���Zs<`j�a4}O��g� VT�-tĝf+��E-¶S�k��Ɯ0cn��	�Un�C��X0Ӝ{��JИ�^t��S�Ap���f�޶�r	~cJ���֯}�MoB��G��-��s�����/}et��F�'�?g5��'� �AEKDdz���!]����Ɗ-#4B#��8���`��Z��Yh�~�&-F=	q�ѥ�Qe�J�d ��p\hm�V��a&���Hˀ@:q���K}5�l[E����}ۏc�!gw���nW�g�G�;��ĺL~���%�epQ���ӷ��)U.xRt�ev� .DPЙ ô,�󤁵�`�C�,,��V��Bц\*��&��l��r^�L��\ߕ���7�����=ޚ�ZY{��]܊"EI�Lm=� ��ex�B�´��g{~�f ��xd�hZh`��%˲d��E��Dm�������3��b��s�x�����i���5��z/�ƽ7n��|�|����G��w67vNMO$����\ݴ/\�Ծz�(,�=�� �Q9��U�vj�I�k���\kc�f�өP��8�TJF���򶧛l�?��]�7�i�G{�_���,랑�����b'GR=�K�{(2']��hB�!+�-fϒU�ù3��&�duS�30����?�~����L�ˮ��O�����j��o�k��Z����+��Vg���������Yrv:Q/�,!-,�`���,>�2��v�k�=k�KJ�z.�H�H�P��q�dFL/�Hl�2!UB,�gF�2�V <��@5�uZ`<�XAZD4��=3{�Y�,�� �����r#5J�}T��� @�Q�(x�S�Il,��fi@X43�E��0l�[�5(|ȑ���֫N�d��Ɍ`	·�F���ٹ���͌_�~�V���pp��d-�� �O���i{���2�a_I0��h��#��I����v�$��Vn�!���������llw����q�ܬ���Oz��j����p{c��h�vi�&��_���_�(�~�������Ϻm///O�L#E)�r���DT��M`ڕ&��@
Z�����V��$�Ig�"0�b(�����<�5�%���F��R�"��&M	s���6p}�1rctՌҵFm�ޱ�7��Fm��Z�,�4��E�*v�'Cb��+q�>|d�Rԃ�$�ۡ�X9&[�foS|�����k����c���[�+��
�M6�M-��1��.?��'�����)�d���lmm��^�b`� !�8��2I1JP�En&�4�B������ک8�OMɖǂ0/�/�_��g?��O>|���|�+�^>w��4�������w������#�����_�^�E��涮� ;�$�q�qM�E�`�8+�*�'r��,q+��LE�f�h�ǩ뺦Dąr�9e����^\�(#P�GT1%�R���9-�
Q�*��Z�����g�Ȋ�a�l�[��NENF������<r�u��Ӕ(x<9&��*��b�<o��b�3XW0wE\P�����O 0?~�\�������g�/]������O��'�j��7�[�m5"B�����@�0�͝]��W/�G�.�`�@|㘇�H�fK����C:� 
�Y�~���WK��]�	�]���4��J�J�@s�2�(]���k��w�G�G��`~~��Bt�ly��9U���o��������ѣG�m0�W�^m6��D� YA}���
�̑�÷�Kǁ��b=3!�4�\ل�9�1�)�ǐ�m�3�:���ߗh�{��׆IJ}��R. �\+�5��.�
�`_R�tg����>h0�\8����,^f�J%�B��3͇~����^zissF�|v`�la^��\���j�Z%�:�P���z0V0ݻ-�^]]�;
�L��;N�<	����?���������|���������n�Z��>��#_�¿y��g/\��կ~��ۿ����]����C\R���:��bJcB�TA!ӆj�=#���z�H����m\�t�K�8�6j�$m��Fm�~զ�c83̠�Nz�1�'K�n���qJ���Cx�"a��Gk_�I/�h�Q ��4�:>i8�T�� e�"���A�U�ֹF0�w�Rl��3P��q�(��A)3��^�`Rܼy>d��́Ր5aU���{�	w�T�(
1�+�}��
6�tj�n껝]�nk
+yi�v?�Օ���͕+�Ｇ��h�g4��򣨷r���굵��ϛ��Rd�N��G��2%j�7
�,ALbX��%N)k@�\+���HF��-��2Ud*��̎�����n"��Jtǀ~�$�ʑahF_�t����"�:���H!L79o5��vT��X�Ċ���%�*�0L�ڑi���hX�Kq��O�<3�6�t_��`�2*E�<��D"����`R^T$��(�m�8+ d~N2a9�z��K3���ċ� �uM�8�Jƻ�m0�)L-V,㖧����=��Yz��t��t;V�4"I�*VZSBG\g'i^&�(�%2��Vc�Gϖd���Lq��6 糱�O&�L���':�84��ki�V�iZU����Ǒ���3P�?�+X	��T%S�l͞*�	�� ����g�=	aiqhz��i�a��� �iv�G/��H�V/
v�6�g�߃�`@���� ��mo& j|K#�4�U+5��n#i���q�0M������^F� �\�O��,� H�B�b$��a"k��[�dj�å�����/�5�(;�H�|���~Y��;".oE�`I��X�]h�sD{!z��Z�DA�<�R0g��Q�'AM�ݍ������"BSL���.��|�ԙӀr�84�e���~����c�`S���6m$AB�-�s.�b�CدX<6[�̰|B�^,}�ࡒ㢦��Å��X�ksP�+ܴ�����.�|�đ�d}b|ms���=�������a�	�./�u�].����&8Z@�=�8�1�LG�263�̉�4wvL�*~ ���{�� >so�G@k�F�����Q{��b֏�2V��B �0oo�#����M���(�F'��M��S�ĭU����@^�gϞ��hmm���H�$Ḑh+4�mǁ�%מ���/�� ��cǘl���f���7P#��_(ԫd���aO��Yp0M� R��o߾��8�cXk���d%�(��w�v��=��3�����׾V7���Y�.SѰ����?��Fƪ�����nE���f?�$1��%�>�yhň����윀"ZAP���r ��:d�tʣ � n
̑^��U�uD\��8�=&}��"���(-�8�)r�$Ɔ�)�7�L�( �g��we!

N���އJݞ��l�0�0��I����ف͎^����)X�T�	V��C~9(�?��.�.X��ᙋ9�P�c�=��o}���_:vl�ɓ'�ӧO����cccH��v��R�f����5����I�յ��^<>�7��qx�V�^P�L�9�q�خ�Ų�B!>��T5��'���LEV��G����?�L��*x�GƮ`}�8Пx≅�ET��v��Mx^f������7_Z]]�1��ql�A�Z㖨c>�:�L}��?�����<,�G_n�o�*|��Py����s���S=�9MNQi^YA�g�dK�bR��N2�@�ސw�g�ݖ.�B�����qʊ���Y(����7��b�U�?~L���2T��bh�Z� Q3���/�|�ڵ0�a/ňR�XXX���ܹsǏ��ʤR��O�WW��J@��+ ��{�����>��/yaa������9�(��(<N277�!�/'���	g[^^��?��?��?�����q
j���?���?'$�+
#l|N���"��Q����U��V�ޮ�kITS�{�D.H��g����=5�e<j����k�ڨ�KRg�9حV�����`���b��JS-K3�YO��H���Gt�)����԰�22��^.��J�B.\�ڵյ��Nԥ�?�@;Ͱ����V�LJoQ���m6�^�@>�q�&�ofnvnaP����^�rEb^ZZ��m��:*��\��<�tl�n�����
�����D#�C�vOԫN�~����K�>���_�t��E拍��g���Ϝ9Õ=��;��gQA����l����fq��Odb�LG�bc�sR��a4��-J��RO��5Be*	�C,x�f`Q�y�0�2Vr�����j�f� �a�O��OO�T���TgU��tJ���g]�.l3�yD0�&f�ۖ�H�r�(C�48@�FY �l�LWt]��0���hmh��ԳA`�b˚3���(QH�ԗ��X�b!�@�K��g������L���Z,���(H�d�M@&0�p!-�q�n�� ����<�=�9���>z��;`9����7O'���f#��i�_0u\��eYE�h"M`Y���ۭ�V�6���G�Ϸ����!���>������iɳDr2+Ns�i��N\�B��|���z}��r�	U�QE����5�N�j�^�-�Z�웟kL��޼��(>[�Y.M �l��pRӶJ���B�J���Ϯ_>s���cGV;;幉��։U{�ء��F��$Fcm��8Ÿ8+��^���'�{ &�Nw�e�n��Zm���P�T��'�BD~�j����h�d9�Cqo$R��%/���TwJ���Q?r��%$�㬙��lͲ��a+�5,4˰t�U	�3�K(�.�dUC�ҍ_���S�������%�*�c�/�
�0�R��C��)N5�Fa��eF�!c~
P�C
V�cظL���R�&�ַ�f�Ā/u���_�"�a����`��[YYa�Ņ%Ԅ��W�@N�,n
�:�8�y*�!���[[�|�u{�ȃ �~}��V��öW_}���#G �m�4��N�u���6
�������dUX'н�gϮmo��o����cQX�.�E^�]Q��0�5�\#&p(-��ہ�'�XR	���9�U���y=�g3GkÎ�<�T�ڨ�گ�FXk�F�Z��p�_3�����Ɨq����VlN����� #�P��1Bv��v�Z ̬�|��^~��>'7�� /Tr�:h1�m�7��́Ai��m�"}?h ��>77W����k�z��������lYD�A� SmlmO�Pi��7B(��l|�(�rq4���ֵ������?��hƅ��e8�'�y��	ok�B�Z���ھt钿���FF�Mq8ECU���NUtJ��8*n���l�d=[W�!9q�phT�۩9$�G��Yr(�)-d���R"1�SMۤ�5 Y�#L�I�\�O�%ˁ�d���)#�4KŐ��v�{�Z*_���_x���R��n���e�+��
r)Ino1�� C8K����Nskk���XKf���2ۺq�ԩS�[�)�?v֪�C6��?���"�I҄���$E-G��5��T��Ky-��[d���"A��bnᄰ>�j�뮻fꓰ 'R4a��s߾q�F`'|��Pk�����Gkkk����!o\�򼭾����L.@'�
|̷C��S����W�6`�=���N���g�}:��$X�޵k�^{��{lqi�t��}���h{����q�1��C���ރ��&>JQnO�"��I�*�'>,W��1/��Ds��Y�⼕�����V�n�O�y���&����K7�(Z�����kR�\8�ư�P+�NRrԞ�+=A{��9J��Rb���
f $2��6�����4�_�Xfp�Z��?[fLy�5��Z���Cr|AWd��#+���J%��w�w���%���{�|������_F~ll���0|[������.�կ~�{������ ������r�
����~6����8w��>�!!5X?��t:pc,��D�����̔F��I���!^��Σ�)&��*x��#�.���6j��nm��Fm�ޡQ�����x肇WNy|����W��P��ڇ�j"*_eY�Řv�b�'��������i��k"F�A;�=�	l�6���v-�Z�f��L��Z�)�.SpT.B-�D�	�&�F���s�b&��K_ �W5����is����0���1C���w�H�\#!@!��ě4LM7�A����
1��9{�������G���8s�F���۷�f��A��U�ow�0���m*��3���Q�dhiR3I���`l� e-�j
�!��Q�`lL�����R�T(MfI���";��F�!O"S�Ȓ�*��
]8AR�RÍ-8E�|��"���V���4���3�L�X���E���3�1(V�HA�R�'����e�4c`�h������"#�ӡ����⯡W�K�(*�6P�#|��~��I�)��V`S�.�g`g#��%
ǉ�D�Pf>�f�|]��Qq�/?��ԩ��6���b�ˍ��a�I�GX79�.ų�,>ϠfXR���i��a�Tf���x�@�_�J� #떬-������J-�K#¼�������J5#t�V���SO><���z���b~K�q��ods���:���X�yi�[��$���=x�x3�Oϣ�w�Ӂ;��jD	�8 ۜD�V���8Ӽ0�������=�:fMU�Ru���sR�P���8Q���r��t �q�DA��ށ��67}��4�Z.a��ǌ)�k����6��KM����Oqy�$#ך���#`��j�����Z��%T����B�����X�Nk�q�`�)k"�F��O$C�����WY�=RY���Hiahz��\&�V�1=��"M�u�	-U��C����¦���:�y����ԤJXL�he/�\����I&`����[X �O���BiV�ء2$� R* |n(�]��0Uϭ8�ӳ ����ٳgYcav���C?�0��gΜ��xuu7�cG���S,[\��X��v�U���Cǖ�H�xii���C������O�>T�="Xv�bZ:�]"挚Xą�EK�y�@?��j��
�R��d���ɽ��TZx�s�s�ڨ�{a�Q�whr����C.�? \�	/!�BP
+��@2N�l}�B�@&De\�	����A؆�eL����K�=�E��ٓ�YOuR�#����U��Ế�>|xvv����r, ER]��PR�%�Xz�f
�Q�����@Ny�$d7*�5�rmm����2��� ����o���֜�ԇ¼���P�+ta�� I1)�'��iip�ݽ�6K
3��V�-�F�ie`�F����q˳��Be�;'h؏;lA���A�a*"���M��ri�x�M�N��u��E�I>�|����;�I��
+_9�s�^\��RJGr�X��^�
<�{�H|iNn��\��,Ƃ�[ځv�F�&���C�0:�"���r�G��#VL����om�+p|h[�f@��G�Y��
J3XI����'W����?q���ꦑ@V�?99933s�ȑ����v��vA:���1�i�Ei)� X��W��o�`Og%�8k�*��*�P�r�F���64&��[��b�(���lIY�N����9B$�/*�f�
?����I�d��p{���h	�4�;�QBAHbqy��Tc��y�uF��vK�e�7r6Z�%�_�?�L�ݭ�����������w/^�x��1�mc���-�܂?/��������Ç0�ccc�W�<�V�i����իW�& <�?~�T*A�����g��0p�|���^����p����8>��-��`N�W����)&qY!�;�nb�`����L^�^	x�1`ŧb�Fm��Oa�Q�[[�Z%Y��KE�w[&��rL��2
2C��a;(0!5/J{��c�1�4]��̲��^�����2���(��&UUuʿ��6GR��¡�j/#���Z$r�cm�e�Nn����}���N��x��e04�>1Uz��Ǘ8t�Hk���[o����ahiz�Ć�����M��d���H�\+�U���`y�� �g\�������-ժ�?��'>����͕����_nmm]=w�Wq�7P�+�",�Xl�4��$դ�P������Y�L��85�c�`���4U*m�jrI�c�!'n�Ans�=�ICU@�#1vH�D�e��S��e�d�����f�~�G;��I�IP7�A@'~/��H&�N�+g`�w�XDq&ox� �4�4����6!�[R��n!2Y��   	��q��|$*����ˎ# i.��RRi�	8���PXb >�֕�*@v��,6c]���4+s�s�Ⱦ�z��al�b�ӹ~�Z�G��̭��^�<~h���ʵkq���K��"uI5
�j̈�M+�b�JX�R05��ґ4����CÑ���-��U����%q/Ց��XMN¤ӝ.�J���Bml��>�|ׅ�7�˟}��g0k�q����|�0��]���]��f����j�:�P�v���K��eip�2`T1W�B�n>ef�p�z����X�_�����j�b�莁>��=�i]7�8�t����#�u�^��=�>��D�@F7�-�2AF�4yR\Rj�oBD��:>J�Tf�-��Z�\)I�_<���ቻ��}O�$!<M�K'M�� 	�W�a��&q�&�S���S�i�י@=ÔR����/�`�4ؑ�@�à��	c����
}�"��;�>R�jW+[[0�<�����׌�-���%y�<a��$ʹ��u��Ȱ,� ���_�ƕ+W��/����¿p��W����W���R��ST`.
hg0�$.>�gas{+�҇O>��#����?��7��� �^�vy����~��Ǘ�������7n�8w�|�_��ɓ'�!WWWa����,�
 ?��.9kkkI�޼yS:�����7�������Y�CZ�D�S�b����g����/��"��w�Ee��#��)�j����(�O�&į\�r�F�}a�Q�wh9	"�k@��@0`��yD�)��Ű9GQ\+��m��_L�� C�
-��7�F�Q����
��3�-~������f���>�P�a�������w��XI�����vaۂ9�
�d����2֠C��`7pV?^��n�	�Az���455�Í7��.3���+btң�@�BLѰ�a0h*It�J��j8zZ�,D���.gN�G.F{E�jZ�o�'�v��S�ɂ	aj�̸���4ʳ�)sM{���%(wG�r��8De�<��t�G���X/�,�� �Qv\�b����y����ִ��"%�\��`Ø,��a�|�@!�*�G拜,锸R��k~}},���9����k���6��� R��)�<'��a� Y��7�/���kU�o3�\<2�S�{*�bh^���#�Q�����@WaA��6ZX�v�)�¬Ĭ��),��A�����~?��T(���4^?��0.SU0bpr8�>�Xan��C�)�[M\ZN}�յ=;v�?�~N6s�=$O w�c`��_wvvz�<vǛ���R�b�9N>����q�z�Bl��^Rh�'���b�*�"�����X]�i���"����p�bB����R�㺗	�9��w1Xf��<=�p6���m��Tju4�-p���^��4�+Ɩ9a9���$y�����?���a��,w��1̅+������F������/^��z,-����--`��ٰۻp$�b8m��Rn �q��:�]�i��5��	~�[i1�w���A;R6@VË�W�RGm�F�Wl#�5j�vkz�dD4iT���}���i4��̀u��Z���*���i�F���e�[Xq�r��^��z�۝�b}��Y�k�"R�I���Ԍl�z��˻�n	�d��AW6�m�[$�"��O��B�/��-�\}��}���ݿ� X���Z���4���_*Wk5>�2�¹hI���X��j���惙�s���ѵ��z�7~�7����7N÷&�Z�q��1��a1[�����0��2@Cz�/� �,�PP��djpHf���T�P��8U�ѬTy�iy��j�oJ�l�I��(E[$J(
��s�֔r�bSO�<@Jd����Z�s\(���فr�pDS	�\T�He�D�_���=ah��Ґ�����]V���`\�	� :z��-�J���/XWR�K�1l) �i�fY�c� ��I�����1`�<c�f*%������Y1�K�Ɣr�X>�@2X�Q�B9A/�w;�խ�WO��؇?�%�n�?{Q0�16�N�_1��W�4��B+P'�F��@"$��8BE �����O轖�@B�\�Q��7<,
{�!�dh��j�ӄ�d���D�<^)����瞻~m��^Һ}��ol��V���}��4�dέ�����T�m�o���vμq��������Է������`�F= ����,�j�:;�h�o��:������յ��_���-rX �_&�����>������#��M�O{֮��b�'?AO�i8H�z�bH���ǃ�J\Q��`D���:9%f1je�eF�_����쭉����:����Re(��*��Խ�w���(�"n�8��B��$SN��Y�"Bt����H��A����a�1EQ
"x�y ��$��Lh2�#�>ܣm��壣n�FhAB�����)G���6����2��X�=���V���.,�"+׫Xط���	�hii	������0vb�I�!����1�P �rKo����Ҿ���?����7_?y������/����^_����o�q�-��'N,//����2l��ϟ������~�O��O�����o|���Ӱ�ള�������^S�^|�E�:`���I8L���]}�e�ʠ!e��E)޿�N
.Y�?Y>��J�T���U�@�|������L�i��6j��_�FXk�F����"fP�H�\e�݇}���D�%ȥ
/l�&R��qd����` |Py^M�MT�*lR|r���mf��l���a��̓,�� K�}��v@۷�q)�/��<��vƳ˜h��R�D�����w��2 ���0_V��t�8��x*�#�6�W�a�U���P�
��a$���� ���'��.֙��c���.yRn@q30W��9�%�a�u������=�rU@�_�����*拤��y�<��i���)��y�ӡ�<�S��a��\K�i�(���O1fx�"�;S �b~�Q����?]�������!)�1R�E'��~��c���©`���]���a����r�0�y4����so�A>!�;����E���/�]�yI�,�+4޾��PT$���0@��H��;;����<&�@�n��(�nV˝�N����wvቨ׫`v�/���~$�@�=�Pp%4�am���3�v��
&�aѼcj��ŋ;�.2~�s���k�>�F�ڠ}o[�yfAoو����Xi�R ~�S���?5U�v;Q$�̓�aU��ű��1��o�L��"ȅ	�_�J�Dnث�(��}��ċ�M���O��&�3�-���}�j�?�ʃg�[���}��+�5���P'�#B=�Y�J�qj0o�>�����˰�av qj� �U�1��L]�u0u���Q5sAB�;�c��wwQ�������Ga����+sk�	a���x`ee��ٳ�z}nf�!���͙G`�ok���t��ߴ["x����n�P�o6$��Xkx?)�.Fm�F����֨��n��E�R`�[+I�Y��b�T�c�^����JHv��V�����A� �,��5۶���E1	kqMF9���1(���9�EY2��C�'�[ۂ^�eĖ"|�1��3]��H���.�ѧN�?�|�����w7`���ה H>�+�	1�&���>��=����V�v�t�^����?��ϧ����ӟ��'>��s��T��k�])E�ofm40���Lݤlx1�2�T^JмK9�Ib���b���F҈Zc g�G������Vo7E-���M���ȫU��ߠ���U��d���+�N0�|G��%X�X&�)��Z����&5��"�1j�fcIes�~��G}�3��q��˲� 6��4��zP �i��$#MK�#y1�\�gus��$�0��2"L���B�	P���#�n� %��H��ǹd�N:"�@Vq�@4�42\o�}�CCaB�4��&��Z�ۏ2����J�{���i���;�k?�ы�2��566z�!o�eękX���չ�*�	"��nzFя!	� 	���z�2ݰ����S)a|�7�'��	.�V�(Ζ�P�"1gGR��D�慧�۴J���Z�ڹ�\�paE����7>?�8qr���������c���;߂)���u��{�]���?����a]�c���\mn��l������Jd=�����2����kfIp��y~�੟~�cۺ�ar|������7�Z��\w�����,/�^��;� �\W�"1�^��j��H�9H��>� J%�k��#����f�a `�>�8V:�,S0�0Iu%��?PZĈG�����1���jv:hK�ƥ�����	#�Y�ᗈTs,8<�0��kY��(��Qw�B����a�Q��b���<11�������7f�Cf��؈̀'��ß�,��5�f��1wOB�c��`�T�K�:���T��4�)��T����v�A�P��>���}�ck�/_�����Ï?�AX	�7��Q��jp�3��"dQP�� G iQƇ��;���z�gy䑿���O��?����������ܹs���'�������>�������w��:�!t��  ������W^y���{am��C�����Eh�����I
O \g��9�T17J��Y8�	nްO+�̄���x����ϻC�6�o�_)|4{��wx#�Q�Q���k�ڨ�C���H��؊%̓��8q�G�?� �kqM�$U�4��2z�Qє�c9x��6
��XA��A�S�-z�n~��
'���	8����
`�٩i�g����}��8�qB�	�D�j��'�MTfci5��\5�f�����
fO�8E@�	0��3O=bG4�Y�o[���9]$���4�@%���`%��C��r�Pc�����N�|���	:���p��cA��ۻ�&x���͵�]��� �����2?Qȵ����""1`�@�BP�w��^�Ⱦ���������v��5H�)n���RT!�@�^ �@���nN��4!�j�o��� �C�Sh�{�=i:����ԮF�?/d�U��K��A ��+L��1Q���\��BJ"~��U�\uS���AzL�P�s:��	OK����Jm�s-��+8&l��j���h10p�#�>&1 �x�HL��u�s�&��$I�9056�W��ġ������Ǳ���p^Ћ���w��	W�#XT�f��t8�np�żs]2ɹdR�^?`RtOŁ3�b�ϱN��c����	�i]$ݞ(&�`��A��隠�ŋ�������YȆ
�Obya�M�����M�o&��"�qY¡��Sl�9��e~fpu^ E�Y,���˛UX���������a� �h��W<C,�����IP�@���X�j0�Ը~�6�cTqnvv�y��q�:\��<x����A� ���o�}�ݰ0�w `�$�TMУ���`%�<5w �,�$
�K�)��w����}8̽xź�n��ݢ���m��5j����k�ڨ�Sz�HY�X�G3L�a����恲j�n�[1��R����k�"od�X&�h�0l�fAioLK��M`:c���E&޳�Fp�CX�E�['ą0�;�&��B!�Te^����֟�[��0�$�8S�eWKU���mR&�mq�EqFq��.M�����y��[7�7OLc��+W�d=��d�*nIz��*t�YB->t��ͤ帑��+'�8�&J`�� ��(�[��A��W�0�����	�R�#��yhRx�?F!�4.�рLI"��U���/�Y3}x�ŋ_���X:�lC/i����T!�z� ��s���০G�%�V��k�N��:õR�N�m��Z|O`V=��G"���:�(�(H ũ�*�T��q'�c�f�k�"J#i�B^.��,]OY�E�e���,�B,ʋ�ؔ�O�<�)�*��#�f�)������bf(���8iX�U�V��1e�a�w�č��~���g�O�}WiN&]@�$3$'��MLN�M���T���B����N�QR���p�t����Þ����`*YɎ����P����u�����uЮ������������g�;�\^]]]�@k���� 
V�����G?�1���������R���?=Q)�������iE	j��Q��=X0k���R�(��'�c�o"��&�Ւn�}O��e��v���J�k�et+$���FI��v[��fٰĆ,�.\���IL,���4Qb=X�/��m75 ��B��XׂX�$ڑġk���J)��1��.���W���0��r�))�H� ��EB�ØejV*�ZQ�.�|�Tb��qdH��BM���oS�r�H7`�o�Zvp��!����7�d�;�f������ԋ�U4��@ϑ�	�n�4e�����8DiT:	�ecS��Q"���&\���C=��{�l��W�^���>��%|�|.��<��'2�b�kG�`E}���p/G�e9�z`rrrqq����S?� % Wn�t򃏕�� ~��i5� �aX�x�	�~0ڀ���N�Ha��l @/xF����{&VS�ˇ��凜J{��cmqB�^��1:�ܻ�w�|/�W�ڨ��?Da�Q�wj�F������1�x-����oG�+�Pׯ__���R?.Fz�lU�Ǖ+��;N�<[A�0:*�چۻQr�d nՏ*���K�ộ�M��0\d�P��i�6���K��80�â�$���D�\��g����������1	�������1�W/��"����'�{��{`L``0*�bLK*R�:h'��$75RNԖ���4�	�`:v��~hG���o�r+�ч?�ac���`sw�0/�R���T4�2Z`=��T��C?D{�j0j�����w�%4Y�������+[[[R"�a!�2tI�
�&M"@"��S\XThǴZp��e۳�0�F�4	cf9P+���B��F�k�G�$¬$��?�СC��:����N;��R
j�\2��d�*J�عE����l�I���j|9D�Ba��r��B�^�՘���C��.���,���!�����A䣍ha��աʳΩHq�C�9o��{Z��t���O�����>�;�IYn(Ä)�?�t��:.������&��e��A�a4 Y�?~���K�v�Σ����y�����ħ���^���ʙ3��XZ�qpi���%�Y0�c$`_�tAJt��N��@-�����a�c>??��
~J	g��m�*-ZN��Sr�Ło�:�	q�q�bA9
z�"@S@'��>��f3lbѧR�J:��c����o#��J�������{`d��/�*	O��B�/��$-0�P���}Rs���:���7ov��ش�	��KH�]h�W�tzp�v�Q�ȟe>���U0���)3Mi�ȴ<��FQ�(�$�B�k����˯����O�c�����-�ۣ�>:77�%�XI����oU4�������u�]p����ŋ�`��$��Y��?~����� � 8���piiian�ƍ�(��|�B�y�WӃ8�\��4Q��;�։^���V0��@�>�>�1=kq=b��b�=6r��m/1j�6j�m��F�y����w���-+r���)/��R�f�����*s���[�J�LL����V�[�T�H�n��5UF��F,� �
5P�@2����ݽ����_T�!n�����/�&N%��Iv	K��o
�ǲK���D����]��lm��Ja$��<�^�c��k�N�o�i�65?L�l|v1ˌ���ʹKG���'�X���I%S��"�.�H���K#0e�\���Ӥ�{J�R�x>XHq�����<|�������Z�U�Fs�#w-.,���[�εt�T��e�:������̄̕�4����T���ʸ^q��ZO��`�����˗U/���om�7S\��*ʒ(��fj�'R�4�8�];��@��3��s3*i���Ǫ5���v{~:c�
 ���v��+0��2tC�K��PV-�V��֒���~�x�J��廏�������o���ͪn���6ڈ�U���^�A��S�I�џ&)'��$L6t�pS�!��?� �E-���eF�@I���l�*�sj�Z�ɐfM�� {NS�c�5Y����R�L3�-�'����"Mc���$�  ��IDAT���z����+E����ȑ�A�w��%�Xt��D�f6�����`���-�_�2�6UK#�9XYYy��~9T�ٕ:i �(�n�s�ch$Ԟ��/��K|业�h�tZi�����u�6� {}��);�Wz?_�qc��5����`,ɖO��)��g�_�^�z�;MF��馥g�6�޵I%i�e*�����r&���Yđ�¸��X$�~{��#le�B눞V_��4J}id�?	��Z�dH�1�$L8dQ�� #	�*�l�ô�j�`���7:ݩ�؃xp��}�檚�#,i!��;���]��K5/���^�D�<�:��A ij�-��N?��u#�J�������~�c`����6=��ȍX��㠇U�žŁLS���!N	 ���I�K%E��1J��ŬUC�� �lD*�X�З&�%Jh��{S�<�aĉC����n!M��o��#�:f�aDzb��,�\�*���3��摓'�x��_��{�c��x  OH)��93��p�z� ����adJ����f�ai=�|�/���Y��i&#�bzA7�=�11+R�X"��������n���)�w��	p#e�!�֚O2�� D��v���I� k��D㇂�X�.�-�L�%3�(H���H����Ig0�x�tL�o��[!Ey��6�,Ʉ���^B��9�&�Q�[�k�ڨ��&;V>	��8H��T�a�������~���Y{���)C2��̉Ab���H&�R�lmm]�p5'��1���R�D~�Q�LO8�3R��Z�$b��
ke,��n�_��"f�:T\���,�Ū���,���#2�f�<Ug~?p���Ç��/�u�ڵ��pڟ=�=�Zm���7����4y���;�v��^yl_��p 0gvvv&��o���g>cZ�{�J�`�;v����˗_��߿��+��4�4`��F�2ee����p�G?���ԧ.�=��k�ٔ�����{_��^y��*�C*F9J�l�0��7���w�2������o���
N=���_�r���r�Fo�d�k����U�<\}�H.�Y�Q�h�P�'����'GAH��$-r�l���f�!K6_~�:�2q͆�瀦c>�G����ڍ]�<S��g?;fU^|��+�ξ��ixp���XE�=����.^}������Zu�l	��r�(�Dg�&%�䵄�x��+�sc�K<���N'��2̉��0�nKĚ#+�]����K���5����N�>&ey�Mⴹ*�s�"]����a~a�81쩧���W%��a�0i���@�n�y>�a&?o˟aV'��H%�8��^����~�K_z��y�/��C��sѹr�k_���0�i!�ZB��c�8G�����_�O��r��:r�]��y���H	n�.y׿
�7ᘱ�y$�L����FE^i=aFתa����w�h������Ȱz;F#>�EۏJH��BX\u(-c%��2l��1��|!�p��`�T�h�����}����<{�l�Z�y�&,�O~���	ʖTT� *��p�%bzy���r��:8n�:Q�JV�8���`��~6-�����x���*��{�]^��S���
�&F�
�!����,*l����f#*̕$�3�N;�Ĩ����	�o���:���Q{_m��FmԄ�eYRE��4�e؏῎����T��׷��o�S�Z�I��af���!9�۠�?q÷��uh22�t���RC���vH�]���
�ff��0�����������U]7{�^��V	�(�a�	ƨ��y���r��{����NN b;��	Q�<	�1yJ%i��d�����
i���V�F�$pd��1���0Kz�_�7��jڑ903�㋍}�S�E�ߖ�q���*zm~"s5��m+?�n�����ZM�X��YX>d-̀u�^_o��;k�
W뻚�E�n�d�}'Ѵ�(���5F�BM:�uw���=��?�qO�/��jin�#z�7��籥�S��oI�E6��LW���O�1<]��������z ��8Z��0`��Sэ��~�I��ئ������Le1ҡ:]0T��I,��&��c��S6I��2���z
Br�vf��(��n�I�H&*�u�\���Z-��E���Tt��,�c?HP�#UU�u܇%ԍ�~�j&��Q~�/��s�m�o���[/�'��O�&�z}��7���P�N۷�Ե��Z#����g��2��I��RD%�ܰ�jN�� {0�l�i�'"�RAibU��xu�(���D�92wh�{��N̬��N[UD;e��|��,��nf�U��M��Ũ�.3�\��.���o�2��D�֠�2�r&d�I��$�*;� M0g�������r�P�,�&q�]�4fW�̙�s��*��R�";����!������*5-6��fSr 	���H���y����z��*��Ʈh�}�o�`%h�v�b顣Ѹ�Y����j��e��z׻�K�q�G�> �/1+I��sI��Ү�c����c�5��t&�?�~���:�y�fL�֡�D��l}}jee��m DP&��7���#�ᱎH��è��RӶ��>��M2Ǵ�r�+�fH� ��:u�ԑ�!�0��*XALC��,W��c�?��{��yH���Ǵ����k�/�����`��"��`L��V�82�P>���搨	��I����N�N��6����2D�8U��
�H	C��l ��8p��l�8���>�O�HW�z�X�Yn����3� \}1�0Jo{)0[��e��$��n1X�P�f��@^1
)�Q{�m��Fm��GC÷�]_[�25��A����v
���F�)�ưz�m�|Oi��V�������r~� �-�K<�k4\&(����J�����1���1� �,�΀-��[+++�.]:t�����ϝ;�"��n�g˽��iε��4�ߖ���k`	U̿?s�X'�s���RQ���������O�{a �nm7��ׯ^�4��EȍT("�n���Y0�v��S���������K`ߌ��a��*��B;,�s�a�9����'�|��9w���p��:��>��S���U�������ti�c�ffg?�я�R��^�:��'>�W���׿	�(�� �2�2<јUUBʱ��A�2&^��*Vt(4�r����*e�d�K�F��Q1f���ʶ>���,����g�y�$v��ٳ0���L���?����K���U�c7��d��Ӣ�M��k�r�$��< ��Hl�����`�K�6�PH̘���ʟ����%�.�u�����~&]11A�f��l:K3�Y�Ŭ-�{=��==Q���y�]з_��sЇ�8��f	Y�R����IFė��&~E��;v|��l.83���\�|9Di��6���C�d�4$2�3�xִ[嶋V<p^�*BG+��'h
�S#MHL�$��iL��sQ���
{�H� �Uh��m�{8'�yii�ĉ� 9?����)�-.fz�Kc.'��t�[�Q���m�a���ӧ�'�����\6���T���Rf)q*uM�1�3�Hה
�i{�ՠ��(d���&�+Y���Ծ��o�|���?����r��ɓ�>���ٟ����q���}�/r��d���
91��(Q�*�D u�𭱔h2��Ǆ��6X��P�0�cZ|/���	�5P%r��˹X<��yRUw,� KK��]������+2uq��ꂬ��.��o?��5إGr�6j��k�ڨ�j��=^���i��L&c�z��7;^#V�k)�釙K[�#
51�B�[ի����Nr���vL���-r�{"��:t���P`X��� Q���pyU+��:Z�� Ƃ4���{�&�����Ϲ��f;��;�VY��8�_�RCxJ>{*�"8z��L~�3��R��1�O��^�x��G�ju���W2�^�ɏv{���i�6�V�\��~����F�9���pͱ�0q���^z�E�Z��_���>_�F��ve#���dy�"�ef��0�JlA�$&�#��{i|���sW�{ｏ�X>��.�YyR4����\���X����°P�?�1��u�х2�o�m�ҥv��݀s"?��v�����#Gȼ�(9h���/(�(W�G�Pj6Z�X�:1t�$8������*0d�C�a�2:�Q٩Ķ�����v�F�u��;�fͳ�[���i,5�-U�=�Q���q�9?h�/�
�����y���i��lmjv�2�Э~��/�h��7�?�O������ԏ.�u���:��#w-�Y��`���ս��N�A�j?�t7���2�p��NX�K�*�0�A��(봽n�kZvOE�&|)������Mj;M�wo�����f�:�T�a�D/߳�N�n���nE��L#3�
\�n X�ꕫ�`[%"�_�����R��i ���3;�/�F�4���?�Nui�#д�7�Pτ)�0�Xπ"��x"����<^+��q���}XP�
��Q�Qv��=S�p�܁���iv�ԁ�-H�(�5#��^*�F3v)K*M5�̼̀����T˄���n�yZ֗js{k�ٸ�����K�ar�T.�c�]�bljr����,J��T�a���t'g��"h0L���T�l<T&�	��Z���B� �Mz<(��J-�TD��<����3�H	+ť�(��@������������/9N�'>�`��y��ف�0�5�	���e�Tn�a*{^�FÝ�RD����Ǭ\��P�Ri~]E��TH^�����Ĥ� aVJ�]�8k�J�@f�^%�4`�qr#��+�,� ��4�<��dJ3���#�(.d�?�K��ҁ˰��"N!n~� �\t1g6��Q�֨��{���Q{^��Jf4׆j�ۍF%�|�7�e�ȱ�������ڊ��m��͂"m�JH)���7�,�?�~�b�&(N&c�/�΢���/�^���q8��ŋ'N�8p���/����A��"'�^��B���0f/u�!�B�7�Z��K/��9����X$\�r�uQ��hV�c4���K�?�^j/K+I�2��+W�'�&@M�n����[]�'m�]�ƣN�"C�	#D��+W�6�	=>6�������F6V
��S�[f����T��w�=�fR�Bds�ԩS�����ūW�^�t��M��dmu&���L�Z�⢠��Q�����?��EK�1&��F�#K����*���ǉ�Je8�:��U���D�6L�jT�����}&.{s��.,T�|����7a�a^XZ ��p�ɾ�9<�^/�P��\wr������j��u-=+Lஹ ��â'�Rv��VNJJ��;S���2ۆ1I8�G�3ک�\XXH�(w0W���x�����q�˶��s<�w�YL�O��	���a�X�����{�1�>Lȡ�dp�~��lX~-�%����y�ÅT��$�?�"7c Spz����-���-����O���<�o�
�xg��y�-+B����Pg�$��)v|	&���6���͛��ډ#p��Ne'CL8��Ȕ�a���ߏ��݀�xw�D�$��,�fb�*����6� ��lA�o�u�%t�p5�Ǌ���C��&����0��J̧��"9��l6���C�x��>���O?7ˢ�<�0w0���3�ȴ3�X���`}���r�*\���Y��b�k����O�^>,���t���A�����-�B<� 8 �x�x���L�Z|_�xr��G;o�������N�.��"��Q����c�eݫ���Q[�6j﯍�֨��m�s���?F/����~?tL�ήt|���xM�E�%��H�J�j&j�<w�4����8�m@M�~����
G���zS`�ú�kaGIjSP��Yq,'&m�ф֐nY^���vm,�������:X��X;nlb�"���,����1�W�O>A��b�t=�B�(M�
w�[-�i�~�&X0뗷�����[?Mk�%���6�yYj������ę� �S�n����̒����x�2v�n��0Y�Oөr9��R�#�/���/{ok�u���3�{������*VqM�*R�Dɦ�6#E���� v��
' �4:P��ii[� E-�")J�dU��yx�|�3O��^��w��d�-���n���=g�s�tַ�Zߗ�v,�XWB%�б!��PCׇ%X��U"��/�����:�daF�)�kԒ�vj`A�f�/��Nǜ���� �8��Q׮_#��d�������{���k׿���=�0�g,�R�T�)���Glr��ՍS��Y���� �
�֕���B#���v�u�]��	|���zlv��S�`�}�Ս��N�-�J�T�Y]���|��ɝ�C�O���z�����r����_/�Wa����X�`j����v���*����ݍݽFK>U�x���[���j� :2�7_x����Z`�VkE\�� #�J-�H��L��G!�w�R�%�">>z�ԴT#�\/�3 R�nDn��;Q�gh�i��������a�>0[�������������~��Ʋ/�+W�����ۭ���/ui��.�գ�W����2����U����TbU�̟�I�@�E��F�\�5���G�f�'''��p��`[�ۛ[n����J�Ż̻�⒅�"��%p��@@�*� �BqJŽ[����WJ�(;^m�����_�p�I�۝��%�d[�6�]Y��"ZԐ8Q
f��a���u7I �5�����:̄Y�s'ͫ�_�m��	�@s=�����e&�p�8Q��L|J5��7|)��ľ�1�^�#��P3�&�,9k4`6M�Y���3!Sф*�Q�E���u5M	z�Q�˘C��)>��O�H�D�n�#��8}�4 i���dϕ"(�t���A�; _��%T����Z��ib�,���O�[ۥ���v���I�T%��͛Gׯ_���G��}�T06ʶa	Ê-�F�U*5R��u��f��n'�I��5��a5,ǮI�/��"<	����R��K���5]�τ$/%%kI��^#g8��%��J�2,��c�!��a�1
����uJ��vw������)���|�g�UI�A�j��`���ߞ�%k�K�����
��۝�og�&�5��i���T�}q�030Ɨ��X���Mڣ5�n:@oE�؝��n!���ݜ"�:ě煢Gt�ϊ[ވ�4�H��V' �UN;�F���B��mH���80k2�q,�tb#.ߏ��}q5eNgMB>���y��\鲰*���c`<�*�Z k����qұ`]�}��p��fI
�IW$��m�7ɴ0�����`�	S}饗�{��G�m7������!�R���#�~�3����x��dQ�#?����1Ty�0O�:u�ɓ8��5����k�"v���)�"G;����Ν�mJ93��H$;"~"��B�ȑ#=�eE9%����0�5����sy�ޣ��g>���{ai���˪�����]XX���Y�3��Df`������? �H]/����I*R��4-��OQ�~��t\"|K�sk(����$��Y��(I�1w_�FҁIR���͗_~Y�$��Zh���ul9��q����^�R4I����P,��{�8s�Q�8 ,=��J/놦�.g.@%yD%C:pyy9���S�S�;k�V��3�wCQ▜��N[���4�4��H-VH��ӟP�;����	|���A�Δ*x�n�I,y9�uӒ�&�w�D�R%wn��KzKM_���8)S�J5��Ԡ��j����ze�v���&5%,���9���=�	��|�FBG�y�qL�*����˞�>W��$I�_�t	�ub��,� y<&p�-q:��@���]��֞�����k7����sss�|ee�֭[W�^e���g=��}���U)a��W�4Μ9��]������1�1�2޲/�>d��&��Qv��-<X����r�2,��c�!��a��<Zʾ���7�4b?���?3;Eھ�-M)�\�#�i�rJ��a��h�e\J��<���߅?)<6X�2�P�{��%l�s�.2� �,�"�z������0!�e�t��AEϭ����x���v:�+��~jqq��^~&�D0��&�(T�+e�)D�E	F2bP�I;i��� ��lqV���4n�X��qc�au[@)�W��.I�6�Z,�9�x��;���3�����Ndp��w�}�qsy��5�4ҜtI)'��O��>�M��I �Q�*�����Y,L�(�f�R;��C��F�U�����B=.y��F�X=���I\,�<ԝrV)��dc�S?}�,ڭ�5��q�	��޻`�� �t�R��4R鵤��,*�4"��UK�;��kIuG1�*U���bRZ�"��⢊}��~Ƴ4�w#��$��7���_<�Pb)�[�KKK�Bզ-U�/]z����m�.Gnױ�bVTqh�vzr��_��q�k��?��Ѳ[��&&�ή�/޹x����{�oMOOY�����ˇ=��k������I'	%�l���8��L�&������z����ׯ_�ֿ��L��e�ˎ���K=��K��ҽU�L��]4슳�I��Ek(��΃�+Q)W�Vw��.��u�����lS<�Ydh,`�)Ȥa�m�ʵE�j���a����w4�H�����^{��(�0��}������=s���V*>���S�r�6v��O�toi�֭�{f�ao	k#�b?��x�R�D���(�P����rh��bO/퉤	Ixėh���x]���{͋�-Bq�����^�����eF������3�������ohϽ�&~:}����8��~��ۯ��;�S1Ǖ��������b\~��\�X%�/rݬ����V���V�K�
)��'$ ��<qo~�ր�5��?rNJ�V�ev;b��Ә�ڄxG�$EGga*�8�#]��N;���CGA$Y�I�;�s�����Ii�`��kT�u���〚@_���"ݸ"���T��Rg~�G0�VV�W~c���p1
�g?���1����������q�n�s��g��mT��/~��_��'� ����Ç�{��$*\Z��jIZ��{���to�}l��,��eFf[��H����(T�@�2[�tD�4ED�$ĥ�2��A�
�%�m�����a�a���k˰�}e ��)'���\R�}D��W�飝~^��/.����Ę�ҿ���0 �}��PzL�G.w�U6q��X6P:2���b��U��_���������d��źRM�:=311��#?=66�;�ݵ啕�.�0@�ʶL[�}q�����x>�H�jR���8��(Q����1d��Ĕt!����A 1�"��pc�B�D�Fǟz��9"wޫ��7���@/����$�B#���s�C3ǎ;|�NXx�뛫����8����	n�D�-�,m�N�Q�W.l�5��h�#f_���I�Jil�sv��7)�����"���T�Ԝo��bG�b�w�|;$/%���=��s��w&VLOa&獠��hs�'�U<)�x����/*!Q%�X��q����t��Q�V�&/�9�.K�Q���'8]DQ��L3N���V,����'�u�����ɳ�I�Q"�rq3�1=%�ڑ�/C�\/ �ӧك�����Ÿ��8��<��|�G1�{�a��5�=C[U�U�{'Wٻ�I>h���i�4��f�Z;�D|i�ifre�%���Bx�y��?��>"��v5�%܌�o��*3O?�����W�766X���͠����ˌ>L�'Np��7����O/�Y���/��S��Mk3��$�(�0e��m���ޏ��~�:0��_'����Bԟ����5�G/�B"�I���gͮ8����؀d�&�4��Ӳ3_+�ݺ���y��o|����a�6Dyz��53�-�]Cæ	�	 N@\�,�VM7??�̙���7�8���}���t� Z��Śo8����r��j��+�Df�`L�'��ј_f�2�b�~�����|?&����VB1,�2,��2�Z�2,Rr���X
�N^��l��j�,�F�ᔕ�ETT�������f�k��0%M�A� ��k���]�3���W>������I��E��i���ҳ���!3�EϤ�T֓)������'2�VA�ƼTk�]K~ФV���j�����zP,�6��o��U��������/y�v�'�����w�,�Ɯ��.�|��WVnn�~�H�f��FS�4v5�ƹ�01��A;�=�:���wM�<v��~�?õ����/�0�5��BK����y$�	���f��.�7~�_�,-e|�_�»[�0z���9q�I�)R�V����+���N#�)BM7�?�L�����jsz�X����:e�Qeqq��y��e�6vln��~�n����Ǭ"Ť1�|���C$�6�������Ъ���I�*�O5H�7����L_��T������j��^���O�.�����[�sQ�֬$��0B%��S5��F�4�;��ׯ�r	m�H�Zс1�8a���;�nW4�L%ѲЮ�ۭ���O>r�� �"7>�r��f���Xՙ�lo4BwB�Mm����{k1e���ݖ����3���Ҙʪ�Y�&L��#�cңFP
F�����������+"��z[��^ٰ��g>��۰Y�c����M��1� ��1��vm~~������Is�nT
v^�0�J2�L� 1�4�Y��%E�
ݰ�]��]U��>�ʟ�ԧډ���#�S�ot�:�[x��b *���5���dK$0�hY��E�d��$0�H�H$2�V���.�fA��Xu�����v����J��]z���KG��N�9u�����.���	��0-��_��8z�:��iY���?�7h)���(����;�͎�_�]/���Z�Ly��_����q��L� dh�dm�n#ZR=����K'>�n(C&�	��t7O�nF1��j*��*�������&����,f�Ha���������)_K��5̋0'ȡ1�6�0�G(�!P�q���� a����	Ü���%ػ�����S�\�q�撡j���w._������?���o��KW>��_���Y[�`ByT��/ �Ya$|�K_ª27��130���J���Ï�ON8�*����4u�xR3�������(U�������>������?K�<��}�yu@x���y���i��eX��Q�XkX��G-�7����ۤ�����YF6�~��"'C��_x�&���]���yM~ k��-ː�Z䲐�Dɭi��fN��B=�� &7�#�ܥ�/���\���࿌�p2Y��fuC�KKKh�{�2y,����{���8�R��TG���)��q�_=E�|��X��k<�d��p~~^��T���$U��*��
x��q ���������� ����UtB�E	�����9@|ߕ�o��ՄYD|��x�,��1ZCc���A�9ʭ/p	S2�Gq��r�.-���^�	���s��(k+�2�J��noo������(p�S��m�&l���q��J�/����8�ȏwy�_�DQ���/�}"�V�Ώ�{�
�i����ѣG�[hsI#A%~��^�W�2�ٽu�kd�*̓v��%����6��$� ����)}�Kfq$����#�(�F��q���gkҾ���U�.��47s��)�4��8�V'^o�>T�i�uٔ�r��[����<�ݡ䤍{�j�F�(b#�
��>k�U��8i��WX-a�-hX�����<��"�&ե�K�`B����K5���Aޣ�dg'pc�O����g4
e)Js{;!�~?NbX�8 �E�G�.?Km�����Z��E:��~�-��SJC��\#�>��_'Ke�,�l�˖7�|o|��;��-g���ϳs��I:fa�~����xR��z��>�Fơ�<�8��N:�8p�/�|��_0�=�����	Lp����@X8��}�c���k���I��s��*X|�����ߔJ%L�TJ;]�vpV.u�pL����>���c�����m�a]��yG�w[8Ox߹m��|�1��[|�n�?��}X�GB�����?oư��e���eX>P��%%��9hǴ�Bq�s�=7aJ�0�u���*��ݬ�Ǚ��.7
{�)�8|�/4ɥ�J�'�/�A��~�O���0	�_'l����5�A��*о���H*J%�b6�a�J[*=0�d���?%fmUp !��Oa�jz�j�f�ձخ����j�"����t�+W�,3���Z_]i�K����^�{�֔Y�]�J2JU�)�Om�S��v�풺�&�S]�U�'�e[QF�9����JJD�ɑ�xYֆ�mY�e�%�4�-�/��zuu��ލ�L%^�ݨ�Q���,�q(f�j�8�43U���nh��hco|��X�6�[��v��a�9%�P��̬RF����|3-R8M$��Pz6:������+aYx _��R�(u��n�/��ƥ�v�0ձcǢ���d�^|���z��M�O:"m�X�E�Z7<�Xܖ���EG��=�74��B
�n�DFh��02:�z�����X'�z�fۭ�,��V��~5W5EW��%�ʍeԶ��	�kIЍ̌H�q�))+ޒ�h��Q��:0gF��8K�0��TS�8Tt�z��Q���(�馩�׎���n�փ&�-�ۉ A`�
�;Ԟ	��D5#���ղ߶�K���q3���Z���C�rQ�j�DӢ4�l]�l/�r�����.$ɑ#Gz��S4��Z�r�<�F�W���-cYMrr	��"Ԕ�5i�&�1t�n&�5]�5(��a�*�P�����q��-��$�LA�����L|���'50]�5#q�f����{�QK�N^�B��&��o��ac#h�PY��h'p�B`���I �RFV�s0𯯷��1�rm�i��ٖ�h���O��,�jY�����3�HnK��ꁱ�c�^�JDy���%$�i�d������{��JO��G�#Wc�byeL�A�^(���z�-09>566Q����OR��:�(+����S*;q��kkk���
j~衇0r:����X���:���=��o:A״z��_G�'�d�$�!�@�_�����T%R��Q�Z�K-�\*�ϲ��wz���DBrJ�7 �2��DU�w�H�m�%��!�o9P�!C�ˇ�!��a�aE��nBz�;���z�N�'#U��ą�X%oh��HD??�n�\O��K��(��������;��4"z����7d��&�#�c��xê5��e� ��}(��.1>�V��`"��3p����ކ��8���J���򗿌�<�NI;�f�9nS����CDj���K����9t�%��v�W�zׅ���p|/-DH ,}q�����r����P,$�t��<#�)�=XT�umk{vv��ųz��U�- ? �$ű��+����Fݕ����[�V�����Q���cn��������d�T�ヨ�>�e#R�����pJ!��&i:'l���SONN��-Sn�Cm���AN��v��;)M�Hr��]4Ξ�L��v�b�\� t���2'�@����6����6#�{O���r�J$�$�ѳwQ�/����O|Mz������o�I8==�D�s��@�/�s�"c�Ԋ9��n�wN���7�/^��P�W7�T:���n�N-�n1�# z��vdCKnIX��DlE�-��16�Ia�%��"��(OH�@��0����{��o~�C�t�̿v�Z�G���(���z��kj�Q2j���C�3:����LF�)��i�1n�RV��M$1Jccc�2�a�KK+n�|27n�8{����#>�`+�ϟ?�mw��xF<i y5AI��"���>q6j2�O�u|��a�v�h��K���՛�L�y5��}���Z�F��~p�7Ve贺?�f�����?[.�@��yD�a�5���o���\i�FLNHN���H.�'�q����H<����)X:(�O�7�/��@�,\-�4������p����=&�@s	�$������w�}?�S?��������/�_>�쳘����h��{��GCAh���/|�DoC�,���Ǔ���^�)��z���jr�K�g���v�T�2���T{X��Ud2Z��Uq��e�R%��gp4�O�ZCgװ�,C�5,��!E��ʠ�Ib�X�:Q܂!��V,u9U�M�q�iD���)�T��A#�i���x���P�>�S�9�{w'"�'���&MM�����ɼ-E����0'��>�V�|qK�0�2��>��3]�?��`I2�A2M��F�7��$U��t�L�J1ɳ���f��떩�Z\,��%���ȱSMxa���]��7w�8��D�J���re�6��f��/Wv�0�,Qd�	�� KL d%�vL�b([�:[cd�����~�/�aw�^����L|��j�Q�kI��"��\J-�M�0Jw�Dъ�jm�ފq�k��<�նH��n��Ԅ	\�$�3�����q�	aW�I?���_�f����'N��;�vŨ(q<�(j��~7q������������{�����:	!3�gG����a:��>���}5�5Q(�(v+��\X5��v��
��JX5-��#�x����r[�n�X��,�$��������{�����Mj�LU4t�E�ȗ�)�B��H	�줆y�z�V���V7���䘫���\j�F����7�u���H+z�b�m�y��b���\,�X�Y�<�-W4W�N��8�9Q1�����b5�Z{����
)q[F�*v�ؙ]�۾p�"�B$�;�s��a�a䚥�Q��8����b�q�I1t���>^|�gi�_;��IM�g�4Pg ^i7�,�M#5r��0�GV;�F���޳�ŻO'q�kV�HՒ�K$�f�@ݹ���'1wh,i�iXfNC�b�TEw�s��MgDpت�I�Zq�,C5�$X�	��m��C�'E�JD$}&�n�,{E�Z毧o�qƑ!g=&]�+�%�^�bz��K9����䢑���^}IG����GĂ5�	�*J�^���x��qVh`BB&ygl��Ġ��%xӁ$�d�3�0�!/�-�٘/D(���n� �� c^�j�����E�"�Z*K�n`�8yqoo��B����`��:c�'z�3C�L;�ZKl�&~N,4擘�҃h�^\ �w*=4����>�m�F�z}���9uCvj(;v��a���k˰�}EQdF>�+���V��K�9�����-@1rD�E�TR`	�/�����9^����� ��w�2j� A"6_}�9����߈����iV��BY8�-�<~�u[c�Q��� � ���.�������D� $8扏=633s��y�yg���nm����<y���a��ܸ�w�ى'"�8w�\}m���%S"sHrJ��ItMA8�2I�6��0V��Í(ۊ��0}��5R�2I�jes��N�Fq�K�T����t�2T�� �dԢ155U96��)?�wvvο����Ҹ���毿��������ewD���T�qIv�T9Ha?0���M�?�U��T����|�,Tpu�.������.�{�=w�ygM����/�)Uu�,����?��#O�>��y��w�����
����MT�Z��������O?}z���/�|��wpK���ß����g��oj�<s�̉C�ўWn��{�;�0==m����_�z������j���*�ɋG��?���뗿��o�]��y^@��Ey��Dq�zm�L���Zx�RB���hP�	Y�y�a�������&�A*RHQ2���s�������)N2��FSR���V��#�Hl7ɛ*��m�ޙA7y�=�������;xRW'�UЮc܎Y�����~f�
޽�D�YK�H�PEp)�^1Bɏo��T�.^�H�g����92R}�ӟ&���.��ƕ>�<q��g�5e�Y�X�94ɖL}rS�/�t {'O����7�]���7�1??xd
w�x�d�"�D�(2�9�{V��F�*��S��1����XM�K�O-���s��A�o`�?GdeJ)q�^�2f8S2NKØ)I���]��AOaR���Ǐcb� �`Xr���7�A��ˊ$fD��0�0�pch�KW�\Aa$lll��eT�!��C=��� 
�ߠ\��s��p�v�W^y��6|������;O�����Vt���o���]�-����/6w�1�~�S��U�`����	�g����ϲ���1�� [�2��<��%z/)��˰ˏ^�XkX�E��eI5��wy�fd��
ɌR�������릎g�cST�(���iӻ\d�*����$9�圶��Vo&M�#���'��~O�`4Mbi2���o;S ��?�{}��c�r��V�4
u�-���O��x��F�$��t�2t�$�0�Lֆ�HV��E�NR2(��"��:�[�#3G�bs�%�"Va��giB��~��N���_�;|�pm|�	̽��w:��Ҹ:Z��ƗS��c��M���_�X74X��n��o����4�A��N/!o�cqde��i�^K4�,�YL���T�̲eW��r-�.�-��~djr�\��B[�<����\3G���t���k�xqzld|d|j|�ըD%�\l��j'�J��+�� ��q��h *��
+)QF��T�O���$��C�,3|<��DH�@�,V��Ov�He(3�#b�����(�-�S��B6A��G���s0��ɽ�x2},��6���Ԝ�C�st��GC���x��ʍ+�4j��]���f�Kc�����lk�6^������7$�}��u7_��fԜ��1a��/X���C��OW� ����x������n�W'&�Çr�Dσ�kMN�q���n��n�cձ�)��|����8�z2!V�H	�8.��6��VJxlub
vmB�i��iOu�WMS�2��Zi��)2g-�1-�nݺ��\2���¡����=9S���_�^���զf���
��hI'IʡJ�����ak%"��-��hn�{��E�0��5��#,�#�M`�ꔋZ$��Rڜ0
�EJʅ��!I,CŲ�J��Y��Bё��'窦�nLn.9fR��B�9�L-�k#s��V��N7���ѩ�X�~�:�ɘ�Idf!�@�<�f��hB�Y�d���������tu�˜Y���Sr�MB&Z.��$�TuR��Q;6+�f�SJ��hE��V�u�#ݠy`j��~�)Xs�$L��(�����H{c��X���$�Y����D>@R�q�Z�<�ni}}��id��&�\;��>��;��� FRc�*�n�[������E��Na�u���g�yƐQ�X'��V�����W/wows��r�mR)m`�v������g&;���޶�+$=�,VU�T�T�x�������DWT��3�G*R� ��	��棧��(TQ�X���)`�����hIO��_���E�&�E=�o��a���k˰|x�yU$��0���Bŗ�rm7ҙ���wzzڰ�C��zRۇr�'G��F;���[پBW�_�� ��][������ܰ2� ��� ������f��� �o�y�ms.�`��K�ѐ�Cq2MV��^��S�(�|��/�r��e�B|��gh˹B�%���7�^�r�ʴ�<��Q�C9�"_[[;������܏��2�gqq�tlrbd�Z���{��]j�d����~����qLi��"�42Po��C1`):�J�|�����ԬV�%������P2��a�O�ig=�*���~����Z$�[��8�Σǿ��/7�ܤ�H��ׯϚ*�������? �w��U�T�p�"[զ��n����7/ݸp�B��Y����<Ξ=�<Z��0����_�y�&�M���c|�7�#Ye������;i�	��	��?��?��Cc���o^]Z��t���]�T��&
䩐N��g�WѶ�R��I|R7>�я���t��W�����R!�HA[7M~��~�я>�}M���ӧ?���0&L}ee��͍|pqa��vk���������Vkuw.^��y�2�_�:��'�8��i��&'E����_x�u�C��j����q���4E��[���;Ͽ��&���ɩ�����7*�w�kyy����u�ԉ�_~y�����1M��'���?��'�'6R���R^�H��s�y�{�ϟ��ő�tq.��~���<���ӳS��h�D�M��J�8�ݟ��������O:�����ku��A�b�^@�g�E��2�NS�=	4m�@>:��@I�q�$�		0����)�N)*3�~*��y3(t׳�����	1��XY��7��JY���$!�b	��L�Q���`��;�-E�)�b9�;M��^x#
cW� {��W�>��Ͽ��w�J������C����>��_��_���1���N�:��q����_��_��w1w�{｟���{��_z�%4��wߍ�Q����(~E=����P���}����k����q"��ܹso�����є��?��CgΜ�v�֍7�
\Ĥ����
�-0��ƴ"~ ��H[�)j�LI���9T��)���e�G�eo1��W������a�@b�a�)�(����X2�B�q�R�I/(��4)�<N�j�"�
�X��b��RK��0��0�8$��ȥ�T&�����7zd������c6վ�����5�"�{ɲwHx�N��ΙF�[e�$����	��ni9Q��H�T�� �7�D$r�VQJ��~��핍�����q6;7~ǉþ�R��nl��쮛��p�1�Z�8#j��[��LY-;���i�5�)hcy����@���]�.$	uZ?�I--O�����IDQ[�F!��ȣ4��h��8�F��]\8>9&,�b�
�m�6/�S���D	�R۲�p
������4	
kJ�T�=<;�n)�4;��8��ő�qE^�Ԙ��Nr�	����mrNO��Xiq�D��i��jW]K[�7��z����V=ދ=�h&�����ӳ^�W��8�|�z86٤^�+v�\�������4_[ۆ)�^R���d���;�~ֲI`�K;MW��c��Mg��'�U�O 05#����EL'��d�ӥaM������c?�4
hV%�J(�QW�̶ɳ��r�h�����Lu)�^�©�r}��ꌘ�Qw�[��5%/�T���Q�_�o��gjF��(���� �Զ�[egS�Dyt��w��E�*x"�E~�-Xj��n5as[��Ju��T�(����ʖv��S3��Dia��K���Hqrs\�y~;ȣ�S,�O;q"�Di���P.	]�0e5Qr�䘹�L1t&�Ir��"J�<cu�;�<Y�Ug'�M��Gi�cW�,iu�VPjerRmd~�3���Υ��ɴpi���h�B�D�ҩ�r�3��F�4������-��3C5&+]ST�`,��8W�H�Y��s�[��(�#�q+#S���'��4�1V���n�|�תfXDKzs3�Y*%Y	w��j�����ZqL�)Ӣ�L��!�n��+@�c�ngc{���X%Y����Ĳ�����OLL\�rm}����/,��^�����kjj�q(��N���.�쓜�Լ:4����!% ���~�+N$aI.����}luu�q8���rۢ��\;�x|sU6M�t]����$��ب8���kV+#�R%�('�@h�`]�Q�(X��GQ��DK�����Z���%�=g�h]��Cq������K1,�2,?Nb�a�)�����}mm�h�|�4eO�C���N��g�n���HB/c���gaL�Ȓ��:X���OH�G��X?J~��� ����qe?���m��|�Ş�T�n���e�,��1����u�/7�U�͞K�fU��F�p����緶�`��rO=�L���j�U��K_��իhfj�Ȯ,�cFF����(�؄���4p��E?�[۔��$�5iH�٣�df�/��Edpc�'���(>���G>�U����;N��Z�ڞ���0�Lx�ȑ�~��t�ׯ_�vա�����YY[A��GR���K���M��-���Շ�����p���)"�k�`���*N�B+9�
��2����6Q����F�]�z�"5�<��|h:���7o��P�]��I��`�	�TqCq�������>����w(���-8��.��ȏ�k׮� ��D�V	?��Fm�!���[�2.1j`�Kج�eq'��G'��]��*b(�������tF�챌9�hg��y�Pa�5�.�i"�����h)0
��щk�%�┺V2����)�D�Q���J͢l.԰����ډ'ІG��c��o�&eOQ�h��c�:ɷ#[�`�<�(�X��<k�z`���[��)�1�6�T�z~=�s�8�ڕaP��dyyC���
�����CH�R�'3Ns��N�bBV�
y�w��+t���?�(��X@���$�!{�:?X1�@bϾL������ w1�̐��h��m��?�e�/�я8ࡎ�_��q��n�>��6s��_���-3���bay�����_�":722�c��U'''1�wvv8h��h
��G�KKK�>�(�����j��p]t2��5Z���1YK����Ɵ Z{D�h����رc��w܁�ǉ�2���������y����k����>p�'>�	t�<�@��ܧ�R�QH;>����Ų���������
�6�Kq��b6������eX��-C�5,���� �b�_��q�Y�{�P��`vv���(�q�%�G	3xn ;;�3�_a��^�+oM|���C�}�h`��a�
�_u��_��>X(�n?{���eR?�{�WM��x��RTEf_(6i�Ā<�u��2��)��,OR%��(1ʾ @Kz1�d�R�*�t`̤m`2���)̊�0�4W����jJV�u����w`�h���S�W/Zjt����_�(���i|����&��~����#i���wqp��o������蔙��IM7�8͒�2:v�=�q����f��L��s:������^�4p��kv[�����ۨo�w�VH�]ur��^�:yϣ���ߐ���R���&��$�ݽ�o}�9��N�%�0&^�z��׶6�Z�J���7$�gA�
��f�n�ɳ����2����tS�6|��0�b(@k��f})ln���٠aJ����15$�9��TOW�����4�r?"��P�B�%)w[Ġ�m�J��X:Q��1� j�B5R�������K��(tn��F��U5�×��o0�n5v�>��]@����������R�1��E�nUM�f���R[��P[S����=�w�dT���#cc��\۩�S�_뺥Jݎ����6.nh
ϸ'�V�-�'f�ZZ�����ŎJ&�=V�r�+��[ϣ�:QB�s��v�ժ��a��\��/���&��P]���ĝ(&E�Y�ّ�n��ግU��^~�۴q�v��%�QE��i���Gˮ�����'�|>X�,'�9Lwը��7���W_Y^]���%�(�F(���2�?O�4�u\��w�ƭ6��TwI�Q�"����D�N�̐$52>�DS�1!��I�y<��]툲|�IR+S��5�n�s	���#dP�4�
����J�9�Y���!��-M��[�CĊ�(�WIY�C=%��<�)�3Q���)�XnP���>MSL�S��@]I���$�-Uׁ6�$���Nc���ZŲ�x�o߿x	���;0b����3�ɏ>�qz��z���������F��=�Vധ�~��G��d��?�����|k�T; ��>�q�0"RR�g�y#$�s���_ ���w ��+�lnN������>}�СC�8sssx_ _�}�c}
s�Yo�~sƢ��v�T]53p=���&�0ڳ��Y4USd:WF�K��T�� ���-d��#�)�eX�凔!��a��2�F�gU��-a,�| �&�{���kEՑ^��YX\\����[��ŉ��
��W��7:��p���Z��t���>��s�#��*��h�}N��%k���o�hQHB<�Qf�P�����y�n"��5ކǑ��̆�<�1��o�a�M�R�
�����R`ȣR*�������,L���Ky�Y�YX�p�7�+���;�0��\�R4
�Z�fw���E{�ҏQ�Y'O�|��ǙUX�Omd��fc���ξ���d���se���B��!������e�M�݆�5??�YN�T��j�����\��������/�������;)%'���g����.�*��Ƴ9i�m��:��13[��C�HתYe!2Xo��8rcc���&շ5���(%O%	)Ɏ#T�	�!�
������:1©�D�_���Ap.��P��ŋa��� ���F���5hF�j��bo���׍����ϋI���n��	K���c�+�{�ƍ�:��S��ʢ���ɗ��;���	L9he��|La
��-Z�����aw
�YV�h�����ׯ�<��#��v]N���QI���n鮻�B��^2%H�k�`��W.\�E���}D,MK.Ӑ1�{�>��O5Z��Iw�f٨eu�/ڑE���g�w7�����Z㹿�ȹ)ľ��CMWg���v�+y������<Er�h�����3����TU����S��A����=����`UTƼ��'�
��INEX�v�MG�����Cq���DV�E���|�6��[o���o��o�7��h�3g��HV����=���_��P�0��u1Y\�����a����v����ijb�5�ĲSĵX��)C1*���X��b���9�'��Mʑ���'�Vhkߣ�����=��x����-<^��k��u~㨚d��zojO����M| g�˰�?��ְˇ�~\O�E".�#�*1�۰<F��N�M�d��w*l&S7�(>�x�/�v�%�E�C!+iw�6ޑ����q�FZI
����:��b`#�|Kl��R�4�Tl��\0����|�T�8EF����o(KPw���fkv|���ɞn7��b��hRr��>Gk4�Mʎ*���F:c��z��\%6�z���;�a"tB_N��}�Lw� T[ĝ=:����/��n�ַ��=^�M�0;�M���C�㘕�om]2�-�%Kٔ�f�l�q
�N�Y߄Y���mvI�T���L9V��w�=�;���<M?w�>?�3?]�����;ϧ0���~g��q�J�������;>3�So�������u�����{챙�C�cE��N�.L��5���^��;�l����N��P6Q��[���:�?���"*O��X�^Ci�jJ��L�n�b&$��_+�B���!vӠ�����^�v|�0�O�3��v`�$����Dj��i��E2%D_H�8i�>��$�b��0�	ң�a>��{ݽZe�K�ƅB%�,�j��� ^ȺI.#�t5S�����Vw�,�~�hʑ;Nmnm�:W��w�#�&mF�� 8(�J~�yH�T��(4 /�����W��P!��������W[��DM/�����*��^g�4<C'�TO�EX�#z�R��u��V3�h�ە*!�B��$ݥ<�+#-�1�k���m�z&�e�i�6ڭ(H^��kv�\�ծ��/��6��[���y��R���������g�'g֛b��{�X��8q7���FA8�C8�h'B5-&�d�q���ڑ���<�X
���#ggy�fb�%�T���f���� %�!p��GHI-[�������n�%N5��$7�,O�$J�<��b؊m��jRз�h��m�Q�� k��t_���c��Ð�>3��lS4{@�NjOq�iF�E�i�<�x��)vI���W"�:�F�w��J.���O�i �ħ-�T]]Y:��v� ������w<��w�u��Z�g`h��l<����c�a=�,{���@O��񫼫���W��1�;z('Zuvf��P�͉���j7?7�+�e��Ѿ�*��*G�b(�l<!�U�rѲ�1	H �T��,��pcN��q�%{�Ԇ��j�/����f�A�QQ
�G"�H��)I��4�?�ib��VI���2�j��c��b`GO�=4��>`F˰�Xe���eX>����%�b�@fc�b���搷WU)�"�V"� ��>��1��O�Y��8�PȽ侰�rW��c��:d���I���o�^��O��3.zm����f�{���vjgs���8G����Yh0"��i�\/�2#�Z��v{�n�v'�L�{'�O9�g�ϔ$�(=?�4YҜ����%;)���"!���0��|bC���@�S�Bw�C��0�p���waۥ�C��]�k~��!��!7ԉ�O��0��e�+¢������o|��Z�g���ܬ��)'��WVV����G�^�v�����
#���}zi��I����R��b�p�%~��:�֓8#D� A�:����I<�Q��Fݗ@c���{��<����ض��&�ō[��p0�"7�� �\�0�Jpd�X G�ܭ����߹�4�M��b�Y"�.�}�Ș۠������?�V�Uڡ�G<�Fye-�f�>{���x3������.�Iˣ�b����V)V�0�IM�g��J�Z��C:i<x��b;v9��d-U�h�R�2�p�������X=D�vF�f����Լ�F��>���g>�|_N�
�������j?u����$����ɬ���M��/(�����ޚ�&5O1�Xfi+���?c�8�$Gb��[>�@��n�r23?��_��`Vz�}��R�$l�O��s�-�w!��w���D~_Y3����>zfzzzk���R)����)˴dBio�xP�"ý���<�{3Q.}�n���r�m�m"��1O^V���;�M�9�LHˏO�"}���=�C=&o���*�c�UH7RT���}�UH�$��R�]F�2ӢUˈv�CEt�\S�&~��@�d�+�2,�?+C�5,��!���6
�Ma�۷X*�?f����T�������,Ls��`�U*%�J\��ua��(���HZZ9g`��%;�����fR{�BŤ��f��ɌL[ﮛK�2Vn�I����A#���v��~`9�<d.>s�	ES��V�t~��"��f�T�4I�G~�2=E�U^$YC�Lq᷾��B�l�4�����O� q���K:��VS%���l>�PBύèV��k��-��/VtXR&�'�]��9��}��Ĩ����˴�B:�e��&���#S��'&�bi��]h䉹9�,��h��}�b�Jm�����}�T)s�E�0u��0�P����\�(�>ۙ�;jwۍ_�th��<�3?�킭:�uO�m{ΦP�w�{��I���ui�ed`�[`��Mô��r��;��<Xjh�p`�e���f�[I��̨o�k��-]�d�F�P�*�dw�d�*%vh�A���H�J�$s����h��H!M5UĹ���GI��ui���F�
��U/�;�Wic6e��˒�N7�]�'�!�B�ǔ�U�Ո���]�u�ݬ`
)Y�{�_��H(m�4�gIqv؇������T�ʧh�A{M�B������Р����S��M�OP��L��F�3s���n��R.�8z���jm�L����bM��n�j�f)�Y(����t�g	4=�H�����"x�u'F�<��g���0eLJ�±���Ԝք,H��r�	���[��i���8B�7}��Jr"u'��G@P�P���\ѡp;�r�a1�3�Sɭ�RT?�4��1>MM�����p�y-Dy�{d�KId6����1a=�t�Z��&�\I2H<��P�p�x �<��/<v�q��^��h�e@�k#c�b���a�E�VSm�Rn�n�ڽ�=`%��y�چ��L�{*�p����>�l�'��؀y��`���Z/�+�t%4Ci��Ms-$jź�K]E�W%�\� A��≤)qܕ�!tES��3�����@�`���j��%C&�o�&���F{F"Q���󈞙�S�I�!�\����<�1c� ��μ��k�&�I����%W�Х5,��c�!��a�������(�{d=<k{gkf6�0�c��|����_�)�.�w�'���A	f�S6�N�>sF>�5Dۜ�
S�����C��2��	6B�����X��8趄����mʼ#\���Ô���(��Sr���p:��/��/L.�S�}����l�������`���ͼ�꫑���O=�Թ���$m]+d.�(,LR���=B�~H>���طC��B�ϘԼ�����_'D�]�T�☢і�Ϝ9��Ϣ~���~��GQۭ�Px �;��Y����}8�6����	�9u�T�h����v}cc��
��̈́"�F
ţG�.,,�ڦ *))�ID�,ݝ�1�o�W��9��h�$7]�< Q�^K�J��W�;<�ؕ!�w��� �2? C�(�ڞ���(�4+��w��H��5��Q��S�h_:�Uɮ)�A���?z�ZVM�E����Z���1h����j3�S8ҍ}rܤD�h�6ZO�)�4�N�T�ڄ���qƎb���N�F2I��
ys&^ɳ��D��n���*E��IQd2�cʧ$����p�&6,Wܰ��B��K`�����������0���aChfj=��߽�������O>Mq�y˛+�h���齽= <c�e!�t;jD����^�k_�ښ���`�&�����W��&�Cp�c��q�>$�N�B�ϖŬzsss<0aQ���Q�i�aw6��B-/��q@%%�;�|���@ˎ�~�9��������gva)�S��:u=c��`:+;���A��4��[E�^�2f�F�� 1�	R�{� ]�D�g���s��F��>al�nd���o��x�=�f�x g����Z��o��|��z��(
w�9�<z樂k��U��?z�I�_���lMZ�����R��ҾϰX�/H�E��0~�*������eX����ְ��_،��8%O�PW�Y�2!8�n!���r吪�SLc�+���\�O̬S���3;�,�M
�<D�2l�2�eml[sm���8�Wx�E����ȃD�i��{Ma�bJ8ۍ�-�`a�����LQ�П���~���Qx[ƺ��{ WϿ�*����������Ǐ]��@-V�S�c��b�J$�0�8���;)�u
|	��TRJ�U-N�@�UCw��=�`�YG�ӂ�)%���t3d�J)^�F��� @E|�R(:k0��{ϸzV��ׁ���������*f��:��d�T���Yz�])�ŒxYS��IX�s�jä��7����;jNq~~~tl,�"��`,�YoLON��H��P�*7�Y�H�䮷���IqW�6�i�ŁDn6��4���)�<-�QwO�(Ո�-RR\ 2r����ޤY��:�>{�o�r��*���& e@�n��	�ڌ;-h2�I�ߠU��BZȸ��E
�6��4 �B��5�Y9�|�s��~u�s��E�@ Zĵ�ëx����;�9�i�@�Y���6�l��TE!�DH��(���:e�2ǧ�2<�&q���NZ��f��l����?2i�ZYJ(�6hb̺��"�h;�O<������^{g�a�Vj\ظ����ͻP�0s�1��8���#M��Lâ;Ȑ�G��%\@��2#M�%�U3	�Ďu<(�q��э\�m���&Q�ٳ��S�l��'R��16㈽!�QD�	�N��p�+��h����I�|��1p���9��o}|��(��oaa��v����&�$]?�VZ���vg �����`}e1Kǖ���B�k�v�Y[^����W�����E)��Sg�?:���蕹���z�GopL���EI"Ul�d�C�euu��!-I�k�Iި{�K� %�h)#G-,��ET���<Gu��,l{.ͼE T�ۊ�
:����	����G��5lE���}T�+���v\�:����,��洣���40-���'��	�����DO� L�<�ќe�g�[��ʏh_��,�{�{\�b��YDh_7��t$���`-�E��+�%�p,�	���r)�*�G�҃C.+�K�t�ә�Z���JzE��D�<vIP�l�0�HI��'�3�2t3�8F���z��E�R�M7�6�tj�0�!E��6%�d��p�/��-�Bgm�f�Wj3�5k���M�
{FYe��0Ix�Fv������=ꖗ�{�{��EEͥK��|��N��n�oܸ�8�~nn�>��;�Hn�$��#\�@�34�.%U�@ձ"Ծ�g��CP��<���Ͽ(�$D�z�K9#2/.]����N���	$���.e|�~�F�t?�^������GGG4b�����������
��O\�i�h4�`��t�u�������r}�@��I����@ ����]���x|�s��$H����M�.�nB��t�֭��}�Nv�U����o�I`�1p���`p�u��f�K����ߧ�ppء�ɪ!|~�{�����%�W�^=��JVr8ӽ��9�u$5_`�i~�r��!V�c9tw}%�d���h��� �HX���T��u�M7$��:Yl�zS���8��^q�B*S�����ɘD�R�D�����l. F8eW�����y������X5\T��l�������,��?��{1�B$�!Wc5m�;�~�Hy�nG\J��4���ހ�(��+� +*.��F��$=�)�
���dzl�$V���ʹ��֡�B���5�A��<8<<��3�p�ŋi��:��]���3���7��!-���卍՜��	U.s�n����Y�9�Q�W���E#CW�s_'\����%h�Q�����F��g����v��P���흊)"x�А�����ׯ_o$`b���t��?ͽ���1^(��ĝ�(�k�'|��/T�^8�Wg65a-�G����
��]:���b���Y��3�:� ;n��RS�ZE^I�@q 3�˴�
���-����LZ۴*H&��,�
w��Ë�TA���O���꩔B;$�&	f���)�xg{�~����O� �h��:����i��|go�``[�<&*�b$5���Y���֚�Y��V=b���R�U��c6���hA�
�d]I �����v��7�qH��P:dW�� r��ZyOU�%�ZՓ* ��a0�J��3XbY@�cB]��UȊf�\���(�B��$
|�:ݮ��/\�@wD�+��`��7�'��={�Fn��q��oy� �tj}qmqcmqee��iQ��f�QE�g�L-$��=ڧΜ��D�Fc�F��`G��d��ۭ��r��^�ȣ�b�A	;��8�Ƣ��.�<�F���,�G�c�Z��idkuieqq�g�r8�_�뭽��3:�kl�:5��=��9�:����q����X=}���!�p�����q��:w�l��N�����NïY�+#�����R9��J�6��<pA�b{m~>�s	��
��CȎ'�5�sd �Rd�2t
�K�>3�� �~H�P��� ��,K`$�ҨσbH�H���+1ѫD[ȯ�Xc��	|��_�3�r�u���F-�<gya@_�K�.~@�,	}ϝ��--�xB�#��I�"ΌL7�um[���Vѝ8��FcGcy�$u����{A] Ije\�6�PwH?��ю��^�k��N���f%�$Ef������n�!CHWJh�޹��(K��,-�{p?3ӻ���9�Y���$4�\T�P�������7
�t��4f:E�Dy����}lF�6� ��|n ^W�7�N�>Dr�!X���ĭ\�QhQ�F�y��:�����~f�$��2�Ԇ�lp��
��׎�S�N�F`/��q�����B�b#�T���M"�ʮ"�V��	�B��\B�Q1����KM�t��e�?v`݂$E��:��D
�N��w�,ZY��}G���h.� �|V�1�O��K�A��G�k�X�U��ꬖ�F����}O��&�m���(�ʗ��	��88����4���ta)��v�s�d�р�s������iVn�9��cg�{A5����B��W��py�MsmF1��s/����3�h :\i�f��`�"C�Y0�fm�~�6�Z�6k�X���H#��e�clee�`��������'�
����ے����J�<�+TY7��Tj�����
��%�@�.�\C�����YfY�W���#@E_M�I_K8Sx�7n�s���>"t1Ϧg�$�Ng��|���?�����o�I�t���|����7�j���R�
]tw"��zPss�K���^�u2�i�}˂ B�D���B:l�
*�q�e"�ӈs�>�l7I��ٌF��է�|��F9�6�MT�Rjmm�kשd@K�&]�np~�}����ܜX�4㯽�* ��dU�C#C7B�~!:=|�p��6���o~C�,I��O`͋û��4ڄ��F"���ի����s���g�-AoB+�퟾����: �����T��
���d7V��pV?��:�L��*f6������"u�������+
�c��jSq��|Q�D���?D�[x���3����nݺ�fzGGG�	�֪��A\���4X&b���f쌓m���餂Si�	c�QyA���U�ѿ1���k��z�f��2Y��9�� �H��Cu� A�1mV�1��������ӛ����������֨�������O�l�L�c�ʓ�N��Yɺ��?��[o��p�0�PZ�� ~F�}��>�d6"������ǈ�'�^���z�֤xL*e<̝�*��ѽ�0���H�0�du2�����_�G��M��S��i��pf9�,SMi`�g�!4���d��ee��3����|������=���B��C������:����V���o��Q��C&�V�����W�XAY���΁|J&Q�_� ��!��
���R?���Ԛ­O7i7э�={�©S�^�a���Owџ_���ܾ#��]��)����q\�6k�r�a�Y��/h���+Ax-�F�$�\���s|L�J��_�����d)��%�Y���%����-R<͡Uu	J���R�@�*jEp�x�^��~ʍ����?QP�#|��N:,�J��`�fa�Y;}��6��6����9�R�1�z֜n�Jr�֝�#��c����^>���s�1��m�^\�֪��s0@�4�=� ���}���B{��-X�Fl8��Q�M����f���KO_��؎�n�������PC���3f?\��F�٧�|��'�	"$i�8�����	�+O���AG����k�\K�2�rk��ݽ�h2M�n�>��=Ǆ���S��b!~lmӧ���\����0� Vh|�>#��P^h�SI/	<�:�F�Q�,^����g���>$H���n�]��L������S���nf��28��<E�T��l? �O�mMR(��#�BKM�q�A�cbD���,OYr�ºe�$��QOe��S�.�%���PWL� $�k٩�������M��W�ѡ����'��V���}Z-��}��K��_�� \	-y�r�@�$}m��l�S��<@�p�݀ra�Xg�ʇQ0N"e^������v�%���8L�!Hi� �M�ۀ��,Qʖu�9���S���e��M�r!ҙ���:��<��|��fr����Q8�����mі_l/��m<<<J����־���L�k�~TY��<�ؑ���"D�B�t�@�(���������(d'PͰ�\��Ɓ�%�f<G��!�y�t�������֠?	[�s��E��"�)��$�g\��s�$�X�� w� VA�pj�a���8��tǦR���Dθ��_I�g�2�\�xU�|�Y�4f}�fԠ�R��
G�ePC10߭�.�dԹb��N$/q,n��6-�,�'4j�-���#�j��2U��e�H#��K��si��*jL!���Vx�iL%�,J�%Q�WS53��4�(�$�����<Źj`��R;��h��+��Ü3*QZ��woj����4(�h����z+��p�`sk���s>[� ��ƃ�H+��l�s3O��>z��ڬ��?�Ͱ֬�����h���%a�M���F$3�,�
⌧�ŋ����=�0��=%׬(,sJ<�3���iŬ�D��˟�D/d�z���p��"uAb5��b��%��S����hX��gڍL�*o�n�޽{�0��O2d�߻�Iئ�����zSrf�4n����j2�tMz'�2 h�ɔK���0Nd�n�����"��+>%q�.j8�ǣXRΦ%�Y���إ����^QRUN������ڇ��n����E߬�!�ȀIe��q<�OPi<��{N��{ą/tP5��DT+����|mm�ޭ[�v�G�;�����+�]��σm���G�����	�9�[�͚��!�fUG��cNU7׻(��ǅ � �(ꅥ�e��F_g�����>��0A�M8M���|Z���RD[�v�����{��ԫ�?�l�J��b�D�q�f.E�b��,eϾ��D�@M%YFapc)�RE�B&S�qʕ�l�f�$�~��� y�Hd/m��W���]��omo����}��-��a�Ly���Õ9�p��(�4.��^��ߚf|cá�6�e�t�|a��b�����(�⤍I+�:)U� R�1���~2�yU����d%�I�Z�W�(j�p�A� IG�'�r�r0O�/c�M�a|H��6�%'F�"���<�b|"��8H��c�8�L����˦�I�d*+j���.U�EfCO�z�%(�r�L�
��B�/��0o³U�@�6��[]<�d(P-�ˡ��z����L��N��޿�p�r/]Ľ�sqQQ��]���L�1�Ƙ�Y�g�֚��얟<A��y`�OGyƐ����������k��q�6��6������6=��rJ����s����px��7Ăpћz�G62��LI8_���R7�Q���@!� ���%�eI�Vy����� �_]�=gﾙ�ed��X�K��:��IΪ�0O6����z�e�>z�='56VV�67	�xR�*��1|{;�������$� SAw���������^����Yh��v�%��`��Ƃ[kݺ���w�����8�nm�g)Q�w=y�R?�S���{��y��u��Y�לO���;�7��K��4�dna<	�ΜZQ��ʫo��ֻV���tjm��a ��_�w`��N��� ����7^x����VfX�1s��ý;���o��3;�'����5�YB'�;2L�q|���˄!\��0 �>�I�Pa�(�qd�N��"wC����1'NݵhT�4K� �k�~��Z�o����� ���05��pº�1�Uz	8U2���q�ڞk�Ví���v��0���ld��+ى(N&�L.X ��iiˮ�ڧ�V?���r3��M�Q��0Z�� ����GQ�����lt2�'����*���ϝ={V�YTm8!�����Q�}�|���`&������D�",�Z�'�r�9���d��Vî��Z�3�8U��N���S�O�:5I����?|�PC[���C�܎��Ķh�&���kN�M�ԑ�c��ȱgt�Hb���o4%Km43,��h��܉�ɓO>y��/����Ր�7�!��o<�������/���O�^^]�	�E\�N���5o��?���c�t�^�O��O�޼�{����>]��w����K�.����]omiyko7�@��HI3�Z ��:`B��	0ҧ�4J�1�*���\YK#�踩��3L2�iG̏S������IEC��U�����6����!�G�ٶbmG��I�5�Z(�e 6�p�D�L�N�8N����`�>Ocös�Kʰ����Ǘ�h7�U��K&S�Y.�4�k cvkRMa*��F4�i�t}�J(7M���E������ O��,]�8�d<�[�2Y�)Z�TZ��wEӫ����cE�0=9�-U��H�)/�:"3r����3~�`��rk��8?�w��lw;�[�Z����Y7LzN٩ǹ��r���K�?T�I3���c*�E��mE�hǹ @���f�YyJ�6k���m��fm־�U	T��`Тǐx��5@V�]�:���E�Y~��$��0"�!.�Ί#VD��jUZK���hD�x19��J��B��H�k iH�I�_cL��ҫ �++A��:�c�=�BR�^�[�ℨq��
a[\�Z �|Ɗ��:��1??OF@u��S��⢙F?�@�u���/?��c ����L	k��d�\�t�R�B��9�q�5*�1��d1�YQ7�ΐ�ɵ���{�W�'!�`�.��t�Q@���%r|�ia&%[F�W�Y%���%!�Bԙ���bە+W۸��&E~dm����;n����7�����,EY���$���Q�!�<Y��Η9*�x���C)���%�3sJBS���Q�����7Ν;7��	k}���~�Ý}��+��@*��\�pN���բ#�ђq��݇HȦ���'��|�'�c�6Lo��]�����Ju�[(�w}Z�����eZf�E?ϟ?Ow������J}ؽ�I���N��h�W�Խ�����\3��������-ϧO�����ϗ/_68�W�%���m�%Ũ ^���⮬EA��$.!���!��a��P�{��i�l���Mjš|��)����/Y-�s5/�  Y�4��`n~�fyw,*�()d!P%Oȷ*���/�D��!(j����d�b�@����"d��¥uR���kժ
2��X^���p�?8G���u5 V)1�/*kLQj'��}S�����[0�Y����hǒÍ�g0DH�c M^pI��9�f�(�ϯ"zҬ�8����.g��ĵ�3L5k��K�֚�Y��V�5a
[�O<������� ��3gΘ�5?^�!��k�0�!&�d2걐�˥N�#S`mm��2���L��n;�7�@1gqYf)�Q!4=OXE�%�E�հb�H��~-�`J�M���Ŏ�z�ו�E�0�tKKK�n��׾��_�����?��;w�,��y-/�~jx�d4A�E��.,�������F�s�`Z\TJX|�LB�l������z���P�@edu�TR�G�4˳\G�� 	c��i��{���[w��z�+ϒ�z���~z�=GÞ��ٳg�6VVVl����&��?н .�ߣ	���מ}��!�a�S�����Q)���v�I�ڎm�q�*߻�p���tgw?�^	��W\=YЎ�B
�c�����;w��BxX�3�s$�QB�$�e����.Q9�9��&�'���_��ã#zy~y�[o��Z�Ng�Ovvv��jB��C�2�Ԇ�!B��r�_t��A�K5[Z�\��H�"�/�G?�����Q�]�ll	t�)�5k��l4��r�'4�y����3�u8tF�>{�t��}p���:���w��w��֛���Q�ymy������~��'���m�e=��#V�q�9��J'M�Cd�5����FQ����
���9a�{����hn�-��!�	E�I��RF��d,�n�(&Vs'�Xj�a j�d���>	c�D���gf�����_7����?>>��,��ח�������z����������)}ʯ�/���������w��ч���\0$,�	n�f������~��/����?|���_�΃�׮]�~���������׃$M���e��esu68h���,� �Q0�'�?6H���8{�0G	�������K��y��+�>a�u�{wv n�s�0$ �H��']6�P�R�g"~���R:<�<��ؿ�h��q�6�&��n��a���7ځ��]�t�g8I��>��^'s�|c��: �%�D��f�T�WF(H���)��/�IQ���L0!�:��yfAD�׏�m���%�R�˘�o&;Nh���'`�x�X��1GQJc,���s���GI�z�i���<FFVҙ�{^���ϝ;���D}�c����ݽ����x�z��Inu:f�5-x��\Y\H�`�E!OzW�y���6k��m��fmָ=}�K�2����ɶ'DA��xX%C�~!�,�0�HB�b�BI!�w¨-����v�M�)��i9�#VM������������f�����ӑ�u�ZF��M^~��\8�%�i(� %����C���_��@F�bK�n?�X�N�����Ө�T�cT-�'Ü�Y
yU�i���Rذ�#�F�.bC��d���G��<L���R,K��6�Mq�:I��}���S�NEJSk�Z���Q�q��w����[�stt���e:�3Kſ���ź�V�eua�\�stm�t%�Tn�r�����/�e�s�1�K��N��4�j���`�ǃ��xt_��� �AW�J���d�� c�O8-yQ��|����7J�Kx3K�IP�<Vd�l��%:塓O��u�J�������-�ź#H�"$��T�t�۵b���j�PA��u�`�=�n���ǂNe\u�p��Z���V�Qy��>�i�~��@�@] ҕ5Y���m�LK��T�b��M�ոs�N�@���kkkd��7�q,���أ\����D:d��RfYc��}kk��ի�[�Yq�Е���Ϟ=KWCi%K���|2첉0��e��t�Q��l�ܦ�\�#/�%бo,�㋏�|J�O��yB'l�����t>����bbCU�v�^^ʱ��j̇C�8�=��%ԇ{��n���[��1V���_Ze�S�U^�k	8�X�R��Q�g`�T�Z�9��Z("��|��$j]�0x�UH-N�)*�Ks>�P�y.�n*�9+�[,��AL.��rf\��J�Ks<�)����)��� �N�	}���F)�QtiJ�i�fm�~�6�Z���J��Uv�X�Uh_E�@����W�������N( ��=�'�^}k�>E ��pW��Pd˫�71�WWW�jd��uVjV ��~�B_�
j� �*���Ht���S%�g���Q��)��EF����_���>����~���{��ntsyyAg	��b���a�
!U��G�����&�8{�au�-�}���]YZ�g��cY����1�26����#t��n%�M1�	���o��j��O>��^�����ߠ�&�՜[Xm����G�ɈL2y�f�����}��b��g_��b0@����{������h(���t{d�;d)�Y8:� �д��Sq�*�	ԥ9a6��H��"Jb2��}�]�k�zL0k�v�"����L�as��)S���f0��,o�s�uz˰$z��an�����P�,G�LD�?/v��?�Jϯ�,�`��T�+ �Εy4�k��kY�?���,�f{޷�4HF�!�4Z����JVd�i\�; ����5ju�^kεe���������淿;�ɐ����Z��z!>-�s%�\-���$m��ky�o��{׮>N[���|�֭��# Le��"(�ln���]V��r���I�h!�Y�W��36 ��KUa{	�C��v*���؊��'`y�^�8v��'?Z�[$�+�>s������wＷpy�:Gǯ�����n�^sP���8CG5�"`�,Ɠ����{www�~���7����K�c_���ww���h`m�:<�T�a���M[#-���n3C�	��\'�R#Ki/�!���u�}q68�ܻu��oY,͟�IFQ��X���R����������ޘ�s0�Jad��An����$)�LM�+�:@n��0V�������p<��t�Cp�s�h�����nwEf��"V���Zi��@�$�9��}�{�E~���9�[��*�P��r���̖)���,O�#�W!�,���bEd ?,��(#u��Q�LU��|ʷ����#��h!�IdHh~�P��6]zܝ,���s�:'���եK��)s������[+k��G�Cǒ����_�5s������Ix8��tG��Y�Y1�|���&T���sRȃ��v�ڬ�"m��f�7�}!,1J���9-n���eUz�� �ecmD�hN<�"_!�W�~��!PD�9�LȾ�J)��0+�)ib�V|��a�ʪ�
��&rJa1��2d�k=��U*�4�9!�@��3��D�/,�g"ыRsL����s�[���f����̵�P�-:�ǜ@%�"�OcWi.�e;UE]���rl]�Ɠ�� �L��iU�����p8�$���]�-/֙d�.��������(kC�O��f���	x�n��;*&B�Zq���`�7^:N���� zn���:fJ~^�WC�O�0�w���H[�	���(��y�b$%�d	U~��q�eL��@��)��,b2��:z*%kz�Wh���H&���
E��ͣKA�ssn}����Is��e��+I8⡧kZ̈� �\�w�9n��3g�`�ǈ�3@���\�7J&�w'L��2�2T�9��8WfzV�$Rq�ذ�,'�ph��_���=|��������Ɵ��8� S��`B�����K��J�$e�+'˦	9^�ј!����E�@рl�.Bkђ�`"�Y��dW��J*W�)�;��ǅ�<�DTQc1�(XM���H։�
��2�����x�sD>�n�WVV���Noh����;}��q���@��ö)K�����g��4�@�2�O���+g�,[� z��X)ź'�L,,��"�Rg'W`N�9DQ�\n�Qe��j��j�ʥ'4��,���6aO.*�XuڬHoy�^ .�E��g��>ܣ)�����u��BRq�d�|rr��Jٝp2Mr���J�k��fm�~�6�Z�6k_��LT��R��W�ڮ��/z\���wZ��'�f4�Ê�;����2Yk�EFXN&���$�Pz�CO1�V"j�!�4�#W��b+<��8U��� ~�o$���(�R�py ��L�j�B;�M�"zQ#��t�#4p���`2v���N�����&�3��NOz3��Z:M߃��k׮e����Z^GU2b�Qf����>�Ǿ��d�a�1����'�I :xd�Fi6	'�_z�:b�B$0����!1v������1�Ԭ8��"��ј�I��9�so�o�5�]8��o~�3�}p�������gB�ô&� a�(�GQ8$c7WH_!#;K}HbEl�i�i�� �"2�	݅��xD`���i4	!a���g;��Kc�@��a����t�q�ˣ(I�è��xا;�e�q��Pd�$J�T�-eDEHZ9h"����!7fW`�
Dʹ��Y���r�'��� ����'k.ک�Q�*�@�g�<P��r\2��6�q����N-�y���n޻~�:��{�G�s���=8HCp9�T#�,P�#�[�5��[{��f�n���^�(}88��:LT�z�C=��2���rV�0�h���P���BK�SH*��C�(�Xx����B<����&��i:l��u�[P�k7[�55�:���m��p7E�'p/�~B�ሠ,����O8-�B��V��>c����,��4y�g�������B�6Ϟ={|�;��P���s�'�|��O/w���nG	jB���d�'l=�OV��'���E��-��[��`D�5W�s3�����(��z��n4�*c��u4��&ߨ�JvR��<�X��B��(_�9v�ռ���/���(x�y�E�t�	��1-�w����ڴc"~56��9�Kʛ���!0�c�k���g��:%e�Qz`�wT\f�'��ӊ���W3^�l��+�K�4l�����	��f��@"V(0�,B����l,���!��(�\"=%|f�h�+�'2��d�j6�]S���]u�t��ң�Ngld�p�����^�'�v>��?��R�[?{���.;ͻ�Hw�$l��&-YM��(8g�yO�D�ɨ��Ff�0L�ڬ��/�fXk�f�۴(��*�d}ꩧ^y����"#��K�m�9�WWW�'���	\]��8��gv��{��!Y�B#S��bH2�H)de��H�����/I�!t�qi�ʒ�*���A�L�0k�` �x��O�������}z����P�������"M�Ԁfǹ�<��ַ��8}���������vv��x�GD6��>d�����p�2��ziR��R��j���Z�K|4A�!�A"r(d#�1����|�^|����pq�N���k��{��?�'�+$��.B���Z"��_��j��Vl�F�pdW�A���J�BR��'��j�%\^4�`c�MK>��jL�hZ�,�@��dve*�.�՘Y���S��j��"[�����5��?��S���81��ޥN�d��bzv;;�Hr�D/���剌�)M�����9}�qgg���Ы��?'�~oY�x7��E������r��}�k+��>���o����.��ݸq�����N�3��
e���]��[�.�-�0��] Wj��C>K�R���{�Yf�F�L�+�/@%�EϰF���B����GK�;�����������~
:�B%1��l4�������*5Q�f%F�'��ν{�>��I���N�A��Gw��7��9��Bj�4�2��)����G*�r��p\��m���Y��h������0G_�4�ܳ�]� �p@Gz$_�:�o`��=��ț��-�Np�4}Ȣ�,B���%���1��?�8�ĲH�OJ���Nt*���Qy��;#5��dW��T���zSN+޲H�b�A�˩UX�d�
���`9C*37V�xV�~F)بK]�{1ἒ�I)p/ə�_��S�8:밻�=4�~�.�#��gq$�S?�1_�{<����ht<����Z��w���۷�����WF~��|R6���U�<ǁ�B��|$�*U���`痑��6k��em��fm־�U]UT=�V���8uMz:"�jE��Ag~~�ެA�yu�l���c�@�z�})�܈c�h�¿Lf"׆2�ς�,	$4l�g���\s��m��1����Oe'ZyY��l�:�%�����3M8,�l�q�Ҩ-.�߻u�^�W�����7?��8��'1�km�cT�J,����q|p�V-f�foo�m����7�N�2�����'o��=�e]r��˕��&��`^>yӢ[6�t��0-��P��GP�Kh84��slP$��MY��v��n��@s�$j6��g�.\���R)PA���,�kuUS�._!���ߣ9�?:D�b����-�p ϳ�L%�M&gދ��I2�h��8� �8?7׊G#��Ȏ���-)0H�0O��X�q�<K�S1hPR�F�똩D��/#�e[F\���4z+�LRؠ�pbڦ�����b�ҒƼvݷiP=�ql�9�D]b�H�+t+R��"�ߎ	���c�H45SHH_�5��,+��=ߴ� ��#��M�{�o�s� dF�R�PGV9�1�y������3�ˉ�����0�y���-3�����$����fH��(�0!krۈ=3]��,OU6%�\iή�͘�� c��i��	r.�[N�`��_ڵ�\��5ڡ;l�Y�I<�Ӹ����$��H�H�����7����B��'���(���m9�n�6��P��M����M���z�h���$4�C�lG��/�\.���W
����D�`4J�߭f�T��%����vn#_�OƽA�s5I��@��a��/2�yN���4��2V��=��0�Wj��Q'��zp�O�6CDd8��	�<"�	�̣;�#��9�Y��e[�J�쐙?��hc��R��&�MhH0G�d�m��\�X�w�ȡr\�l0�f8���g�H����VˀBpg�L4c���Yj1�z�uJ� -O(�S��u�q_�ep�5�\G�1z�o��C�a�[�'�0��M����G��L(65��(��	�&k&�셩
G:�}��Y��7(4K玡E�fJ+aG�6�L���0uY��^3�k�f�K�k�ڬ}q+Lɓ�=G�'D���0�W�$u��ܾE�tz������ea�Ӧ��l��&�\dDfSB�b$e��\D�s��������u.	6��g&��Ν&I����K��W_}ur|LVE�u�J�=Ĩ �f��^�p�ܱ�^{��ew��|��d�̖��ݏ�r4`�zswww��i���*d�A;�5�.��A&��E��aqJ�F��AI���Dp�3uC����c�)�Y��a�����N���{��b�����t���������{��w�z$��,���-���qĩi8�|��}�0�x�$Fm�������w<`E�:�������R�azN���U<�V'�Or�b�L�-�3��d����t���5Ķ�L°ץߩ{4J\4��f��d]�(�H�%Fۂ�X��0�E��t��NZs5|�NO^qml��xH��9�O��d+x�����ۄ��ߎM���p�z ᘫ0-, <��,�&��L�LN��7���Y*�"g)��C>b�Eɰ̓�wlQݠѠ�J]���r֟r̰�cbNg7Mk��kF��˚�`6�OA0�U�*��8W��N���zo��[GR\�A���uDI_d��h�~3�-ʊl6��h�:g���6��	�Tz���I0�!�ָ�,�����/�2Gj*mI���?��a����hss�o��o��B�p �ϐ9��%���q�R��� �q��� �K+����pj�90��imz�k��՚�(��'K�v�S%�7T��& ���EI�\\\ª�Ɋ��&�S�H�Փb��!���(B��?Q�����Q�
��VA�T ș��Dt�-s��Z��� ,i��������#�o�����/��&�b8��¡8�dU���T����s�R�}�e�ڬ�s�k�ڬ}A��!����{�vv� ��%��+<�_ �����bY�,�3�-��X���y���*M��t�HE]�ȃ���r.&�-ǩ�\syu���ӯ��|2�8v?KLC�B�.�[�9�`4��W��Y�����z�a�<3-RԏԀY9�� ���ѱ�ϟ?���WOQ{������������{��ȣ(h�i٦A։F�{��x÷������6���!+� `}�6�$#�7� �V��5�'���\ȇh����
5CJ��h<N{G�;��X�����'�j�!Q4�UQ��պ�j@ Iqzc�,`�-��g��&ҵ4����L4����\�Մ���n���N�p�Y�|���T��l��B�B��'�]�*D�}?�;�E�󬰧l�Fb�ң�����X2)��q FW��6|�-�8Q�7�Ө����4Z��f��ni�pujS����"�����h�ڈ�c�Ǣ1�U�D�ȳ-˘mP&yu��Gm�r����������A�n�i�o?|�r�IB�x8���t��2|�"�'�$c=z�tMR��Z�Rk��I�rL�7f�]��	F�D�ի�n&D��HBX�,�h��ܰW7֛i2NcB�#���hzM�ԇ��%������;0Y���8����� �{���t;�I����r�`g���o�P��Fa
Q��#Z�0�	�!�@&3h�G�Q�q�n՛�[0�3�$A��H:�u����?���2��85h��u�flB���Ylr�-���jE	��Ƌ
1����q�vñ�ц�_@%��� ���Vy�VV�2�v�]��n�(�0�������tz<~���+W<�����t�A���$b�v�X&��:3m۬0����Ձŗ84��W9!|�D��4�C�|�#,A��J��j\z1�vŒ�tuڌ7)s�Gz�[���ʲ<��k~����U
�Fl����ze�m�o�G�qs~Q��&�q�KZ���?�9�Gv���<�J�Ѝ�-m3�=�P��2��v�%�Q�����j�ڬ��m��fm־��27��h����@� � !��$�����³E� 1B:5\��1)}Ut��������B�t���VaE�Lc�
��z��u��#A��������W���믿��+�'6ZOj�p�-�2dн�.��{�[�p~ii�A�0��O<A�����v��{����ٟ�1�*�cɭ%��e�<Ѹ���
�U�B1�
l�f�_\��6YK��G1�Յf�!�G�-��ܹ�/�H������MֽT�B^ك�;w�����Wz'���7G�Qse��9�soooĒ�"��s,�C90�<Ϣ��Cɲ�8�IT-��G �Y�Z6��\���X�lɣ�RSP�(�K	�*�ݵ�|�!qUey�w������n������b�В,¢d�Tt���%kni��J|�HHX��3r��R�ey�F�ow���9� 1�5d�<�{I��(++%��M��Y�U�M$+I�jX�ɏ�M�.�Ӕ�J�9ɮ�W��ICB�2N�s��!^c�Fq�����!i'�����3�H?M��Q����~�1}����]�vog��W_�S��~n���/X�Ԃ0�rk��fI;O�v��U���~��)��������fj���B��Cʝ�~�Ԣ�̊5�x�jт�6�rg���j�O=�����v��a��}�՟��r��h5љ�Ԫщ���7����K�TRh-p�n�Y�J`4x!o�x75�Eq90NI$k�a�o�F���R6Y���Y�,$A?�~MtS�ݤ�T+i���;����*�4�B�KQ��٧8�d*3��%�\�qU��3G��|c/�a�w?��՘S\ސ�#��tP?|��5��W
Kbk�!�:��#��/��F�ڬ��/�fXk�~��4.�~�L�)��a�5��Y8���x�&��o@’�W���"x� On��%�YU\�*t�,M+����U����B�|������)�j5O���× 42�"�M!&5�4I�5����Lxr8|��g�^�·��>��!�B[��uA�R�r]o�����aw��#;3�> ;�Ɂ������ۃA��h��-,�h�{qg,P>��Ђ��]6
jOK!����	�3H�Z�I�aaa��L���U;t�$�B([�5��n��M�����է�!+���3t� ˸�2b�����>�h��,��=�L���[X_$3�e��z����t,��\�Ϙ/֥�cC�5�X�^��Fd���M�\�&��u6L���1<"���E�m^�Rs���.<ϼ8��ёp�Vn��M\(H���L/���W(5�'�����fs{o;7�ޠ��װ-�+��`�iĔּ�h�y2��z�"J��	�پce���./T'C�X����J���Ad�~��f�â^{&�d���ALv��;��&��ƩJ�^n���l,���\�o�t���&��$#�!����4�l.����dp�%��ɖ(돠�fP���7`�<�Ӝ�4匟sm�Rو"�����?�����L�����w����Қ�֬$��̊r:cB�z���-����R�*?]�<fiDӠ�2Q���4���>��s�~���48�����~nBX?� �s�a��υ�r�-�\���ݶ-X���S��w_�&��݇4�g���Xh��=�Xpo��?'C�}�=G��xk'UF����GN�|�d�Z�٧�ר55M���Fs��g��a�Qa���P�2��V{r��m6��c��yĦo�4J4�e[������	o�l<�����u�Ąoh^�Oc�!��ͩ�����L��A�{8�S*Yi����pDEv���{��J��AP��jZ*c�傘�-����.����!�K2C*��ޚe�Pj^c��C��B������4Jk�y.+����|D�w�ʓ���o�Y�����h�:�]I�4@of��9'���ʱ��|���(�����ڬ�#m��fm־��|*-&3�b";��a�	�����gE�����JnH}!����Z� O�4��'��^O5	��x���*��y���ת�W�Z�V3���K��Խ����nñ�{,�t�6m���(rPe��w�yG5���8�F����>Y`ɘk�$в��΂Q��+Y��I'�b�u��ē�ye	2����e����Ng�D�P���l2Y�������/Un���v{<F�Q8	Ț��$�|�ep�)!2�H~�����3s��:p��Pp�Ղ�'l�=�~���$Y0F���Y7�T+(���8�j�"�6�L'���(ӼXiBR��T�=��ODM�����q�P {T��.I`�f4,X�A��T�-L	$R��S��+�#���\����۷o��.2��B�L5�R�x�G̰$�0��)s2_:C+MY	<q>�§�gi��=�L)쒙Q<�<wE��IޑY�¥�M�0�c�����i�ߺu��E�O���!{�l�8��z��m�29�]�9s�J}�F��sqĀl1� B�t�_&ɍ7����u�R�g�&	`�n��S�h.�eA�$����E����N���?��7]�V��S�Qa|4��z�O�(��$�Z�'��t��P�u  A_�����?���{룏hS�Zt&��|��'t}ڳaӗj~���pUwi�;w�ʕ+F���jd� ��P�Iǔ[ G"m��0g�)G}gv�B�r@��L<,ۮ�#�d%��yy+D*�U���&�\
ٿ#/�&U�!}�3=�ώ�:�9؀���Cs�1!� q�
�&g�wf1�3�N�o����}����%�q��Y�d93��(�C�w�T�Ŵ{����5k��˷֚�Y��6m��*�/��m�,�yYx�GfZ���n��gE]�@��VE(�t�ִݬ˦�;�V����)J�S���u��������}D,3Oam�}�Lz+��+�=��o�����;4�v�VV�x¾m��r)Չ�I�dqq1q\3GIz�̹ǟ�q�̙��<Y ����ϴ�vvv>�����q�.'Z���5|/�3D���넮�*�:�~0Ա��x�L���8,��Z_�X^^��s!*����t�	5�|��� �e���{�g��<Bz��{��w�B��!�̑Fsz���s�֕K�h4j��;�1���n��~��:E �d�-CU,ef1 -��s���y �q�w,^�*?�f�@�r9oG>i�O��*"܄R�F9��/�c��"ؙfQ��3Z�:Ecif�"� �d^�e���%�٧i���GI\��� ���Udv��#�[2�:�^��X���ӱz�%��z뙆�9k�� K����ٳg��/~��;w���ןz�g�ã�Ǉ㌾4�4�sX���l2χ��l��h�6d&;>���T��ɾ���'Fi5����R��>�JP<Ό�l�g8���1�Q"3~2����g�3;Ђs��Rv���/~�+�j�"�{t���777�n�%�s�n?[��Q��\�Ys`c _�U�O&藣˸��w}�C�;�ծ�^x��瞸6�w&���Z�w������_��_��X� ?d1�[+;�F����&c-Cg)ݔ��b�w�������cB/����A�J����x�2�3J5��B�S�Y���XL%.�j �IK�`w�4˫�$\l��-��չEknyk�x�C��9�o�Yn����1-�2盍ǯ<F���\� ��?�|ڑ\������U�Q
�ȁ�	~�D�����4��qЗ`E��(p��9�^��E
�D�M#�D�i�^��p��2��&�ȥ&�b�ʟ5	RZKQ�54*�	�y�a�Ԩ�H�lk!zR0 @�g�BK�%��j?��Cȯ{��X	e�h?B<�j@��#�i �nV����}�2QO�ڬ��?�Ͱ֬��4����4Yq��"슝��F$�J�Vz3�.�bYY����kN{�+�$�Ӓ��ο���x��i����/�ZEiN�m�~�d\�~�:��+����*��7�M��΃��	F�8��A�=�CA��ƍ����z��������O?M�?��?H�a2��Q�t�a�r�dU�9�v���FK�;t��i25X���t:�d�8v���*5���aa_}�U�)���aE�먞Ŕ��2p�x�B��+B�3!�~_ZZ�ta�:�2J�q����M���'�\�X"�*��I�YYU)�(#�FE�H�Q�(�e
�{�K��z�^)*\+��3������"r�-��O�r�ք(�7뒗+Ĭ�<�
{��&;�um����]&��#�V+P�O<qaqycc�~�`�Y��x�����/Cs��z	u!W3kS�,�4�XV.�\���8!�O���0�9E��ɮ)S%Jʘ

�uބ�WÄ�Y\���I�M#p��%��pإ�J��`n}���J9��r�ʥʙ{]I�4���r�L�*EA����H�b�?�<}}{]��ơu�\�Uӥٟpe9ȵ����KB�B��9����i�?��cZ�����1Z��� U���!e��/k2����N����h����;��,//?��s��(z�����[��.�A�=5i|��_��}�z��{�A��uL�J�E�$,b�F�je��=�ܕ���V	T
ʒ�8�p�a��PLȊc��]&^���.+%ʴ�q����'�A�˄p�gS���+�o�pC��Mz�^0	Z��ˏ�2��ܺuk�߃M��lCV�pV&�`�٧Ak4���B�^|+p)��-ϓU�C�����5k����֚���V������+V!3��HH���Ϧ0�g��4=7�w���!^��90:O%�,Qfn�6��Fi��2��ړ3���N�i�pYՋ�u�^4��qh~���%og�����H�Г(x��gO�:����v�G��,63�a����
*d�l��2	�Qͬ�ܜj��k�}���w�����i6̕�����<{��P�}#6�^�`qi��w�!]�n�d��Q�$�$k,�@�ĩ5T_��$v\��$���GF�6N�����Ked��]_I�0#���0�qa�T�$�s�λ�����o=s֔7Y@��&.P-5�,;�R�����-��f�g�N�違��
Ñm��&+��ִ����b�M�e4F�1�A`Ϣ�,m�0�`䑅���N����"�lR�0lc����!vU��$��[�b�n3d���IӪ��bt�6A��oO���PH�\���1D&0k4�y�#.�Q {��^O"�,�fEf��"6����TԦ���`L��(Yq��`h�������A�&g�_�w�\�G��z�ݶ�ƓO���߿��.x\|H�Tm���FQ�r��s6��J�[���Il0S0ySe�ma��̥L���&��r�h7-X�T^��M�`u�C�T~KSZbd�b=/��t�`� 1BMN�s��[g�.�>��u���	��5W��UFY�mAW�1�4�u��b(0"elah�x+3��iIx�sZ{@������l����De�+���C��kô��M�Qå��,��3�(���0�I��Z5��lt��?>����h<{�i�Ԅ��F�$D�fZ��g����
Dٚ�Ia0�ɔ��Us�킜���3�A8��:<�������� ����M&�6���QfX����{<�/,,$.��lca�vܿ�?�o�ű�S���D��r�	���əE�9H��AZ6�JЂC��$EP�	�#����4"[R�'(5�E���*O�r�[�a���71�)�s]���|�P�s�\�8Kc��yB�>���� �ύ�R��87��R�����[�n�RI�Xf��U���8ɜı���\���9��gp�1�v�����-���J���[[�[>L|�-�)��.���nhH�W�౔�ek�ڬ�cm��fm־��i�pH���T��Sk��"��<M�|*C�W�*$�T�?7���p�Z(�Z�j����v{���^�7�v�I5-]�,I�K�y��S�K-�m|����|�;/��q���6�Ж��sU��`�r̔�v�����4�Q�]��R̗oa����(�d�w�hk~~~=��]�;��(�I�5$?^���Ru\񢣲6��E-Y�A���8�.����GC[l���[�wϞ=;��
T����7k������g�S�C�(�0	� IIF[#�i��A�c�^쇎��?��?�Gt��h���Z-Jju�l�I
ICU�ʬ���xƽ����9y��@�H)��YLd��{:k�o���V��G��
(t8�Is~�э��di.����Yc��b�`�1+�I�*b�7<
%�O��$f"Yu°2�`���r8U�A_Y��6u8\���/�y�s��L5H�\�u�2����ܮ^�@c��o���*=�C��Y��
h#)X_I>���Ռ#gU$-�L{��[5,��fL5 ݱ |_ֶ���9�s�D��%�_vyh�h���,���X(͚<��k�,c�����޽{p������k<�ɍ�(��]�vM��� @5%vU#��}� ���DaƂ��j�����/���{��֭�� �+<E�5D;�o_�`�<|�a��B+
{�:+��PՌ���S~MP���Q�qr�v�mh�����ls�뤨�"��O��	�9�M!R�\���t���>|�L��A�F�~�eɻ��%�'�AOb[�<?l�j�;��z<��ú��&^6?	3g��l�>����6(c؎�����)��hQx\�<=/݊�H��?�
;;;�{�;�X����IM+e5���R�y5��ַ,��H܈P�q�{oy٢>�G�����R��h��I���Z�E���5�E��"�{���:�f&@��@���p]5��Ⱥ5����ӟ�k+TYۍcXZ��t���s����7zZ�{�D#{Ǖ��9�mfW��Y� Xr~0β����~�;�O���>���#J�)}�{?x�׾KVW:�����\�A�l�&�Ζd`�ݸ>蛲 ����4�� ˊ�o��]����מz�z�3�=�t�By�Ng�l�=��j����?K}�/' �S��:qjs��tN?'*3�w���d����U���D�kt�x�r�������"kJ�dv��ׯ�=��ʫQ>����Tv��jyy�zx6�G�%�	_�g�O��eb$��ᘒu��(v��灶ʲ�_�_�B(��d�&,��T �p��ħ�#���͂�eY�q=�U8ik������^U���X��ƌ�*�b20�4"dD�*r�f�Y�w
�܋�q6y��-p6t�����/~��͛~V---��%�9VH�L�Ph-ǣU1�c"#V�F�c�~p��GTF��k��)��!�B�A�J���3��4��EPsv�O�R�B�ޯ��i�����撝e��i|O�'�_���&qDS�޽{��qfȏ�_�˿�{qӔ����կY>=�\z?�:Q�����(�Le�	;�����7� ����xE|���.����{{{d�Sg��%�b.�5�k��(�����i��!lfsGQ��镪��BW���٩��)�,���z�jk�PI���|-s�}h�9L�:���f��g�x�[snv�L��F�ғܚ�n��''Z�W�v?�%G����#i�;�,Y?��Oi�q�p��=ک677�7�{_�� ��Z?������:�h֔`�>0���M�.G�pHTh:]�S��N>�	W�&v#�O�^]������s����tG��EY+q3u���q̛0yD��{���3ׯ_?�&bH�cn�r�M{-Y���h�D@ӟn"�BO{����x(Y95^����~8,O���tXt�_��_�\�9��xZi_�/(�4�ju(H-ڢ-�ǵ���h����&��UFJ�`�p�n8�8�/���os��G,k�I�S���5�Ԓ��U�����H�J[L��ͦd�)��:95�~��2��z�kѻ����'?��#rv�8��$�q^��78Ksee��x<����j��q��x�[[[�B �_2��*%�Q���%��4\�PW�aL�{�a-�4��W�4���4G���u�RQR���n/�0�C����,W	iӭ�OǨ��/1��y��Ӳ��F�*�Z�F��mb��qͥC�'�C����F2���1Gb�o5ǔ���|�A���rY<C�u��t���e�.J��~��~�݅��ז�"c49>E�~|"��@����@!;��[�ʽl:����n�l��v՜���C�d�6���1�j_W���666p��M4]ܮ]�H�{�7��.\���3���t1����=:[�Ϡ���,�G�B�a��
y1��+�$8�Pb�p
u�|���vY}�<A�*���r�s�\Y�&�j��9��E\d�\��6�j�3"��T��X)�&�Å�GT�>���B}j^,W��l�Ws�v��t��4��(�%R�]��0�,���Kg)t#����,@��� r�.�w)���	��Hkܩ^k6�+~Bq�{��Sf�%�Z�P�O�y����u�k*�d��MȌ��;�]o2y��X�+j��HDQV��:j�"���!��y�Lz2�u�}ހ��PX;|�6�:�"꺈:%I���Oo>�ye0�ȁ�\xV��h��-|�E[��mZͥK��eX�5
�_VK��2uX��n!�U����za��i	;��[��Iƈ�B2�FczG�f`�p���kd�����j6�=��bܥ��o�I/�n�C���.�����b���'�'�)b��),aq �dЉ�q��(��!b�F�9�q���nB\:�P�F�3���q6N��j��wC��1[����Vn�ѿ�h�L���a��_
/��X��N�^W���+J6Xa.U�� �w,�TT��5��&��&b��svW9	}�AVF6}�:'�&ʅJ䡅�<UU�m����f�]��#ko�3��%��j_[�sV/L0 ;(�
2��jCF�q9���,O� T�v\Gk�A��I,*��M�ٍ�4�/UC/Gv��� �*�AQ�ȝ#���#+����D�s��ں~��E������G'^7�=>(�tfK�*�*V̀;��f��� �́Q -��XN�KYs���ђƨKI��h�Q?1��ZX�g �^�`w9x��:W�Ґ�������<ɒ$��Bcr�VW�W��ntzxҋ�'o<Fl��A.�s��ۓɌ~�iJs�A܉�C�d�Sh��kZ��ʇ%I}��'�='��T�T�����FaAn<�G�^`�3[ ۍ���rS��K������*_;aԈ�Y���8�>��f)�RiC�� JZ���k�k/��Inp�=�s(�|ui)p�=Ȼ
�Ad+HS_��Þ	�G�Xr�G��,Ŋf+]��$��{x�uW�V����;��6#�
��5����u]�H��GH�3^\�e2�������o�T?����q#���b�G�
մ�zJ�5 t�w�[U���.w��V�,xh<�	�Oߤ4ݧS�F�(�g�!o<��B*�&��H3I�e/˧-1D����pۄ(��x�6��:�.�����7r�j�AW}8˜N� ��]e��ŋ��<����hk�4y'l����@[0g,ڢ�ȶ�m�~L��sJJLef�ᇌ�ٞ�+~�V��rs�d��}*���&�wŏvd[��V�}�����Z^Y7\J�+��$�Dd?��lv||LEt�������J�7�w��l`la��qRq�&_���¤3f�l�^�Pg������q��0�p5�@���7A�����F��?�rI< �(ᵫ�����r��֚��4tZ�f�&Z��b,�~9�/\�`����qTC�b�(��U��nd6�W+��\*���~�G�:�A�9�HA���YF �%�_���a�|Eg����h]��Bև�28���׮]������۸�y�ҥW_}�.����?|��'?�ff8f�ݭ�-�Aw:D,?͙��=f��:�%��b�*6��};�
��Z��W<dF�z��RQo���:�O1.A���O?��|t�ʕǮ^�y���_��ۣk��=�r���!]9����׿��o�ʙ�r��X��K5���"Q���hDw7��{��QP#���t<o�>���uMa�����|&-�<.�yQ3�]��·��y�%F?��=�}�51z{^�T
�9ż����Nl�����ż�}f���8`?ϧ�^|뭷&��/� �!܌���28�jg,5�p�L�Aw��uAjA�
��Y��k�ɜ#G,�ײt����FM��ôK�&�Pg][[���rYqo��Gj-�ed h
��`zt���+e#��Y&��p�*.���L�l�!"g��NX�dDh�ќ�@��{������_~��kO?��et�/�V1v��Zm��Ƕ���h��c�<��q]��YP����r?w�t8���A�YZT��s��'s�L#��R�{YM5E]p����>�B��B�`,�n6!a���7R�m�K�O��Y|,�å�Оkjf<�T���)�o�%�^JH	����Y��*'s��t�]�/�����d�n�"�L�kcٻK:!�7k�^'���XLF����P���]�<��u�����������NpE1S��eE�
�ah:a�Q1�t�:��:��.���2�s��UmИZ}V��n`}$M�8� e�AY�6�����؍���
�n�7j��O�>t �Y��r�����Do�䨾���ԥ~���"S�cBM��K�/^ȎFGG)G��s��W%���y��Ǽ�Bo �F�u�I�C���lP��z�?��q�a'NP���fe{m���ƥd/O�� ���N����A��H����;����+A�a��\��5�$��3���7 qd-���dxEsf]�� �iQ�^7���'4������'{|�����y��ֽ�ڷ�~+���� cu����^|᭷��&��nV�p����:̾0�f[����f����f�<�DW�|s��*@ƜIl��_��tV�TErEdȅfU��%Ϋ�/�tV��Yp���3G9Mlf� ��xP`7�G'6s�{��)n�'�o�
ޢ7�N���1��M5��������"�2���e�8�h�v�w���ۧ�n�����'Љ�̦�t�n�<��ҌR�	}��Y�YU(C��4΄���Փ� pֱ������$�Wy���]�69�>�<Z4��N�:aJ�$�jS��J��m��֎=?��(3:�`�FwqttF������8쌅����O"6�O"�5ӢGu)�5`q�=,�������h/cu�ީ�L� ��K�Ԁg���[셕O���P�et�E�uu���F���-�?��m�>���<�y=��@H������t��8 �է��	n H�X]�.���4Ao����D���,����y.��لu[`S�2���9�O��u
�1#�ӏ���WY����!�4e~d_
9�e��˽%D�aF�Yՠ^?�#�� ��R�?���{>g��ǔ�%��͛d�Щ���  M*E��jQ��~0,\cbĞ�ܹ���%�1/O�{�Zj>\�N��,2DKb������; ]̟F���[YY��?��p���}NKs�����8�na���[�-r�P$F'5�}d�J�hW���ÚM���e�����W_}�[߽w�ޅ뱒�sp�P�K��r� ��D��@q<�X쵪��̸�,��ȫ�S_�ti��@�ީ��]�7�S��666~����G�'t�"���t�?����o����P� '${Z��U��+̈́"�͡.������4�ə�]��Woܸ�[^�x��l���Y[_�_����=���ի'''o���� q��+i���Wi�u��������t:�^�r��huu���>�Y��/|�R�կ~uz�N�>}x�����
ʹ���_�O�g��T�eԜ,�k�dB���a�G�^p�
�̖���p\�)EZ���'����� ?��R�6���"��n��p���7��b!5W�%7�^������k_�#��G��n�&��'��7��f��*�����Ĵ�m���V����r�G?w��S��h���]�;��J)
�����Ց]K0%��.�T^�Q���Vҁ��ԍ�2׎2�+w�D!����!J+�(�NW�񶶶d�n�n�C3m0��'Y;ĮrZ_V���pV-�X�ڑD@��O�h��`i�җ���_���6����f�%e���<͏TT[�E[�����Z�E����Z-at��ef�,�0����~�w�Sw� @"\��r�G�'�^y����V�x���5��X�Fb̥��F]gߋ˒̷�,Q��l�,>Ʈ8��ru[|G��S9��2���H���*1sd�8.���L���F^TYN��M^:�9��ex�vyU�.o��-Y��Q ҋ�D��0�*���� �O��l�Et}��HY�gf�ѭ;ЫQ�[�(���(Z`*Uy}���]�t�s���W�����Q�G�
&StG���F�l��0͊��iVT��̽�Ƞ�3M=���d2.���)�{t�:�������t����t]���p�U\�a��F���䱲,���С��td����ٗ^�6ɞ;�4*t%k���Zo}����w�-�!9�@]�g�°4�(�Єԕ���C�˫\�*�3[��@hh`��ac�<�8Rr#��3��yJ��KsP�AQ�x�����{;��]��t������{�~b;a���)�W_щљ@c�a�"癍ƒV��Y���5b6��"9턵�6�W�_�t���p<�.���5������//�M��d�V�~؁s�2L�f�[^��+{J�a/��p�I��>�We���["��Ц�|v�[Y^�Շ�}[{毶�ȹe�͒��nK5^'��<��*�ʓ dC�g��}���ǔ�Q�����`�S��)NZ{�3�I�cb=@���(1n}�s���E�!�Ig��p����1��ԕ��Ck+�o���ɣ�\_�g���ձ�pr`�n��	�P��X9��͂�+�
W�U�0�EJ�Bt�=^��Y�P��d���G��Ǐ\U��ů A���ȼr����xg1����M�b�[���t��� ~������p��h�4M�$���i_�tiy����!��YQ���#�&*��O{W��"���c_�U>�z��M��&nYD�Kg�����ݑ���W>�z���5�	ݯ�1Kl�f[%����v&��h��h��֢-�'kb7p0�+|E�Յh���(��N���o2hz��I�1���6��@T��zSR�P1 �ؒ��	X9�Hb7DK��p=�
n.2��t�<���qR�ۚ�fl(��~֖`8�
�>y�]����NB�j0�cz�ʫ�`�[T@]�1�¤cR���%⣑��MP�����..3D+O�����ׂ��Z���T�s||<����˽�sc�C�[�{U|AT5:�Q� y�>�;��)҃���ZJ���ݣk���x<��>f��Y���N!�6u?��v�+++���g>����۴G�N�����{���z��T��d&���]^W��Lv�dne!H����ɤ�80?�&�	�Yl��-��g?�ٕ�M��|@g�2�GK�֭[KK �����m���;w6n<K��ɹjI�.䣯8&����D��^K�q�,�z�����F׀�G@�.]�J�������o?����K Og��N����.�h�!)�t�J���Q'�x���+�~g49!�{zt��w�]���ח����/3-ex��퓓�k	4�d���>�Q?�fYD�����XY��{G��S�p�v~>������~v����J1�X�/����sS�4��1���T}��ƶ厂��2�H[s�^�x���<�-��n
���������i�|��/^\c��N�w�޽�L�t�;-�	Ӯb%f���^�M��y�N����N�+|HƴU�m��3"e���"Z�AVзF�����mл����~�_����z�z�I'���6�����u�H\�E�dm�k-ڢ}�V���!UAV��5K�q!tbG�zIM�����ԏs����ɬ���^b�y^b�,��sV	�
2�}����,Þ-<�j1\#G�KB|�����R6E��c��d��N�^0bܾ�(6�������M�'�R �w�
�jQ6=a&��
��&:<<�M��Ѥ� "�,���м�1T%P1mџI��r��J��{6N�hE�Yf� &�OM���*��\c�F��zƳ���z6��78I�#�h����j8L�H3���N'Y��EK�]�(�=[�fy9��m���K���L<x�X��#�ϸ�����CZipc�Jƴb0���U~��	�"M��o�����f�30z#�CV�R��YGY��2��� "$pӡ+�P!!���-��_
�A5'=*L��|F�ݍ�% �yl3��
&ɠ{�#d��t=���N4�y���ׯ����0=��S�$�Sh;�B�~25LKgkRn�+VZI5'�
O�>ԔP7�"�Q9ٯ�cU���E:;ػ��,���u�q��F�'�lJ7eA���.���r�i�jj�4/��IJ�+`��AQ�i�w��fE>�fdگ��YS�(X��غri#9V�!�/���Z����3��|*�i����G����p&�}���B�:�aԁ�@O�d�h�v��lV����S}�T������=F�LZ>� Ys��mp�:��S|TW_K̈́�yʳ@�ʊU���#mn|5K�B&rʈ��R�J	6�tQL�) s*(Tm�T��'Z3�L���TUY�(�%4���VE�-�*��i_�$Z��4��

�F��`���v������%X�^�����0�Ӄ�|r�!�ӱ�^�aC,,�2ڋ�(���\v�(�[tG�.]�����N�.��q�<�V�yt��=yF�"�J�SF�I�zpd���6?������WTy!�
�i��3���o�բ-ڧk_k��4}�A�S�FO�^/.3�2SMQ�R��j�z��-?��'6M�E���:��϶P���t1S�.�B�֕I�l���C��n�2gk�J\�V�L84s<���x�N����4�>��)�C���X���(��:�9�����]�W�����f ����NS�ً�R�ɚ0��Q�Ug�:�|w�r��*=d7��j楘� �#�E~pp0����s�H��20�<1��t�!�kMN��"��Wa�^�p�����?��R:؝�7���&���uQ���{Ã������c�E_z
��cW��:��'5$E��H|�CբXRIh�^�3�@H0��a�qA�x8������?����,j��}?������>G7��%�����铗��_~��1�?�O�<==q�*�<��Ҋ�*/�zC,A#+H|QVF�X��?@ݔ������q�(�666�KP >ợ�#��Ν;eZ2��q�H���Au��mr�8�{��P��˗/?��㯼���w�!x/������]�pL�(h��j��J?ť���9������1ae��.y�����5�x]�$3�VM��*�X8}�j�uS�&�6d��1�����ܫ�E�b'-$����l{Ҳ4V"���Ȩ�gvV-y�����+Evxx��:�yꩧ�⪊v��d&��49� ;�+u��C�(�>�/��|��ȹ��#ͪ?x�m�i:���Y*1,��D�S5�P�2����O�W�}�YЇ��{eV�P����/ڢ-�#���Z�E��&��QeS�̉:X�GY9-�	���D��'1��\��O��2sq����PT�s*�q�M:�lR�}P�<0zBV�%��2����-�o�ҝ1-P�i�[(C��k�}_W�E`P�P9�+f�O�W��/����`R����#;wz2$Cd�����t�Wк-����I�< ��h�+���4����LV�I�LH^
�=�,CVxGi����uU!,����+O���#�'�&QXe��t<:>*�Kc2M��aԏ�����xrH.*�F�s2NmV�G�2�����Z�z˽��X�6@�EQ���|0��y&�JFL�sޏյ��]�}��8��f2�Ġ<%ñ�Ku0��wwWVVN�J�����`4�8�#?�(M'�� �%���#�lbX�3���H��B�J83Ѯ滋*{�.yQ�����������IJ����/g��ݛ��P>޻G^�G�;�}mon���c�D���7�*9X�w�h$�"��[*�}��#�`��S���W�zub[A0`�Ҹ��e������??Q�p8���|��x����Zo����!X:<?���p2+�ܽ���_�җ�N'�"���rw0�������;?�.\���ǿ���/��t����7�7�d��k�э/--}�^�����w�n\���jem������ڱ���zתs��k���.�|Ius��9�J�@�N��:�M�3�ڥy�Ǆ;�7���m �?P�u�A�\�S��5|Y���s^~���iQyVr�=D\2�l�|�����6·Q9��`-*�Rs.+$��,��W5�	�p�5NKR��q2�~��yJ��"��6XB�D�ߔս�n�ҭ+�ț�9?P7�}��_�"�ҘD�H����4yv�>�}��R�W�<���xs}eus�:��ｵ�4��8�y�Ng��\�$�OA�1@���x*:Ѵ��"�y�b��DA>~��ׯ���U���}H���3���D	���v��v��uF���P��h�v�-|�E[�OЄ؊��d�y�#����&�9��K���[w>}�}]��maw[��Ƹ惾��C��4sD�毹�A?��*'a���L�:���R����j�χ��aδ�`���QJܷE�f��R���PyU"Z�3_��	��,��t�K�.����|�o����x4�}����17�<8�aZli�:�Y&�{ty������`{�3�2�Q��8����&)�-?X'gFD -��Q���@w�퐥59<9<<ԍ�ƾ��ZZ/��s�.�'��*��:%d����$θA������t8�ǾTV���Q��j�]j5Q�l��Bs����)	�nzF�ߤ��˛7o�% H��C�Weuu�>������"��{�:���u����)���5�H�� f��B�,N<=�T(�����}	˕Z����GP
`�ݹCg�?<���t{\l��uR���JB�Y��Ic��Uz+f�x��٘�ёaL���۷����/����iX�o~��4���k#�x�^��wޥ���:S+�چ�T�L��/B��rT��F�����WRj<����9�X�������!t"1'v�n3aȍxN	j�.��7uS�#��u�
{�VU�%�xUT�/�� YrX�)�Z�F��N$���3Jcc4�t��8�0Mc�W'����v�������ވq �dd��=k�:�d�wi���)-MW�'���h�\Y�D��&	�m-8YZ�'l�xs4����sϽ��˨ԥg���t<��pTi[��s�l9mdg�m�~¶�m�>A��{�23��r�Rǔi���������N�7��Q��*..���#(.�ݭ3���S��e3sG���+L�{ls����Ĕ9ʰ8΢d��@�Ԑd"���;�@_-r��X�*vg$���Lz`3����ԕ�T֘`�� ,�i+m�_������j��]�8�Lvv��E�z��{G'ye����4����卋����ɬ	�w�ڵ���1/�c?8Ms��q�
S��%�M�L�f�4dݘ"���B�t��>�̍�<C����ܽ{W'd�3[]utpD_]^^:Tf��8�AK����I��4��>�����~�uW佐z2"�e0�h�b�=ͽ���k�-�O�͏,��C�	��PχS�OJ;�F����`�z�$�O7�CTj����k"/�ږ��ʲC,R���a�*ϊʃ�KG�o�8rUe��CU�#?�u��;:P37r#_��)���`9ˊ���K_y!�������;��?<^�u�~��۷���ɚ�,+�p�fIΰC!
����-�B�^D��k~�K�mm!}D��
������h����og�������["/~pr4:8:,���w����V�p8!�W{>+�A����hPeE^o�^^���
�`Vi=�g���I}����4�k �;�:+޵K��7'��j�qFi��A��g�(�C�s��x)�X�J�q�
�|���:0�2/�ҽ�˫�6�o�#!��n��a��������s�u��y��\���U�ڟG���Y�U@��-,$ř���lA �b���>;��+���E�}�?��9��V6����Z��R�,���,\ż����^5��֢l��1u�B�S�e�O�*��N�qD�����;��VW�������q||\�4	�a�A�K���JN�����C~���s�����^���B��)˄}��+}r}̚,a-�*1QtW��Ƿ_��_{��/n\�`����VyVTȼ�'��
�پ U;H��E[�O��֢-�'hm�Tr��aH��Ĩ)��	x�*�pT���=T�$��b�K� $(+4Y?mI�s~ P��ϲ �Q%=��u��,���k�[R�C�,zC�r��6J2�wZ�Cո�E�>���'��W�9�ڐ�HĐ]{��E�3����P�w���c���#�(���u���}�Dv�S�����---����5S���]y�^�GH�Y���t���F�t�����p<���A���x���^{�#N���}F����m�.3W52�V{@6�Ѻp����Ν;w���O� ��1U��L�h�=�����43������i�b05C��R�i�	g����*=�3`����z'˼y���"�I��i
ܠ��Yֳ2^�]D�9i`~˲ruuI�6runܸ������T���+_�ʕ�K������7�J����"S��s�-8���k>w�5���2Qt:�~h�)��0��W��{���t₫8�R��޽��;��T�z	�GGG���hr�^XN�Z:;}�l���[cW�4������4���?x�7b0���}����^�����_�7��QǺ�H�/+�?e[v�=O5�V��돌��m�oM^�{w�ͣ����L��5�m@��Q1�籯��`>��U0~U0Z%��l���z������v��D���Ҝvge��,1��6��Ɨ�^��J�s{`�GN�G�(�U>=c�/�ړ?S�9�:�t<���[���ݻw�%?>
����~�.���y��s�A�yss�_�����vf�$�&��� .lюN;�k��S����h��[p�L$_�%�8}���Ep��V����4�Sr�?%��\,��ԥ�4���Y���޽c�
��K�!cQ�^y��C����X7���੧�����߅�����h2Xά1���ּ�椉!��Ugy5�l��4�V�	V�}21�tzr����R�DT���ŉ��$7���������H2m���D�>��'���_xv8%��A�͝�4���a�$��T��˷�����
=��,_�ݏ�?��:�ϾDW�w2��Nm��D%n�^ٺ \n��ޞMOE��<Mg�=P��{$H�3��rol���d5Y��Vȵ\�!�3���\�Y6��Cf\�^�^���_���k���c��7�\�n\ݻ�c��v�g�?Y��Q������(����h��q�[�-���~�P�I��"������Rz,[�u�a�P~矕.h����b8�eEGC��Ӿ��1If�w�7V��^����(˳.�����JClLEB(�P�d	��
�_�D�U��$��lB7R�h�f��QP����h:��`-��ڻ���V���u/!�nce5a>}.UUyq�||�n���ҕj<��;��B[������DA��)k��3M]Gߍ-�ݨ.gE�,M��������W_�9:�u�٤���`�߼�+��:H�����?N��m���t���Eʼ����.} ҁ2�����U��N�G��_t�xV�
��In\�|���9�}ggg�4f��?y���_��?�g�ʎǇ�����&&>�:6+��?P�*A��U��i��|�M7��8o%�lFk��a���G��s4��m>2��<�3����z���N3�DLxYz,����G�"�����pr`xE����gYit0���t1�N,�C^�ȸ��D;xk��������l)

��RV�b�G����4N���|��|��ʖi?%�T������w��
!.F��g�=�3�dGscU+�WgQ3�2�0� ��V9��i�\���LG:�_�ZYi���YID=b&鄜���3F���*iѧP�(�J;q?���4+���g��2w�cϋU��&�Z����W����^*L�#���L�w�D:�\�8�i՜<�|<ͮE[�E{�-|�E[�G4=�����---����\��N��y��(�Rj� ��f}`�˨��Ķ��2 Qj������ݺv�} ��i���b�����ǅ�� �S%�*��4MC~�K���T���"E8�[�ت��`7G��հ�9���\�&�e}I�}���"��y�f�p"���r`Aԯ�%s�N�~��]2�m�J  �VIDAT��!�UʊZlPJ�4#TA�
�a��p5�c�pܠԄ̹��xc��q��ԄH�����ҡ�Azwu{[j��R���� �0]p:F����Ȥ1��-���<��{�i��6��ǰӴ�l+[8��6:���1%�R���z��͇�� &4�_y啪�­����E��N���զ�}��ko|�����F?�}#���8Űzm�����C��h=gg�:������jw����0.iz��!N��/~�����g���_�x���>,7�2B&0\]^Xq|
3Om#vxxx��͓����t�˫�tw� ��6	���k���q��I{`45{Q�+R�ɂcŪ�t*Q*����v���U�g��qm>~e.}��yw���}.ԧr=�	��!f��Z^�E��Vg{���s���B gJ7��x�/������ ��Ɯz���S\Țs�/��J�-�#(��h"�l�8��%!���N�Ѧ$��9Wl�
���M����nܸ��č_|�w�:9�y�sf�l�Wa��<����-ڢI[�Z��h�Z˧�_�����:�$��<�V7���N���GPL?	|�z:��n�;����}��iZ!�@��)�&�lee�q6]VB�����!��K�1�D��a\��Q��������x�k�[;C��3XM�a�)�D�T9�E!����Ҫ���xډ=#�ammW����T��9IAa��H�O6�jq6PJ�i&�Ж��: ;+"��4��I���*=�@�~p<ɫ�� .R39�g�1�4N�"�($Z6��dJWٰ�po��5���T�Oc�i��Ea�t���H)V𔣞��,��[�i�ϊ�ޑ��z��$�y��oEI��JS���MjÒ|�*����ɸ�8�W�1uKY��q�/�P\�3�iۘe��C$��'Z_�5�±s�����ޑcVE-:K���/S�
�&8�	Q\�W�鹺�Z��چ���ƚiTp�
�8��8W���8�L�A���`�l��VL��t�Y�s����~PU޺ss4<�׏�bo����	���dmN��O�2Ǝ��Z�������7�w��dFA�^59xE'	"2,����\�X7�}񙧟~��r��O�������MZz�G{��IH�d8>�#�(��A�BOg���Ĩ�Ѥu%��~OϦv<:<���g�����w�z�e�˳A���(ց?O^�\g쓯I^�c�S�SgCl�� ���O�i��3�Y�����Ԛ]�j9�b�H���ì��f���AM�f),�b���*p.M��2A��������z���u���JE���\��wZe:�2��`HӶ(˼�lg�[^���1ai��s��D!����۾i
Q2XI�����M%�'(��g\�`��$ȥ -XA^���Lۼ��#�ޑSQ�=#ЇQ}v'���5�k+�++�<F�Mӳ#�%I���`y���J�*M9�z>=q�o<� Ho��|f��ŠߟEQ@`�g�0��01�'��vgU`�h��h��-|�E[���k'��?��E.��\�rB��Ġ��!�+L��w�����NG�������~�{ߛr#�J �^k�d���#�
$�����G���u��~�����j
x�&
ӊ��+����� �"T����Ub<�#�	1<U=�|�hƈ�'�0�W5���R7n�Fc
d	������>���	E^��!���W&�* �l�@��)�p~(�м����j������7(
7Ge&��\j۷����nĈ�ƞk1�@g���͛���Uy������N��;;;4����'By�o͊���V\���5&(��는����+(�N�|+� p�"o�&U]�a����w�Qs��*��w2��1�t��|�ey��di�p�ZA�S�8u�5�c|��w��84�~�A\OQ����y7N��2@��&I�	g��H�q�<��?�i��2Ґs����O���O^���*��q����?�i���;h=Ҫ�u�}w��/:��OJ�bnj����z*���<͠\����;w�Б�:ɀ�LgOOO������;N��g�j�����>Θ�)]�n0� *8O��$�
x������xH_i:�Z�Z�����"8�jH>�
X��Z�S�>�zn��Ҕ�K�U���p���9�TG�5��y!�=����t�Y�4��і�Q�y��ܩ��\`�R�g�.����)W�y�@����f�xY��,
�$�h&W<�R�Չ>�hk{cc�~�wu,�{Cټ,�����ǌ���Z�E�۴���h����ؤ5��y�*�B��>�q5��e!��8�m���ek�5�G�x�}��1I?�}"�\�ߚ��4��	w�|��"jk<���^T�8;K	�Ш���-C�Z�v�y��5B�`����k B�Z@NU`4=�-��xH]�j~���pU��4�ހY����' ����"��}�B S�sn�g�kFX�̂����L�!�b+䕄����d����x�#�������(��┙�E�*}[|D�eɶ/sY�� r~�a�U�K��M/�����(��Q�f�L#銟��C�ٓ�r�i��ݽ�&�/��<�u�.-�(����3�-A�r��ةu�QaZ�:~�Ș�\7�'Y�����I?�|r�mV�U�Sq���tgC��A�%���\�:�V�:'H�R�+����y�C�-���Io�yͺPL��׵מi��*���a�OgY��U`RE��:���@>+���Y;�ŤH���s���CM����匵���_�㪔�Q�J"�Q2�|a"t�C̿�D��:[<�k]l�_1�bi��w�4�v?�C�RzX�����{o<����}��wh���/�:K��~o<�'���`���
&�k�O���h6=�_V������w<V����Nh�wn~Ѝ�����ӻ��Q�X<&��ὣ�c[�q��#�yJ�8�_ݹ"�X�~D�����H������Z��ك�?{���o�s�\�x)���G���9��j
�E�X;8�G1�Nɋ�G���2���<�e�hz W<<��q��K0����	}�=�\���S�P�Υ���d���c,����ǜ��fE6t��N�h!҃@̌��:Mj�N!XCO��*>�F,)Ks�f�E�X�@t��D�0����i��Z��O�|B�w*2x��j+���c�<���sa���i-��.�O
@?V��@s?}�E[�������h���$��x�j��0��O��baGf~@/F�e�"�Wz�<W��~��ݻw�ݻ����+c�?a�j�.�a����J������~t���1$^���
�-K�[��࡬a͔���+�����slb�+�j! ����g�l7�qe:b�I,EٗR�UGJՊUJ��9	��j�đ�A/~����L ,)��U�p�(�@8<+�d�edL��&��R��*��9���k�dj�f]-{*>����O&����.�f7�^�s�����t�G������2����i�V\k2�����q4_$Ngf"�K���qHhu9���&M������9�g��˝aS�"?lkK���3���;N=-Ū�
Uv��K��
x��t��=�\|e�~?��EJ?���/_&W�^x��u���{4蝎�˿��e�2�͎��N�ez<p�g�����aQ�4�kL�����������/�长����P����7{�1������eii��뭯'��������ߡii�>��>��S��#��ꥭ�����Z^�ϫp���-��o����������*�?KT��}�!����� R�FvV�٘�zǕ���V�ڌc �ߧ�eL�RAi*/+�Q����&UW�[�JȋNGX�X�A��{�����e}1Wd����7�, �)yA5��k���J�d떯ԋ��[�MD��A��C�n/��c��pH���Sr��Բ�"�\	#(�w]���It��݌|��d�	�J^���J|��GTfon�br@Z�g<�xy��>ך���ڭE[�O��֢-ڣLp�9��s�=�Ǥ=��Tf�rΞ�'m�x_A�ݱ"$�c�pqki���kE����?�ַ�u���w�}�L��dH~䒕�DU��YV	ك�:��C�'��PcUWo�,�C����������� ����j� �U�0�`�x��Z�$%8>��jz\Z8���]!��Jd|U�ټʐ/�\�-�Ɓ��q�V*E�]�_�svP���%^�+�{dX|�37�ѡ+"�"�qt�d���z6�#�A�F���p�K�,�h����T�ޖ\�^B�V��覐��zE�=�0��/Cq��PZS��@��o�(<t:Ti�J��N�J
��s��I��@M�^(�`F��p�	��Ȏ��2ŨMF�B�~�ӘT�-��"Q���l�I6�:�����8��:�>�(�z#����jB	��V���Y�&�	��� ;�q;]:�=�!2<���xB��������;�v1���޽�Օ�<�̅�mZ7oݺ{���V��w>�����67�"���;$�e@�*k������Su��k	]�nK~���ݫW#���C�H_x���^�:d�?�}����;�����[w�I���:�����������U4d��>�g����F������N+}:�NO.�W/\���yxr���~�HA�}Z�~���+k��QY������π	��y�;�=�P}�<�ߣF�c��G��q>^��y`����>�%�b�s��u�K?i�������6�$⑧f����)��L���_}8CN��*ñ��)gp�����v5'� ��_2� BH�m�E� �X4ďb���$�ﴉ���A����*�}e5��c8�x>ŗ<-&� p���볘!�ʨ�,��r�L�3��%G��2�Kx�T1#���ǒ5�\�@B�<Lr���4˸^�c����l6���J6W�B�B%ʇ/f���왬��>/�9��'�-ڢ-��m�k-ڢ=������`/���O�6<�Jf`�>'�ވw�N�<������mz��^�w��׾�5r�>���Ȇ�I����Z�����<&�����.�.{R?2���Rp�A��@�e2By�#��2/�XU����t��*Q��u�g�#����k�,�1�ru{�T!G��2�h4MZT��U7A�@ލ,=���Ϧ�=�9�7�������x���"C1�c,K���HՓ������[����ͥn�c��$5��/����#>�~
1�^Q �����gѥ��M/h�#�J�>K2�XB
�NAF�ؓ���^oe�Dg�~cy�����s��j�#08�"�S�r����ZK��j�Wt]<�Q�@T��� �r�8��n�V���������Ԁ��FH�r�1=�ڵ�Whړ#��ߏ>������#;�^�$.0�T<��??:�[{��õ:�薼Hk���ܾ��kW�^}饗�|�Ϳ��_�8����_����������	��O������l����>~�*]��o�C��,�U���/]�DJ��?|�����kkk�c�	G����7������G{�/_����+4��$��^��#C ��)��ٷ�;��!�&X��I�)��,��u�����SO~�_����}�K_R�ٹsg������w��ўy� )fȵe��\��7�)��Xe�27M�V�%X\u&L,y���C�5�[ӫ�IN�o/����x����r�H� fm��`�B���*S��r� �9"G�N67:�d2�/�I}�"�S��Ui'��[����������sUN0@������G�ԃ0�k�Z�E[�O��֢��ocF��ۡ\C+A\��\T�	$�0=�x�@��z!�ǧ�/'�yd??������+o���_��_��N�=�:E��69:���g�� �Br�Q1�vU�p�Σ	�Z�v���䵆h���S$�ą�L�tY�iUXq��rf#=�˼9�w��t�5qlUF,��[�tY&��S�Y'I  Vt)eQz�$"�z�,Ψ5����	��q}xB���k����(J����Gw���� w��*��R�4�B�Q��N�s����i֕���c� ��
�/0�3E���A�����	��3�k�ge3L�Ȏ��R�{m����D�U�^]�r%*�t�`������T6
�ge�J�@K뫐�"��`N�Ғ1E�X�l��*��6��_Էl�V<�d�<u����ՇqFBd����'���u�*� E*�����\M�_c&��6_N�9�p����j�����]���_y���� &Òp�b�O���;�/�_y��lн�u7��O�ã��y�g=Z�0(a�c�K�u>�X[I��� ��4�&�8/�ON�^�XO���(���k+�[4́�E]h��5�A���ɤs��qd?:����t��Ku��OA*�gM�b<�a��6�����[ [�����B��;@����ш��7o%^��?�B/Q��紸K��ρWZ��и3?��z��}2\K�GӮ<`]��=�����P�˖mӈ��N�1Ȍj�\��+S�ʌ)uܡ?Q���W���]�c��z]�	�׼��W���%�u��g�����zzz@���L�W�_CX��J����0eT	�_@�Y�����e5M/#!�����-	9MQh�4�2P %7��F���\f����-�<=�nݕ��Ll���$�|U�f��F�-���[q�!�tT@��V�&�����VG���NgYwJm��M�N�GG�W��n��^AX��{�ս��賩8�X�E[�O��֢-ڧl5���o�&4� [�L���9Q'''dcM����{O���i�1y#�"䴠p�<�R���#	�<�ۧ`� "A�<�4��_He��Y�����+�p�9��3����Mr5���r�R�˾/^@0�든im^��,~���X����;�y��r� 7Jd�	f������u4�P�F��j�.z7�lOW-�'=�Ҿ�]�OƧ�uc9rW��؃0�S��a�,�{QfX����0G�ԉ\�	��6%�<2�eӎ�������Տ��<��p���^�-�˾6�X��壣�����rx�'��Ȕ4穻����l�ш�uY)��ԣ&��]��O��b5�Rp-�Z����}��`����	��#��.ͺ@��������|EOn��9>���V���!j����ׯ{�I/�w'G�t�t��6����bL�a�z��>���dA����q���\����/^�r�ƍ��2m
�%ں�>}`{{{ww��{��+�<��SU6��t��A�)s~��CF�*�o�����h*[��5��\1U��p���-W^h�,�6�%�m�W�"�~��[/��H>�h���=���V�P�{u��3g}����i�`	�1��"����h���o_k��q���CL�N��v�%�J�̛��Z��pu���&�~����������*Y	���:y\����B���tx��
O�
F�0V�
EV.�@G�S�x���L<..��t�*�	T��(ͷs�c�_�jd@�%Z��\r'\!Cn�F��	��F��Q�]�{�	�J왤�p�U���5����q�G�=z��tH�Fv��3O2]�9��N��t��F^����/Y&k}k����~�����k6
6}�	=���*
��F�T��)$1ા;)�ưsf+�cS�+��oq�d�1˕�G�re4;��>�U��YIc�|����eo$��U6/g�R�@�RV��3����&�3̯hK��kn�9>:�Y�&J�/�!PL��/�{i6�sZ��ߞs����:�;&O|��k�K�%{v4걪0S�sy܍ۂ�����9=<�뷾����}�
����:����z��ޣYqac�3�G�Fn}�̉�����xyMu��w ����2ywo������ӟ��̴��t~镟�3�����x㍰����M���p��������M$��}��V1��ϥ���O>y_��;��U@��h��ԫ�������W����?��P��:�Ùj����n@h@h�E���'�D�h4��9�s5���Nh��Oqx
B�g��84��L=�{k8����9u�n��{��˶�[u�>�콫j}�[�[�)େq�;v6�;1R��g�Z��H)Zf�	S���@H9We��!=����15Ae1�g+��ո�B�����IK�G�1��r��Vю;�)V�֫V�m/��z�Ӟv�A=��`��:~{P���5W��o�!�o:��V����[�8��^��͹}�y���q0�9��#�J����B�b��g��p�� �5C�iNj�?��H�<��#�އF�_��#��S�����4 WE��N�I�
�)��[^
�P9~��	̊�>:����P����^�'i�g�39���y�cҴ
Q�p����mk9s��|��W�Ŵ[+��
�b�*�" ��755�/���ܱm;z!����tS�Z��h1dS�qs3�p5dh���%$	��rJ��e�T9l���z�U4ZAQ^��Om�J��@
��@7��ݥT���`���Aڛ(��x��LWz��
v�c� O8&�
K��3�v�
6i��L�ƃ�_I�-e�po�k���[�yR�ّela}f��-7�[ѲV��bMjx������(p4~w�oyƑ�T4Y�*�cH�LN��j�c�1�{�Fu��<��~nh2[�6(0����Z���^�n�c ]�k��6l0Dg�>A�pS8�f_��_�}AY˺�1�=�����D߶m��
��٪U� �@?�;�3�k(���!�f{B��ls�x`�TQv�I3X�ͨ�����`w�0�^�����A���bt⍿�Ű6��T�G���K,��i/Sg��Jmw����I{��Ӎʨ��S@|8�������#��9�5Eu�h����	����k��֭[{�L+�ނx�'��X���~� ��	1�r��1i�Q|�P?q���0�N��h�@������jZ�T�Y�%�l��G�YE@�XX��Fx@Xd��ը�Z���1�*��ᩓ���9s�2sX˙��/R���"��q��Av���[�n���/�|t�A|�����t������?�ӭ����]��wp��)aj�*B��f}٤?�]0�_�㑊��<'�i�x�r��R�(B��-�)��#m���Q"���(���ce<�%�ác�������ߏ3�E�el��;�ۿD���T�LKj�ٮ9pMnZ��������5��8�dP������.��С�1^�d���3�x
��8����J9/˸�"�����i��v������$�U�KB���pf��!��J��͚��6t��yp��.��s;���f�� l��Rd�2��Z^\e��;�q&���g��!�R�Z���谒�7I�:��Y�o�����g�$���kyl��R�u��S%W��E��z�I�.�6�N�pȩ����{���M�ճ:���W!���{ٕ1|M����}�	(���ź%���0{��M��%�l aF��k�?�ٱ��m۷�t�u�FuJ/�1�;SSS���I�W��,�hG<�N�j��=h���i��y^������� ��D2o�.��ww���SN:�������l�~gon�l��K�j�|Y�")�|g�����'��n�ԭkY9�ײ��ա��>fP�Z�ُ��I�'��QO��΅������i������=f�m�a��>��ns�&IJ21����/��_���];�b��<o���PP���h��<������f@Ѡ��*Qy�i�oVI�,e�+Pa�"�YS0b�D_���3�/���h��8jR���g�3��弞1	M0L,��R�bV�N�M%e4P��M�ܛ��~��������kU~�DY1���Jwm�r�l���ZΜ����0F������-r�t�t~�C�ƛ���f�37�y�f����_�h+|D�Z�o�kL�<t��W��:B��AJÖX������.,�qa�ݕ��b��V)7\���L"�Rp4#r�9=Y��Y���1Gu<C�]w�uU^��	��@�����Ѡ�3d-Z.a-���6�yx'����9�Z�&���ϴ�n٣hOT#W�?�Is��J}2��_W�H.�9�j��[<��H��g#�v�1#��K��:��U#K|k�n�v�m�gff��9�C�=@�rcT�.Q���n���q��ʴ=I�����\ЈhvD���J�Mb��	Wp�ZF��	QDǙ����Oz��/t:0�V��n3�O�M�6�=���H�ԫ�������������Q1�\HF_\p�i���P
�s2Ou衇~��VKX�x��\���fK��Z_b�-����"3���33\VQ��bt�o����b=Ծ7XqP�tVQfV����<�8aRg���n�������,�ZG��g��`UVXu
]�_��;ڵ�f�!y' �T��Y�Ω��+m�g�#>cO�������r�l؈8�{��X����=�eN���~]
�����\Y�0�ґ*+�JY���<�"�*6m~�s�������Y����;�3���A����*R�h�!UQ�bŜ��9T��K��~�IX�����gY�C�D}���%�6��lV��wQ���^l�iY�E�L&L/M	��a��Q�I2�p��cY���0 ?%i�:=�ӟ���S3k�@h:��ލ�Q�N�zwj��U�<?�X�?�$k��k����:B���+��'���!�b7�;�c`ʥPL$� i��:������#��,�l�V��\\�<���m�»� �{4����Q�7�����G�z�$�8;�� �o�� '�[�Y\�Lb���+̢wk�K�Çb)Oٕdej]KN,����W��)�J` �tR�9�]�Z�^��ܸ߆Hj�X���g?����^o�ڵ׷m;�(�L��H	�Z�Sِ��5o����wE|�./}<L����w�u�U@���l�!r�V����4�v���F�Qq�0�"�m���>���$�3���mz!�/�����2a�Fh�q�F�v�i��6�ဝ�w�Yn���c��c6�� �����hd�3S)>�U����r�����+V1P��D�I�����IId�񃽘�+���d1�^3�
���}
�)O&of���ց������ꃎ9��~́�ظ���9��n7%���<�3��������h��m�/��A����Vy�=I
�l�ݣ������$RBt��r[�dH�M~��4kب�]���k���	y��k�&#����V?������C��z���QZ/��6����;ŝ���8V����*��E�Ń� �F���6�1֯�h8��U-A��g���氖3g{Ɩ����NM�>fA�xE� 	\��$��u�;�-[������Y�$��|I�X���\��6jI�H���\&[*��G!^,k���m��{ُgg.�l[nف(
C�����:���p؃� {�.NT�����^V��g��m%}*օz�t�,g��D��� Ry��+��>3�CR�/��X�e�
��P��X���sZ�Èz�9M>�k8_�$YB����E�U8�֒'F����^�H�+��b��X��G����q��q��9uf�nݺ#�G$3�e҉j�����9W0��ʥ��S8��}J��!��>�t:^Ɣ<Y�zI:��5�'��E�@���5�-z����S��)��I���Ƶk��E*ֳ��ׯ�v;��!�2??�-W2�[33�*��yY��r��[��n[�OD��S~=�0�I�O��a����p�	0&333| p/��d1 č�����X�.�6l�PLP���O�~��,�#�*����ʢ�E\ ��>��Q��{�j�[�C*�}�A��D���^P�!��X^�a��L�0 � _���(�5C��Ga|rz�+mn�ej�c̆��+�Z�/��ԫn'�כ��4�5�?i�k������HΜ�}sX˙�a�KEFb�ϏC�1�׫�*Q�K�x�*z�S�dQ�+�cn��������o߱-��3?e�E8f/��7h��	܄�D)��G:`�P0�jkD��R?)F�1 9��9�ݷ��F�E8`<Ew����'@�Qb��;s]�ыj'�AI�wBI�����I�c(����s���;��M���n��ZvS�����c�w�c���lJ�i���.��B�85���
,���oC,�"ƈ�Ps���q>��z���^���)�@}k,����C..!|��.�&}$'ՔM��4�����¹k�t�O�<�!)�p(�$�y0�A�V�HW���!�Ӗ��-�*�LRb^n�{j ތ����:eU{������V8U+�+�[c٠�U�Ԫ�Q��+$E&�͜�嶛�o���oܺs�Y�պ�*;7}�%i@)�2�PvMP�M��B9%E��e?)�>&v|q�IaH1�?�d�- yH��s+�2T��.E��Qn^��QpB����Y(����(���7������Ɔ��$�����;#x?��;v�h�i~�i�t7E(�!rɖ��Fl?$EX�%?]���`���u���׭�Y�G�[��Z�Ȱr�Gs��J_$l��)5�Îy�"�D�4���U��;n���ظn,&^�ְR�O���|�k�y r�K'��u���3�n���$W�~��e�5�8.%L~`R��p�j���3��/n�4�T)��J���|���{F��p��Xx����0|X !k�v�8��?r`$����+}��:�h+Q��u���,��hk����WP��Hu��{.�i��S�c��MWO�c{c�Ǚ���9����=`��Y�cq�DQ ~ �����>zӋ^��u��.�p����ܵ��D�q�H��R4�YF��&�����{�����b৹pgAge
���S)�LQ}���L����m]/��R�L@
��<s���}f����:o#�
FQ���2�F���03&�� E�K-ʘ5zw�((���Gg�1�1]r�ܘ���Cb�U>�>����q�1R�\�Y2�U�ow�E���!M�#��&A��!�]��5r��$���C�eF���k�q�n������m۶�B
���,����c���41��/�?b0�þݠWK��q5pv�M��VEy7~%�҄�=�A��O;X!���u�j��Tp_�^s�������o�yǎըm'�]�v��v3��(^�&M����>}��;g��W1�A]YwNSd�V��.%�4�
c�E�u)r�(�{�^x�)���јn�hMU���S,L�TM�� 7oތ�C�_����a�DHWa{�|^W��
r�zR��q�B&���1U
�`�6/��r殉2R\� .�Qp�^�٭�j5�U<�[���ϝ�����`N��B��Μ9�'�a-g���u�?�(����>+�~ܜ�=���[a�\��G߾~�WͬF�E<������A�2��iE�����9	m����Rȹ��s�����QCW�8OI�>��`˛΃4U 8[�m��*�����'j?ˌ���W~�� �]�#�]�F��g~��`�Hd)�?O�4�>��E��x�8��7��)KgE���)�L1HYe^�B����x���m�p/�z�����^�~�k>%�S�2�� ��&��p�<��<��vh$���9^gJ�\C�i�nj�D(Oy\/���C;⤈1�WD֒�*ƹඪ�U���0e����W�n|�E��|����ktCJy�OS�����(b�����}���Uz�IR�S���j��3̏��c%9���nZGYě�:�8x,W�=��TU���a%&��*:¢#��,�{��[E��+�D'��$�@J�8�I�Y��ǞҞ�d�~{C��}�ٌ��[��!jr&]�m��~��Ɛ�b�zP!���0�C���ɱ���
�0ߎ)k����1̊�/����X��;	�'z��f擰��M�]��a;�������s�v��c�y��ڱ�<0!:]^F�
�)�y����=�q;w��rZe$|�1:j�Z���h٣�?]�0Q��(H+BZd�@K�,�x��;&���@(Q��P�_��r��H�J�gd/Fפ�D��"�b�Y{>�[A2[t̓3g��9����=luƖu��'1a��?��c���[ny��o��o~N*j��R���(�9���,f�#�&U�~��OXK�`x�b�fj�Q��Ln_��ȷkU�HE���[�{0[@y������=�����?���nk3^��LOOwҴBY9��t�s��^��;W(����!U�z����e���h��aܨ03�T@T@��C0�ܳ��dq��	�Z�.��Ԁ� ��|�2��ɨ�2�(t��HŢŪe~����"��<�~�ܞ��b��u����"�5̡�JJ��R�!mn[*v�2Ԗ��&�}C)J-�r�yg�~���\L�&k�~z��6\����)J�ɲB�OY1mM��Q~�('%��a;Y��{Ɯ"c�mۖt��$ź۪���Y?�MR������Uy���Ѱ��b�Z�O���۩�h�\圇��ޠv��8:J��h$�4&���H9��>��O9�ݳ,l4�Q,�hpXpA��]��kY)Щ�j�t�I��0`��F#K�V�o����;�����^~NTZ���0���h�**,
�?���2�������<�H���DՊ�kX�ə3gw�9����>d�~�5TI3���'ɺ��Z��ɧ?��}��߀���6U��C��Q��!��ۼխU��T�V"QC��F^!gG8J�B���{Y�1{j�hA�HAߴ��{�S%B By�W�Iao���G!��J��l[3��1�K'9��8�� 1U����T�H{�@����!�l��4왕7#@֥ ��c��`<Po�G�D���2@DnR�2 z>ʍ)��0�\TY:Ԃ��X�g�?�B�!q��~�"�w6�oOE��`j��^�Ie�
�r>�T�6�p�M�ݬ�i8E��q��Y=lS+yT�xvQ;�M<��t�=���-J6�9��,S�J��0@�F\E�5�l6����[�㇩^�	28�E��#��`�[�q��C���V=ѤƞH���+���V�s���J�����{O��ʍY�3in�L�t�����ʁ������(;���(��!���|�:����뙦�+��~�'&Ty}a�<Q�����wܱcǎ-Ǟz�!����?Z�V`�,�ш�Tb�a��,�nlY�]1�&pkL?#���I�0��`B�'*(�=.(�	�")[ք�D��XG <�ƭ���Y�+YI.��
����Bk�>��"��A�`g���ɇ㺡јt�p���^3���9����;@+Ǆ����4՞O�%*�s�y�Cһ���n��?��ޡ��Z����{�w��:`~�����K(�`օ����@[���6W��x��K
Ub��$k6����צM��,kP�����Z�E���,GB.3cZst"���Q�}ص*����L&j,�#��u�Bd�F��h;PbT�L?���d̺�]��#M"c�QH<[bH
΍�3���euV���8Oh�Wyq�M�Z+����b�c�_�sk'[�����v��O*[f�y%�����(��*����aJFVW�U�?iK9BL&7�1]�k`q6NqbΡ���(�GN��t����*ɕ�$�����%�J��A\�:h!E�%1�r,FI�0'���ՐN�w9cL����&��X˖�?9����^z�>�����u���� ��eqB�����cwQҡ&�^D�,u�$ĸ���5���_ :\�S��5�3*c8&g���yY[����o�"�RTYXRʲRV}�/�t�p_��Sᨡ�.�A]jR�-N�\����3g{��r����?{�b*Rp�� ���k�e\3�����-G�;��S����}�?��*8a-�e�cw,/2(D�t�o)��H���ʮ�_Qj<�̀�fE�~ׄ޳x�ǻ��>(�S�8G0���U1:m�4s�m��� ��/U�}��m�Ս`:�����H?�a�]$�D;2=D��f�4���7^g�r�j�x>��E��ēp~�a����_�(�^���y���)9��B88��#�}��P=[��P�*��ʤ�j�ʼ��kX!���.��-gR���HY@�r��]���/�>�i����QJ�a=;�K�ݝ�������/|��1f�:��V�&e��ŵ�4%t�4E�%i��?�Rݘ�zh���{�,�R�Q����B+�"�bM���w8�u,�M>b9}>|�g|�UblbL�l�a\�%��|�2-�$Q&{�vT��#@�"��T�o;
�9鲮�(}��	>���'9����@}C(d*��c\C$��J���i̪Hwm0��?�䣎:j�)�NOO#He�о�d�$*�UZ�*����͔R�hAp�e^}M�%��g$y���S,B�����B�� K��2+�de6���O���B�\�y5�p�F���Հ�ߴU�2�zh�e�x�G�NO�2m��Z�n�̙����r��������^]Nũr,�i�(4��S�����c�]�j����s�W�G2��]^�PS�)Q�M����ж~�0�P�k�2�Q+8�i�v�`�wx^�q�L�`�BIi%����۶nC�f��o�MV�+�zX�[�;t#]�5Wu�#^�Eɛ� Y�Tc�\�� v��8ʨ̑�4��G�L5@D�A+��y�(G)�PE������j�["F<�	.Yو�|Ȑ-?�H���3'k�B-l428�HҔ,%;*�d��*�� ;�:���{/�r�r$�b���P��m�G^e
�
4������ʨ
�G�R5�<�ZsH����Ζ�h��8P-F��&b��-M},~����Š�9��fgf����?���Hw��$1��4�%(N/7PT��YKQě��J%I欘������.粴�L�
�U��W�*+p(��7���4vdF>�楆W�2�wc�۠��c�!�_ř3gw�9����=oՏ��u�ի�O��D����}?�y�#O=��������Db�~��qGV�)�4����*�6qb
�X��0�Z�Gvz�ײ�X��c��#]xf��e��8�Dm��zD]P6�?�cS#vZmz"a}�]���A��h���g�	j���SG�SzV+�H�F���L����5)݋z�YNutY�����̡\�"Z2ϒ�zR �!�o���2�a=/�է���>9Kui5I|]wIr^&0�i�u�r��@�4!�L+j�K ���0)��SҌ*�fɈ'��(P"9��p�K�1��0�q4�G�1`��h�IR���es7ĳ�
��8��*
@SqVWP��[���0$���fyXB�#iS��,�=�kG(c�F{"8���`��#�U�~#��80 ���&�T������
{4/p���.1Yj?�@e+%9�`��Z���E�Ѐ��9���%I�K���a� 5�����$�UŨ�2��\
i�WTC>t5΢�"��|����{�2�ju���K��$=�L-�`�(��/���ˬ�?��m޼��'?Ƴ��C+hA��z���h�<�|�`�hw��%����� )�^��j���YĊ��R���))��
�Aq�����[m�fQE���C�n�K��07���I���� �3g��sX˙�}�Ɩ<�4����X�'<�3:�k�����_(�h4lB��ȒϩG���%�����c��x�x˶n�]��H��Hẏ5��4=��C�]��7���o�V�ɲ,�h:Fq�_�R]@�.<��߇�>q��A]�k
�ܔfb�n\�eC��@O���=��diB�STC��F���I���P��F4�J.˔�ڔe0A�N����oC(������þQE�h��RZü��c�ڞzm%,��!�j�Ka��+DiYc����xE[
�s;c)�!߱����f��P?����9�M�̭,�EM��#�"��A�ܨ� �[)c���.�B���-e%+K3���Zc���x�y�G2 @kd�m)^�.�9H©��j�E~P�2���6,��^����y]�|*���e�N��tb�}� �v�ӫ����>���<�H��VHu�
���c첩cM�5��d��R�k=^�e��KΜ9s�氖3g���Z�|�����y�T��ǟ�����G\~��7\��xڍ\L9$@ZJP�TQfE�Ԥ�/�8��A�V *�U�D%�r��L"��$��(����4�w�1���k�̀o�ymK-�o�}�_Υ������̀TUJ��-��8A�C�o�6��ܑG�RI�v�2	�B1���Ǖy��93N�	����:�=� �[k��:�^�7�M�c)��w1�(�3�#
E��Z�X�OK�VQ�aZ�M��i˨T�>�S����iL�f�1�H
�w]�#����iBE�^t�G9��-+�kf`��IF��H�E^P0Ld�4�`�m��ů�1~Xly���^�-�9 )�B�"��`tyu�
�|X׾'����2�b`L�0dI��X&y�x($��g]���WohR�0�&(�|�"6��`�Cٔ5�����&Hσ��(��H7T�@�a�0_d��������Ƥ��@PN�Œ�\y��7��c��WV*�9����r�N�^�sb�����������Z>Y���4������𼛠�_�
�J��욙�i�:�μ��o������q��c�ǫV��u�|{��D5���)�\����:��up��Q+�D<J�k7;p�̙�=hk9s�O��)M�"E����q,Q�,>��#�l�2�s�7ܐ	Wޙk�ۅ�,��ÛӪ�/�O��Bd����1����"؄p��e��C�,�k���i�&ս��[o�5o���_R�iI���c���;����O�x��'���礉�U��/����
�3�Wac/���ļy=�����pd��0ښQ����$���)�/,,�� ��?��GCTO��:�;�s�5ֆ���	�%A5b��f��OS���Y���jK�DS5M��[֪z�yc~J�^8��
72�gI�p���k�Y��zh����7+��Sx�`�U�2�Cz�*Pq��
x1Kpv|����SY�����!b�9G�
�HJ<k�H��͋TA���I�5��f�tm4I�$�R;�n��YNP}4*�E��@�#����-+���b�'�h=R[��T-�HT�|Fv.tp%�[�w�Ƈ<�X�f��l��o5����6��%}SY��/��ǉ.��dǝ0��r���]6���9̰ۗweעt2T�T	Oiz�`�j��9����xԃ>����o���l�ݹ\�<%A�qG�����K�: �G�k@�X#5����A.���:�6���Fxn{g?��نӿjzv�:Q�B'݉w�S�_j?$�O`���@�t� �������e-�����=~vUQ8����[�ʅAo�#k�LW���i�Q��"15�����L|�6DV1���~��g�S�=G:Bl!6�����ιm?�ygn'<_���o��v�1C_削c.�%1UbE����Z�/C:��ڌb'��4��S#kZ��mm���j�Pqī���5�S���g�~$��w9��jDʒ~[$�8Ԉ�?C:��� 3E�_�z5L���<Ҹ��u�-i*X�M�4ȷ¨�"jΉ
!*�+�Om1xk�ZA#���ǧY�V�����ff�V�ܜΓ�ߏJ��w;xd�V�"�$��4�Qʋ%]�mQF�1E�^}�'- 4o"%���lV��zuT_���Jǂ�︇��hL7`NaEv%��N>���<��?�5�6��(Oð	��"��@(�o#�VP��e�BF�N�]�x�����r�Μ9���a-g���U}*_=�<�H,�fW�>��c�m۶�������$a�B��|GC�6K��V�F�R�T�.U�Y��*���g5�%���~����w���.��'&�_z��$ɡ�
�tm����#Fa��X�y{�:��j�9���KQb-Q���UI�U����,���ãG��/�
$4�7n��*t�=�)XՂ�se䏰qf��~��R��8����J��`r��}��E �����|vv6�P�N��{A��^ZnEEj�x�ƛ��EƑնN��E�y���GY	Xa�����Fڑ�V�0ջ���"̆��jHڱ�(��W�0%�Z'h1�C�c-���a�[�e8� ��۷[ʳ�(Od��߀�m��E�т��%d/=Z9F͵���<�r���"��ʎ�c�4�y5<�U��y�ؙ> �$��>R�i����ӕ��[����O�����`NKxV����1�W��X��U�O���Ы�*>p�U@�!V��)�4h5fffڭ�q����#���$���g�Bb����ڒf��������9sv�7���9ۗ�آg����sP�c�
J�t�S�,��AE�vt���I�7�މ'��\�Ul"A�U<>�.�>Y�[���+�K�؆z�U+X��h���3w��7��'?Y����κ�>�h1��`^`�_�C%=�'�����Y�o��{�dh6��UM<�
mbD*J*������i���e�S�#�,�z�ֲf7��Y5b:a���~�I��*̂�a$��#���	|���}h�"��	�K�'��=�i*��dY2{P���C:� ��������&v�H��,�A^�	�[b�(��k�)b~�\\���&�N�U1��5|������H�2��T$
�4��fӖ����
�Q�����Qp��5a�	�S�e(���Y��^=�Tp��"&�������S?�A`$�Z	�a���*�"�z��0�H�(j�� @�2
U�Bh�Oz���b5!UCF}x�rb/ϛ���#��=|�פ*�-����J�H;L��2¶�H��8��Y�g�y�+��_W�k�p,֢폁UW��g�X�[��jﷱq��8$W�	�/���X�Lk������Q��`�"��`�`͎���㻖a+�ct�̙�=hk9s��Y�I|),�Tf,e9�z+������-���N������D�i����1�P�@Ԝ�°��W<�,���Z
ِ��۷�����|����)��/��D��*p�D�����r�-��t]�pay���k�tU�Bk�̰)�3cirL�)T�-g��u=�������"�����;�a�^�|�cE�"REP(��[:�����o���ZA�#�(�.v�s�L�����En��� OP)b��S�K#v�ӕ��ޭ�U�݌��.�E�e]=|t~5��!+�ƼX��p2�R'*�aëK-(�*���*aX�Ac���T჌�h���Zz�bbz���P3`v��p�B��j��!��Ѳ��xJ�¾aZV@�2���=R��}�#Sj�/?\���GSӳ��pn�XɡYm���>�*��6t�t��P��� @��A	�ݑ��P9��p��U�V%ac�ڵ�قe�Ѫ:�1�A3J{j�<8��{`�9�˙3g�.sX˙�}Ɇ$���SK�O9W
E2d,Ce�D�2XS�9ډ�>y�u?��̲>�/��$TX* M�n�ϛ�(ЃoU�^����E�4���;��o�,�>`�+���|���`�����P���Lz�:0�n#_��b��3���R׍���.-tDy��wC��� ˌ�}ҁ��ef���;r�w���j����"��$Geg��zd����In��J��?�8>����=ю���ȶ����M2+�%�����U$�����}��c^돪%��މ=E��X��%6G�6�N��9�Z�Vd5�7X�HǍ돲X���+�4E�� �R9�:k�RQ�B!���}��6�KKW�Z������yJ��{w�l�0���9����R[��Bֶ�y���YQ?~�˲��5�b�9{?�;&	A;Q\�%�!��$�x���#Eo$a�ME��4�+��J��V�=�Ǎ�O��0b\�I>䪦�^Cq�+�kt#�7`�X�^�>�6UT	�y�x�	�|�0+�q�0,z�4�j���Ϣ�	?���Ryd=T�31rr�V�>c��ͥ�j�v�)d�?��˚�C����T+��z�'��0_+]'�^ϽASE(�����������3gΜ�O�a-g��5��GQEQС���ne�>������hw�*���zl����'q��Y�������x��/h6��о�=���kVwp�Q"����T1������;�4������rȇ���ǉ���U���!�WR�^ŲDy���ӎ>����	`K/��{�Q9��^�
ǶMjgfX�M,��rO�Ǫ:�˼n�b��U7 �*�OM�Kb�1�U�K@�_���	^:=o�̢:�%�;��j���K�?�:㫡[ڝA�k9s��~hk9sv���u��]km���4���q܈�����nS7h�x�/x������f�=���v��ыNp%��r��q� ���^ڊ�+�����ǲY�*j�2�X�Z,��5�f��w�&;�N��UF���L�G�g����E,�2�}= tla��C��Œ-LZ�#��.^`�G�^w�fI�X۵ �P-�G��]R�p�̙�{�9���ٽ��MrV*����F(-���W|v�Rbc���N|3�Ʀ9U�Ykא�A�f�/�w����D�T\�	3=�$����(����X"�jI_p	/y��bwVw��]�d�KYr+��a3K�h�ƀC%Q�Y/vCY{C���;�o+��'�]uhG:`'�N�Z�'a����%o��5��rD������m>��Z-C/���Èb6�O��\���R�,��r����4{�v�9s���fk9sv�4Y&E��x�[[�7Sb2aB���"�N�zQ��<{�;��CD��!�j|���f��Y���d9�%��O��h���|�*�p��	{�ح�������ewz��P��8�����6G�s�5C�����ޟ��R��7�k����l�ڙ3g���氖3g�V[�,�iF|����\T��J$Q�],r���j���B����=���<����Qb�4��߁���4�%�}�JTP-��_A�����u~��cB.>�b�&G�q�e<�㥬��2�� ��
`<a��$PbW��&�sIm��?)oj��j�:�����/�g����%��V��f�����j�l\��d��������9~"���XJa�,����u�9s��>lk9sv/�I�# j�L�]���k��d�uf3O���a9_�O�y���T�c�1�-��C|U	�$���7�� �>Ok��j7X�h�:�R�1U�YD?x��	B���#vO��R��L�?���=��������AP1���6��M��fI6k:Wi��-gΜ��a-g���[e/y0	V7��JEZ���R�
 �61�߽��=v����o<��]ԙ�����XG5�Q# =��6���F��qw����=0>v�+�~AmY�)����>D��u������+<>\�a�-��o�}���a5��i�W��>2Μ9sv���ZΜ9�h��a��^�ߋ�H�f~~~:I��V�$o�{D�Z-�U�$~(��]a�(gΜ9s�̙���9��̙��֠�J�1W_2�
E�!����5�����9az�;��_��7er?OF6�Ӽ��Ʌ�[����bðQ�~D��U{��
ٳ��-JLڽ�x��o�[s��p�:{{�h���a�<�J��xZgΜ9ۍ9��̙��L���՟�7�I����]�x�Ϛ����V˛i�@d���V�ۦE�N*�{�3���p]x�3gΜ9s�l��r��^l�^��,���\+m����Mv����.��?T��i�(���(`������m���oE S��G�%��'�g?�cV�[b�ڊy	����'�<΂b	{C5�,���௽��TD[ʕf��e�Į��=9�{�V������?˻�}��9s��n5���9�/�^�*+C���3��y�;��=���р���_�� ��Z{؍\�:݆����TX]��>�Ef�r�+R�v�̙3gΜ�G�a-gΜ-a�G9�/%�w?O2����ͷ{�w���i�Z���v��F�`���,��(�6Fh��F?�)1����}ņuǍ��c��RI39��`k� vo�޽�S�Ԥ�Gr�̙3gw�9��̙��f�eڒ��AKS��W�
P��M���v��j�e�4V�%P�5�s��eZ\��:�ʙ3gΜ9s6��r����}軶Ӽg�Y\I��2&�P���}U���#v�M�ʰ#W)������?Z�3��jJ)�!�u;�_��c/zс��0������.���
���M-K!��������������H�}�B,��1�;?�v�n[��N�9��x_Z��F��P���εT�$I�e#��T��,��K��=N8|x��+��Z��ׇ������.�}�x*gΜ9sv���ZΜ�u�K�T���iGK��HS�����c�{^��J�秦����w	�Gh����:�����R�ZZ�4E1���}�	�ٽ�"�~��3gΜ9s�l�氖�}�����g�Y0�>�$��$�^A[j�9.+�x��� �j��?��W<�����Oz�;�����F�~dD��E�-�B[&
�{�z�ϴ���O���z�s���k����z��0wyͅ���㹇m�<�أ�<i,�����W8�̙3gΜ�%sX˙��n���e�'mu�]Ҍ�*���ã777�e��� �D��5�ZX>���ҩI�J�V�����J��9�Z���&�f0�|����e$sw�{�ru%Ey_T�t�̙3g���9����]���_/�c���S���4�I+��"�l25��+>��s����5��5�&RƤ�������]�:WS�)��c&���F.`qd��y+TY��򽮍|��1��7�B�mM>q��`����O̼*{���Ļ���ZΜ9s���
�a-g��Y���ӌ5J*$j"p�C#�>�!��f`Xm�
��i q�ZQ-����,��}U,�,˭�Z_����̙3gΜ9[�9�����e�%�������w��]���ʴ�̰\T�pf:�+ћ3�*�<���@�<��}�޾�&�Z�J��!�������Q��H$D�J�F��K��U_�������=m{J�����K����3gΜ9sv/5���9��[UpOI��M�$��������E�YD{fV܂w�牮�}��^Ѡ�\���%	~�j8Zw�Μ9s�̙�{�9��l߲z!��y���_�eW��I�g�$A�����,���+_)��: ��r:��H�z���D�~��K����U���6�u$io������q�XǍF��s��?�0�?�Gn��6[{
#���^A'������B���\h?�S��/Gb�0PYx�k��QkY�*���,�A�r�l�H�ֆ8L�f
'��y���<<�n%�ل�y���.#
K����yI���,�R���#t2�)Ɖ�=>G��e����������?��8Pp.���~������(�C��}�E��f<�}.�ʣ��1��vT
�(�(D+k"k�+�Gc��ҩ�N*�n��h69";	���Z�a���������Cݍ$��F�Cx��:�����,l[�<.)����5�D����)���mӵ-<dh?���::s�̙3g��a-g����]9y�ՁO	����0lC肞"���s{�����$�3�A��	6b\\��tI�����XE�$M��g��
<xV�^i���SG���Q�ŝdLȷ�@��
�o�����2x0(���ݑӯ*��N|!Fp"t)���d��Y%x�42�U�7@�!ޚqG7"<�"I��T$� � s��÷��	C��|���)�p��*���`��(BhA��3p7�D)W��������?3m� ��9S@8^�(�a4��f8����� M Z����*��<	��i���4�U���]���A8/!�R��d����oN�yj4vF� �	[�1Eu��>	ȅ���-F��f �,`lq3n�s�c�;�%q���� ^��X-���+�V/�:�̙3gΜ9[dk9ۧ��4�j�c�*�h�qSY���� )�{q��0@�Ʀ)".v1	i���3(��9r�a�{U�����A� `U.K�]RrU�n/nD!e�I0�#4՚�{�b��4Q�%�F#���aŉ�����]ml 	��#���} Zq������2LpỌ3��	���M��;��x����f���{O%Ƹ!7�g��>Q�1ދ煁��%�>fh� ���:G�&�A�ˠ����X;\Bj�Ы�e�9RL�0�%a�g9��Z8�L�2<C��yI��19Մ҆q�%��`  g�:$�R�pX��C��+K1�$J����B�+hD���(�Ej�(l�^.�![e�<h ��
*e�����N͘�ל�
(IM���T�$�;�VeIZ`Nih ؇~"�A��(��nR�����QR�g>�] l��>�p�}Bq��a�JŴ-��@�D�Ъ�[��PRgΜ9s�l���Z��9����Na����<c�����>���'�.��F�t*�#��u�z�ad�y�7R"8��o���L�}����o�� q5Bkn
|T�ks�<	�N"�׉,f*"���41��(��j/7��;�^�ـK�}���9�~η�qb���$��C,f��p� �Ka�KF��Ơ񄇔��6�Nu�?��1��,t*�� <Oz��{Vտ9֘��B��L�T��5G)J��,�"���@5�O�����0q�������l4�����DOz3����8���IV���A�L�Z0|��ς���x	'�)�L)�
��vx�pM*BS�`�`%��?k�0�6�ab����H07+rO{%�
x�1��a�p
?D��� |v�O��=^`@�����ŝDde���7yqV3[1�.�Й3gΜ91������312K��0����IL̃�B�H���r�KwBb�c�щ4Y��	��~�IB���әo�Z 3�+E'�h\y�[h2
^�I�t*@(m�用'�����Q
.�'z
0Xh���O��?�Hy�)��Y
 U��P2����&�a7E�E� ;�K8Z,I��؍N��������Q`o#��c�@6ii$��0[�h6��ވ0~�X�z0n;��fff�ZP"h���,6��(Ycg�^j�B��$wm�E�7��G�w����e�C����*�Eaxx�14�����C��Pv�i�Ի�����|�ӌ�0V�:/O r(���pi��<]�PLw+B-�#�������m�V���E��׳)|��9K�a>,*M+������V� ��E!^ �-pl����0� Rx����}�K���,&P�.��m����ǠY\�7�$���/<��ݴ�t{4ڲـ���i�.�Y@��ۃ����3R�Y̚���jgΜ9s���ck9۷��Q��N��朢}�C��{j�i��>�5�y�k^��W"#���o5��gZ��V£!~������?������.:�	@��(�������:��O;�K/��S^?����G?���>���y��e�|�|e8�U�s�`7��?��ON?������^�nc�4�֞�ԧ"��
~�S��ԣu֪U�<W��>��?�i�$�
q�l������===ͺ`�6mZ�~�W���vk��xWn��g?�Y�ρ��}����% V���Ҝ�ڂ���Snٲ嵯}퓟�d@ �`��ª�ٳ�<��_���O����q�����.������}���5q���4�KX�W�s�%4��� �zF�a����5�}ի^255�����mo�u ݧ%#R� ���A㱏}�������w�9�s�eW6�~l0��-��r�:��S/��C	�N �c:]N�;��#���_��b$���@[2�y3j�i�ʵ����u���ܰ�~k�&�U��~��zֳ����,��%�����f�`� ����1IZD�!c���o7�x��l�+(�l��G��~���7H2�YkO�X���O|╟��B�`�/��r8����b\�s��c�7����g��G��C�l�^������B$N�>�|h�1����?��~𪫮�yA�'�Q[Μ9s��Y��r�O�$-7i��Qy�4Q�9~j�/�[���7}��߽��+���y@h��"1�+\F+l�����I���+.�����O:�X���a����|kj��l��e/��ߟ$1��:���s�C�3��8�}9�����d }�<C��_�җ�]��	�P������}�����kb9��O��O�����_�v}��+����0�saa�c��>�������o�� �t���uiL(���}�c{�Ӟ&��B����?�y �0V/z�󡷘�%d���PCh��O~�-����? �`�m��CW�k�.�$�������/�������2�c��S����cox�?���/GM
QLP]o�y{ {�0���~D<���ka���0&$��-I°`��,���4B8m����~��?<�製��v�χQ�X�fP�YLUj��<���O����o�O`�k��{��J�<�u���~�O;�������l"����������`x���g�> h���~�����Sƈ,Ҹ�	`�fk����������c�AE����(M�����,���g��eVQ *Һ���g�ϯ|�+����?�kb��\��O����t���5P��c�:󪫾0�9>��=������o�@<�O��g�x�[������֧ҙ3gΜ9sV7����Ӧ1�*U�#?�O��<���DJi�5 �Ї^u�U���'�������y�;�Ca�xĺu���o5P' 1`#fr0�?�������I�(���9]333��[�|׻�=ٵk'Fj�z˖-_��W��?�s��#1t�*�r��U/9�����%(U�#N�޵�?�������.��bR�@Hs�/o<��M=�Q���w��y*�/��/��O�䮂/z�K^
~��_��]��d���F���|�)Oy��矇�@�W��U�����\xᅹA˪p�3��+��,	���:]���u�����u���~���tӦM�]z���'O<�H�W���p�c��<�a'�Z�n)��*�#)1F�K.9��YX5-��|��a��.�����p\容��;n���0A��)$�t�i����n���׽LH7��֭[�h����y�����}�K�:c�B�~\l�0��o|#�_�B���Ff�^}�ig^ ����κ�+T�tV"�W����߾}����l6Bβ����G>��'<�C��1RO�{�����������G>���j	��&7��v>������>���|PjL��5�z�[�������~04[I�1F�w�y_��g�gKO�P �5�\s��WOM�����k�õ������7��7�Η94�����>���A�̙3gΜ9[dk9�'l��ƞz��Z�*�΄o�饶1�x)`0���ϓru#�������z���e�h�"I����m�,�*H2�Mt��	�yS�����.}�^w�qGڸ7՚��9ݟ�"J%B{�]��k��oL7"��A�˟��駝s�����O8'�Y@Z��	<�9�`c��7�����}�nF=�5<o���g�_��?t����2��������w��7���O���ӟ������s���`�����D�.��Y/|����_����~�ww�Rg�����5�Zk������)��`f�����S�=2ͺ���,�F�uo���=��O;�<�������Y��^�������9�s�z�#����5�=�7z�o��?�\3��v�ՙ�I���/�~�_�ԧ�DX0�	���>��o|�����\���D=t[�%֭�'IG��6��	qX�Kǽ�0�<��aX
"]�-\��>��?��M�J k�XLg�̲�P��V���RYh[g~>�R�4N�|��o~�g�u��G$�Dp�,|+E�L����?�ɏN>�����'��~�6t�ơ@���%��Tm�i�Tj}�Ϳ��G>����������O��g	~��~����qN�r�=���;�m;�q�}�W����O>�"�-�q�o5�|=�Bi�S��΋����~��K>��7u����ʴ�/}�5��B���g�h��W}��c����V�w�����g<�N;�����<��GM�Ӎ �K�?�� /d��N{�W��#��T��7�����j�.���ڭuJ�0̻��k�������kg6���{�駝��w����8�j�s!_&RMr ��q�.gΜ9s��~kk9ۧ�l!���.0��q�/�~�d���,o����$)6!�,��2�$��#,C_����E/z���}��W�j���.�hx\kh�;�e�v�~�f�R�J��?���N��g?�u������BuuP���?��g���^�\q���}����_<	G�]����V��=|�K^�_��c�A!n�Vd���|Q��.�+�F��͛��pNq1s�y(q�O^z뭿{�߿n˖-RRY����H{pӦM���������+^�7���������j�p�_��s?x�X�C����7]7rƙg�_��R�.�ֆ�>�h�rss��ٖT^��y����g>�뮃�iD!xٹ�9�l�9<R��r�X�@z�'�v�M�P���,U�95|��;�v�c=�W����?_��<�_�lzj���qE�I��̼�5�Y�zn���y�Z�^�-�u�>��+�z�&�/���m�z�|�#I�"��?�я�y睯x��?�	O"A�3�`��;SSS�/|�o�u��G?H�yAҗYV(&��'R�
��y���?�
f=f�X��+8�#��^���u�Q��c�ic%���=�C���7��3����.z��^���[�������������?����f1�>��0���o�?�a���Y���$0�}=����я~t±ǹ�AgΜ9s�l�9��l���E�ҳ)����];$�=�EI�-���O�g���
�:�1A x|r�-jes�)�ڱA|$��u����uo|�3_��+���8����6�R4�H��vKg~ב�#����׍>��#7��~�֛n���i��dh "���a���u������:��n�~��Y�~��-����QxPǨ��]�L�>��}�����;�iWi��)N"��yKOu���~�c? ��7�v+h�\w{1�"X����y��g?�F�l!
"�b��/�~�=}����e���w��(�3��K/�\Sp�n�`j���TK~��c�-,������P��˨ـ� �gM?��g����3�K.��JN*���:�iR��/��RQ�I{�{_&WU���>{���z�221�GD� �4�@T��@d�`�Q����A!!b@@���^�1���E��:��Z{Ww*ݝ6��}Q��動�S��T��������R9V�l��DR��^#'L��&-_���Ƅ��6~pB��Un����)��g�]|$��C���o9���g~���ｧcJ	#C�̨Z� ъ�ܧf�+�W�m}F��#ږr����TK�%�W7ݼp����7�,�&�6�
��ÿ8	��{4'�P9�V���/�A�{��ߥ�
H�aA��T���	Sp��d�k��|�-S%�r�zWW�C����z
_���������W�`�a��=�d����wР��?��*���s�������G*�	���/��F�t��6*w�8~��_�����:���;���c�8.��T����r�ҟ-�c�=ꐬgw�l�
(P��*�A��	��U�#���{<`ڱh��fH�8Z��|��{�[������i�q<�[�R�t�1�\1���.���I kr~�q��)W�S
IVG+<�qת�I"ؒ�vLr��XX%ĪU��x󿧌�m��I�u#��{��ԧ>e�	v�E�"�Q�V���)�����P��KƱm�d����J�袋x��8`�ͷ ��:\E��۹G���+0�-���*�<�'kYj}�M7�9���0�r��e�`���=�)UyfÍ7�����Gmm���7�xc�ʕ����?��>�HtH�p�رc���s�=9��&���>���Rg�>}���N:Ic�a�i��5��F��F1��o�k���F�v�9W�����/���k=���ʒ��TV������+E��;2�#0�g�y���s���r�n�p�`` �HA @N�'F�[���3t���|�Q�����a����P�����M�t�M�z����M���(�T��/���e�7�-����(�Fm�z�j�H�{��F�1�l��Ԅ��Զ�z��s���l�˱�������9BPᗰ�BDp���o��˗Ͼ�BW`�����@�
�(�V�����rE��]�m�,�4pC��»<�/�&�<*0�z����|�(�	
Z輦!���g�_�ꕗ]
�-�╽�g:gT	N83�j^�a�W�j[������Lbr�b4�7e_�,}���>!;�9�2�&�?w���>��Nۗ�ʌ�$��1w�r��g�]G�FL�x�G���t$炜0��d�LNa��y�qs�e��4��x>S�uC����{b�;���!���T~H�"��L�k�:j䈧�z
�k"a�B�)�C\n2]7^^�ׁM
�}l���	��ݟ�;`�?<�$.a_?����jh|
�1FK{�6����'�Hi)�e(Pג�jҵ�k�7Z�@b3 �k�<�P������a�B�K~������7J52	��@o�m�4��3R*�2O%�@W��J�Λs��O��uןw�U��U����=t����q�BQ�ǙS���������@d^|}�������g��'2�O=����oio�uK����M��ߛ��s���ۖM��S�,����$��;���O=!��m����A����Y�$>���.C/��L(K:�O?����vo���bO/<��S*'4#�ki�Cwr��W���{�l9�K�*(S�kiT�K(.�H��p�}�t�er��`�ѓ2��_$tF���m?�Я��j5�Łbg)����f�
(���kؠ�C^���l��r����S;�&�Og��3�q��z�ο|�kk�\.[���I����s���UN�N��hѢn�����S�Ky�7��ˬ�4�1����&�s�z�hLK	��Q^�\�ֱ�F������]�($9���B�(��ۦXQD��r��8E"�s�nuZ�3f��Y&�T��������symcƌy�w��\�@�y��z��tȐ!vq���g�-Q[[����/|�'�gϾ���Z����<��ȑ#O=��[o���$I[9HIZ��t���_�k�=�޹��ObUg��rw�]��'x[*-�9�̳���l?>0U`���7���</����=u͝a�Z|׍7�x���?�AiE-ݘӦ�t٭˱��bbu-x0t�P�����.<������A�D��-&��2 Z���y���+�C�BiWI*��^�D�F�]�{��'ѐ��<��R	���ٮY����G�^�Nf��с�a�k3_�<�����Oz��7wc��ʸ��N�]�d�?����λ����8i��w�ɥ�μ���'O��h����
WV*b�^}��������B�*P�@�
�U`G��#���J�Zے<%>�0���Z�z*���t���/��?��t�7���M7�����n�l��X��D��E��[S�D���Gk�w���-���[��zz��Z��h�5A��.Z�mja#��6ވb�a	B�:Jk�=�e�p�i�W��
�I4���~�m[y��kolٶ��y���ŤiS�=�Dl�$�����رc�O���|����&u�,IkǄ�Y��(3Y�	����`���Q�Q������j�=v�ᓙ���y*l�E_z�����V[mD%�e��q*u�q�V����2�K��t�V��?�n�����B�~��/^��k��f��-oD~���
T� ��2i�K���8���]nQ����/�{U�T��@8��ʉ�w�7_z���ߺ��3fTʛ�&
���Q* ?�D5�M4��������<�&#�;����wn>�S3���p����CX��欺�=��'�\��$V*Gv�<8p;n?�7>��[���I��è̌�N�1����ɫ���縃>���ri9*f/�y��wL!���V���W�2�	|�ĩ��<��jo/��C�K������{��BA�N�o)q.�������<��&�˳�P��2�/c����
S��h���݋���g���4!�P�4��Y��3���Ϳ=�j���$Ak�9����"5�7���zr��(P�@�
�U`ÆT*�@��p���ʥ�&�1	��4���a�V�X�zS��(,�Q�ܩ^I��>z��I��3g�6;��H7�Z\����a1\�!�P�֪/��R�T�T*� <��g����ۇ����;����ֶ�j��n�uv֖/_>r��N1����j�Z�\�3�#���EZ�O���Y�ivӊJ�7Hd�g��Z��]��]�J�ʏ9�e�-[�d���ÁJ�p�c�v���0���vuu}��ڹ�[�AB���#l�)�m��f�+��\��*����FG��"�\�,�'���m'���n�m'�t'W@��	&Æ��w��y`-$˔/�0i��� �V�q⤓�\��ȑ#>�૯�z�wt���U2��s�	5O|��5�~�m\*�����X�]v��$�{K�%�))�4E	��W�V]=�5c����ZR	��!��Y��8*���k�Z��y�0a���X�l٘��J3p��C����Gy䣏�i�8���f��I�y�n�]�a�����{�1cƔJ@�	l4\���ĉ��+�Yh>�jøa=�����(P�@����od�ػV�p�O5��0�FK�Ʃs�f��Bl��s�%[KBa�&α �Ѫ��EԠkv��'<���=�l����W��������Q�UI=�Yp��_�e�/^{n�F#G�P{�ͷ�z�����M6A���xGVX��$:l�D��{qםw*�����Gs�9�͹����<y2�,W�Q�E+�^���Y���3�5���HY�Xp�qvƅ���Hcy�f*���,O�t|�M�tĥs���˿x�a;�5=}Oj��<��^��9sY����)�3[Sc-뉴�}�1E��`�9��M<z�/���3��)B���}��7�<��[[�@7`��%�y`�s��r�{�i���o���(N	�B`f�_�OK�;�ڔ�������^���)qAYFL�ċ?��3���\�"0��5G���sN�uW_��g�����4��" c(@��,��Xt
^�Tz�ҭ��P˵��n?L˟���S��:X�Z@�ࢎ㏻�+�\r��;ns�Q�Z�
48�V����8�g:Rt�cE�K�T
e%e��-a��-��F䙺���J]��p҅�_w�s��xԈ�eY����UE�7�z�왗����3�b:ɥ�!f2O������1LM)��+h����jlP�@p���Ȣ{�f� �2
���lZ&�۝w��k��B7�1���,+��
(P��?5
�U`��-�Ʉ��q���ݒ�Fpd\3g�|衇Ə?hРj�V)��).k�N#�a��q��Ps���[o���q��~�c�^/�eW�?���n�ɸq�]����;��C�}�]x�c����LF��b�w�ǫW�>ꨣ`�݆aLoѢE�rȴ��t�M�?��\�����N��v��W�F��f��rc+a��yX���迎DKE�0�60f[����Dp:~ ���o>����{��&����eI�`��%�͞=����������ہ7!S��m��
4Kq��I����e�| 8�%\CZ���N�8�s��#�h�RX}��%K�6=���Jݛ�#7 �ʺ�W��l�0R�'�/�CR��_|���+�t�f�m&34��.ZV�s)��r+`\����rT��5d뭧O�~�uױ��i����<�/wwr��\�:�w��;������/ۤU�,=�S�q�c�=܃�"@�ۖ��|��r:�=��Y�6H�	H���J�ʤ��W!�xKK� _�|�ҥ���gF�}���r�ρ���&1�fͺ�[`��ba�TBY��Z�<р1�l�W��U���[��~<���)����w���ͳg.[�r����k�Q��v�P�[�p�СC���[F]S6JȚ�

(P��?;
�U`�F=W���֊/xQv��B�"��C�a���Ξ}���,�aȥ��cY�C n t6�
�e�T�z@�P��fJ�ʴv�W���w.A����ZV4�Ǟ����=�m���8������t�a�<u�9zo0��/�r؈�o���x�i���uB� ~�1�~�h�AMx��'�*m��H�B�G���~k�Ɩ�T��N��S�����J!3Ld���_�'�^�3�Ж(
��0l�DM�����oW��s���oX�v��nX�,�$��̞u������F�Z���8(#��|������SO�ʭ߽���.���90�,EJ0{�7�1\�Dfq��z��k]��c�!�����mXp�s��XK���Ѷ�z~P�V�GK���vL?�DK��T	θ`y%j���˸Q��q�+`D�Lx����\�ܴ"2K��a%�V��ʗ~zׂ��}+�z�#lE��;���+�)Xk)ݵD�Xfz��F�3dp���`��%W9�%$H��>r�������g�}�A���5��A"Gο�R�CΣ1�s�yi�xŵ4�y$�!�Y'�3��̲$��:�0?$�����?������������:�-Iռ+�9r��W�g������c8$a�絠D������ǎ{ϒ�l��/�ZJ��D���;�����2%\���u��;�(��,-��6�vC2G�z�
(P���Z6h�>r ��Sʏ�t�4O��$K|k)�?7�N;���"�u���셣6`+�0���T�@Ȟ[;�n�������<��믟1cF�Z-�e
a��/]���sϽ��� �f����{��P� ˊ��B��W����#�����o�����6�[�7��|�������tС�#<6x�9g_y�5q�T&�����s5K�o�=[��2N��}��z��*��'���41bD��_�5���_���!������xI&3��xk �@>���Z�V���j�R�O�]Ady�ݧ�{뭷��ʋ�E)�az����'�S1�=�cŊ�h�v�U�5�[��X&��J�����κX��r�I��i��}8���)��7>fǱ{�d.�-���$�}X
X��R�͝;���Nw�\0�J�R=⡓���=#7��MC�B������{�-��vo��f@g�1̓`ԨQI�>�����g��q5��_|�\pA���$5�+h��&`�=8O����|���N��˔с��z *cƌ���<���o��� @�v�n����]@��-*�����,&��019�z{
F&��l��vo��椣��կ~�c& �e�.�?���Z38�D�G}�>8��#aJ@�I�
(P�?\���CT�?��.���O>��_�4-�`#:
���:���e*�w^ւ�Z�k���2l�D��	����͹����j���m"+��oS�=z��S�$�u�6v"�yW^>���8P8d80���A0��@��:�4&�}�f����g��\0�\�8��G��>|��ѣ�]U�:�LD�9��~�������O�2y�IڐLc4oR�Q%��
{gRo �?��K̴J��F�|�<t�T`ޜ+���a�'��qEh5"�P�T*��@`PRf�vҩ�N��d�Z��+��o�<�~�?����j���繖6�O�ngi��}�^q��	��5
Ɉ卮©���S���Ѱ�:�w��`�߉3N>��:�q�5l#H~��I,�R̭��+�G~{��+/S/����	̦cYz��]1�:�o�2�D��%��N�8�)�D])W���r���nM?��'���!+��h�f�V�3��B������n���;f͚EC���:�%��|�]w�����B� �	T�mC��ʇ#���q�I'�
ʤ.��.	���ݜ��K��}��,��S�KC�R�Z�^n���������e6§���\ea�::���F�����U���m��R�L˕�e�R��_�˻�#�a�g����>I����CKY�˥~Ȉ���F}���&�v�݁�е
(P�@�\�������!hWT�3�g��عI{6�D�&N$z^[��8s�m2'�1��+;b5���s�	aph����(�e`SRCH��A���n&
Y[�@�@h�k�I-���z�iӦ-^�xֿ|=��F��͎�P��vP�3[�ݍ���s��6)�Z���-c��}m#fbl����0��^��si����>h)�m��#��4���rl+� ���G��b�^�&N�u��+�
��u�+��p���V�uz�~��K��\�2ÞnZh��v�o�u\=����= 8娜��}R��p4��X�Fe�!�u���fh�a��l�S��҉��7�Pײ��5���Y/I4��3Qd�,
�-�݃B�ț;��<�q�<l���3g��
�^�	���U��љ��I9�`Òz�/���<[��{~�� J�YXC�u\ƾ۠�"<�m��}�R-�8l�l��	$�\��IՕrYY��p��A��D�4u��L1�e]�4���Je�RmU5X�$C����1��^siOZqF�ѕ�,[�l�c���]�rP� �>��d�
(�ρ�kؠA3	a;��� �P"��k�J�"x�b.�?���r�lC�(����(ϱ��%P!E!��9Z�{@�j]�A���X<�{2˅ϱ�z��H|G68 ��%H��h2mC|
#��L(q{z�U��nǫ��a֬Y�UҲ�����!��b�`�0¸�p��m�?F ���(@�8����ڱi\MQ	�7���<C�aq�S�~}�$���1ʑ�i�m-"�~	� ���-0vg�j���A(�U:�1�N� v��@��H�d����
�L�]��9s�5~����'�9uv���t�Y�r�Gk�Y�6���P��r�6W�>���)�w���(�g����$�&��@�H�^�RQ�C�׈�s��<E/GT�<�2K�*�/*E�j&�M�m���V���D�"f���рњ0��3��+��ʹםu�9�#�I����U-MemgR ����*�Jp�l�0\!�J��Sm���H�]Ig��|�w\ +���º�4��X0��1X�e�5��ȇ9�3U󨟫'M�*�J,.m����5����'x�Y�aD��ˏj1�1�k�tB�����<�=!�^9o��CG�g5�U��Lg��6�S��)��*�
(P��?
�U`Æm %s�
R���1��}��mX�q��1�Oj`цQ������2b�t<�ֶ���>q��pq���l�cB�,M��P�'dy�� ε��G&Q3�@��F�H88������ �������?�3�ZQKq����LO�S%"cSc����YhIP{ �3$,�y��F����5ϔ(	$w����V���r T ���:�a��yF�M��)�w�`�P<���^���և�(�Z%%�<W��9S8$�5jk��;, �	����Go�����y�J�8e\?+��٥��O8G��*-~�ı��;*-�Dq0(��$aȞ�8�[�I;�� o�m}����8��y�֏��Y�0r����,�%������	�F��k���y�����n�8q⌙g�r9��rXv�t��J���2
�P,�C�.<e�Z73��tb���2�G]7��#��>%���ϹV��9�5]�V�n؃���4�#a�m;cT�|,��J�"���jZs���E%��d�6�'\������{�=���pfZ��L���=�!���"�
(P��*�A�`M�#CQA�f+��B:�购Sb`< 8
�D�8��c��'b�*<�FB��P?��B
1+Q��8�j��]��SB{xf�� �U��t���!
�	�>p)�Z�_�)�:f�54�g�n2�t,��%f��=	Pi��]������̅k!������.o�
������P�F�/�d<�u���Z��:�/�p��ؙX
c���|�j�"��-P���{8KL��:"l�[QZ�8�SN=���" �@��u��pk�? �C<�-%>_Ci4��*%�Z�ex cv�;p@X �Y�u8 !��r�>���k�[��/���5��l@y�3C�����!���1��`�׶�WcL��Z�ۭ���$UFY	����ύ��o�1�vT���}�'�:�1��_�9�v+�y�������A_�ʡp���dB�k�(�A��9	���(L��7�_|����ZdV*�b����V\�Vq^%���Eþ����P�T#f�v���/�,�̡�wʒp�
(P�@�*����ԵQ"�zH�3@Fz� 5�bo~���zi���ʇH�'|���t�Z�0z�WOXڍ���X#5X�g�GA�W���"��M����4�H�;�^z=&k�FϾ���g�{ͥǲ����/-Y��Ycqw�V�`��@����U���44�9)�t���7d�{7�����Q�X
(P�@_\����Fr}�JO������H�>���|����F�^Q��}=��}K����4ϫ[�an�Ύ�]���מH/BȚU��wT����6s�O�h��ԗ�Z�^�j��u����k�������a��e͑�Y�Op�־r�c�{o�[=G��W��A�n��Z���A�d����ҝPI
(P�@��(�V��3�
p{1+k��Ⱦ����7�����>.f5=�E�}���R?����w��/{陵�X��{�;������g��|��K��\�����Π� k���2��70��\��]���{�En�����a�U�����5s������c�k<Yõ�G��'kݏ�](P�@�
\���VTz	/�t���s{��\��l��n��i0�W���}����x�|�{��L�/��.5�\�^kz�{�J׬�K�t�i��t�(�O�����Э��㞦/��}�u���޺.����A�ٽ�x~/Z�|Zz�Ԣ�O��ٹ�3I�
(P��*��^z�'Ni[����x}~�o�V&0͡���_��B_A�祁y��p$렸�ר>�뻿�:*����`��t����+�o)Z3����{���y(P�@�8
�U�=���|M��h�D�qD�О����׵�&�p}@]���Kq4}��z?��� �5��Kg��r��ԗ��0\�O��4���/o��F�\������=�,��b]I���͢�gF�)��!)P�@����� P�~� N    IEND�B`�PK
     �8�Z�GR�8  �8  /   images/08988072-c7a8-475c-9331-8aa77c72a02a.png�PNG

   IHDR   d   W   }nw    	pHYs  t  t�fx   �eXIfII*    	      R	               (              2    z       �       �   i�    �       2020:08:13 11:56:58 t     t       �    0221�      �    0100�       �    R	  �          X7  7bIDATx��i�l�y&v���ګ���������%)��fƴdy��M����'�#�d3�`��N��q<c)�eG"ER\,����w�}���N���<_5-K��2��@�ѷ����=��>��|�!�e��������I�|���<ϣi�2,��:$���ť���_����bY�w���}���W�9�K���E۴�������{�G��$��0�-��i��qDӌ$I�=��dI��kf�N'K3�e�Ca�[��μigV�����K���'�/��	��عB.��(�x���G�w߻�~���-+B�a�$}��c���^P,����/���|���}ٶ܉Z��iMNLMOM��V����V���VE�0�8̒��ϵZ����}d�>����ph��h�l'_, FX����Sd�S�7���~i4��0t���t�0���q�`	���W�zg�����(2��)Jok�������`��`ɲ�ﺮ��:��Vd���r�z�J�� �|Q�� òY�"]ϩ�F�hEQ��,��K%�s�X�o����!�I4��Ngfv��pA7�*�J��Y)�,�{���[��s4��,���P��b)���wF�*W�e)h�I����c��aD�x�T�ɪ2Y���������A���Ƒ��$�p~rN�9-5��Ǚ����7N��i���QO3�(K�Tq�F#�S��������;E'C+U)�c`ȐD,��᥈�hڧR��5Q���[�ɕB�z#PΌ�7��g���?� +����~���HDe�/>���Gg�֙�G� �I� ։�8�ș	^q�;.*T�tf����&i&K��W��u��l͍=�P� i9~ pQ�M%�����L��~ gY'���)� 
%I���[��w��]��a���_zAd�Ʒ�"<iSY����s�gWg���'1�@%����2��J � %�E� 0t��H"�2��q�QF��'�JrQ�ɱ���s_��+ł^�( �P=߁J`8fDo9�\�o5���G~x��P�r�b�<l"������%�U�,?MC���)�C�2�7�8�2��N�	/'`h�"���C>BS%Y�&�u���0���	z�޻�����y�J���j�Q����{��Jn1g��ngc[ՌQi�$��8Ψ(9��:;�>�'���t���ƑEs4/�� (��&�B1�?��Yz>Kj�p��B�2�\W2��	C��t���Y�d����y��We^���o��?wu�2����v/��Ȏ����������N��|����ϝg�e3�A�Q��!�!T]�5Y� �*τ1r�&@��	�HLJ��ѬZc7�J���.0tc������|�{aJY�᷾i��;��蟬.��տS����î�9-߿��_M֊�Ԋ�!�c���8C�{f`���U�I6͢�G�Y��8���Ȥ��'��'�8=Q��b�K��9�8��r�za�-~p��?l�T�Y�s�i���N�(�|L4r�������F�K�2g�ƳLC�D���s����WMUP���h��Y�y�F� ='�R���8�\3����r�*��}M���S�֮M��5�ze�7�n���,Neϛc��������W��TY��8~��o�'M� �)oH�pfm<K�<�:N�U.2���M�bM��4!�YuM,�d�#��!1j}� *"����p~�_-�����?��_�.�]�f�9Q�9L���0���hY�r��i�zJ+y!�JK����`}Ñemi�|���Ϫ�gv���-��
#{���]\�����G�L�e'$1�}�K)M�j�u?�˭��:w)���t��+2{���I�ēf9
Fdum��v�=0d%-���c�H0I-�RB�iF�Ad�RQ���:a�<�<�6�XD��*C0���t�t� �#?�4�L�B.Nѩf��^��)��e�2Y��ؖ+���4W��~Y�O��U�x��oMۍ��DA�-GEa@ѥh�!G'4�Nå��k+ޫo��Zo4�ի�gYc����b��,���Q��09��LC�OB�S)TEړ�Z���5y�Cc՚�
3��ҝ{��5A�1ۇ��</x��R��p������X��)������p;9�֌ݳ2���E��6��o;C�̤)��������=s���/���?A�n�춨s���;�LǻQP��z�?���(W��ݜ%�f��Q��#N�Ó,���`�F'�5���������S��89;����,��O6��㔕鴐Es�h捎!�']���u{���e]I��(Is���7W�h��Ԋ����9����G�Z��}ߵi^���3�Ϻ����_.,���Ȥ��(#dd���,����?Lҋq<-����:>�,Ñ5dN�t۶�0�X.�#�0П�9������1��
,��%�Bfn���|���+K�9�{��Ӷol���b��s���d�:̓�dI3�(	��]�b`����,l���Ku*��Ӓ^G�1F��R�4GI�@e~�Cs��!�R�����I���X^^yp�n��+��G�<�l�{����*��W.U��(�%�aDfc�p��Ж�֕���Ԥ�`����0|�hl(S����m��ciqᆬ-�X�_�aL�lD3��������h������%����{cHH�e�ë��N�䝘2|o�q LӤ�3,8 A���?XT�XaX�0r������zMv��K�(z([�
G+�α,'���,钐W����T�8��[#ۑҌ��tC�-�l����E�]�.0�Z.4{�9*;�E�	p�"�a�HC�y��Kl�i��R(�������7޼kG� �Xi,� H=:�y睯}�k���ի�juuu�����(j�,󂠍�a?/X�{����n׵��'�����=��ù�y�����V�	{�F�(9���29*�_�^�@�fY�5ç�@�Pt����`(�y")��I���@A常�	S��HWyF�Ћ|��s\�Az͠��~�����k�-̌zC�1\��K�O���pH����wv��$�4�X(Vk�l`�V ���W�����Xdn&�fgf%Q.�ʕjMU5�T�1Ib�0y������2	Fa����k�j�9:��8�CQt|����{��+=	e��[��{�)N��[�nwt���?d�Q��4���x�k4� I����BGMH�0u�^{�I��I�����~�V{��gm�m5��i`!��~�k��K�!�W�碋D͝*��H �V#�������4�Ty9�(I���]_��n_f�_��1 e�����J̰���|j,1�1R���;��n�x�q�7l�� R��A!'���rx���U�Zy��oC���_�VΟ;?91�q��q�GK�(~À�5C�zF�G� `Y��Sǣ��}���
�mby��)�>��'Չ�ÿ����R�OȤ��&�� U
R��8����~o���(AoL�8�v�4*�/�	�ғ��[�;��}�N����C* ΧTq����y��t�0�TRz�\�E���Ȳfo���4��v�!<����---�z��{n8�D��$Y�1�ƙf�踁�e����[�n:�[�T�S5���+o����Isbbb80����j��<8:���F�dU^���-���ZI(US&P�8YrOlˉ)��2Cy���l�3��X��v�{e�]=���u����P
LeP���۷��k	�+*�*�S$rz�)u&���Z�p�jVB��+s1��|J���t%>�1�؏^{�UN�ȹ� �ڝ�^�9A�񁲾��EɥK��Y����Z�ɺ(J �����b����;w�X,˒8;3�jZ.��%:��eE�Q��gC��>�dFL�斖����!�f�AV0Eɸ���(W��?n�#w� ˦h�M�N;��JR��q��׎F6;3)��/M�D����
������-s l\��P���L��f���
F�>�
��AP�V�� A��*D�RA�i�:��>yBj3w�ʵOI�8N�)���p��������'tF1KG��F������UӸ03��~q�9><��qb�Q~t�_������L$)��F	%��T=luP�l����X�NTG�
(
<M��f���儑%�P.�U�C��%�ˎ�2!K���0�ꘌ���?�y^�P����硁v��tM[Z\�q(>��f/�P�o��o:�=pF�����9ʪ�"゠7M7x 	�(+f�Ӳ�zI{��fWs���lݼv;��G'\��{TD�j9�lK���_>��..TeJ�|A,����J��d�=�O|�'G�RiN�Xi��g,:38�X`M;N����^Vڣ)��L]0V���V�@�xn>�R�$@DXA�J����nw�8^�-.��1S��޻�����eY� ���z 9�������d�$'��ŕեZ̀B&2t����������i�[���n$��!v�$#OT�0B� \�{vfx�R�g&�~����Rm}gW+���C3Hv�����a�'������{]���e9M�r1��iV
�8��0X��(��ן �#��qm����;88(���������\�]���b�4:�8h��BR|"X�.E@e׮^��Pv��Z���\�x��j/���Lς�|߃U�9N��ر����,�u�%�ȗ���K��:l0I��I������b����%��
ͣ�ߦ���TM�"�ݼ���g��!;.���y����������g���{��|q��h���c��T��CNբ�H�8��o����B���J�5
�vٖ],_y�eQR��|�ݾp����"~���j��w����Ms���8^(K��.//C%T*僽���F��b����&&��.d��bL�z#m�4ke�
��Ί�Vr<��Rf��/O�E�Y&2Gr./��qpD3#A揺2�(�+�I��D��{;�����������8�����K�	������>��޶nD��:'K�v�8���Hf?�@�����K/yP��O�N���n�R�lmm����_z�%���t��}6g�:�'��Y��q�ɩ���J�12;;�3B��kr���A��\i�l�4u�-�a���s<|���{a�KPq	D̀+�%�s� D��Rtx�L_������ �-5��b�tҔV�'%T"(2�0�P!4��}��^��Q1N���=FVJ���Ri9��OՄ�����[�Ls �W�Ȓ��\=���*BƉs����� ��q�>g�Ï��i�����6�P8v�wA�(� Ѳ,2GfS��K�<�1z��|�5������:�9������<]�+Mk
+�mwo�S� K>'��)�����s��QԨ����)?�u-�}��:�Ux6�������[H����R%�����-8Q��6r�,��y�3�%�ea��`a&>W��j�40GPKd�J����D� �8A{�4�-������o6�Љ�R��?��d|?��������hنs�C�r���Z�����#��l)�f����	/2Ղ�x�GN��� (ϒQ̐Y����|?u�$�%�,Ӄ������vx\U6�"mU�R��7wUTZ�O s!�6��e��J�3����@�i(?0f�ɲ��Ίv�����>�܄������C�A��u��Z��2KL�DVH J�UD��<�b�T�N�� Ppw(���脙���i��� <�����b����D9��ZQ�jB������j��g"�����₏��YVU���<��eWSzFӾX-1m�r��u���G뛾9��WI�[����G�#��2hmn$�ջ7���n(��~����ڦ"�\�&�V�a���)�KqD"�����LϠ(��\�x��h`�Xh5�/���+W��4<=���!���$Y�V��Nguu'���������D�A �g��������Dq��'�B���t�v#�kzk��9L(h�A��Ey��K�My`��ƾ����N���p����r�*�hw�a���ۅ���I�Ѥ�D��)T^���|⸨"�������SQ0�S����x����Y�u��D[�rpx �utt433���_|�y$b�����4XKK�иS�:����濅]__�i�ڋK�1��]��|��:�5�u,;�K^���\���|��55'�P�3Ϲu���&�	�ʞIH��i���v|�Ix���;茡���hii|�~�)IF��:s<�Ő�%�FV���	& !��f��9=ܧ�k�͛7;�.t"�[�%%��-���6�
��˯�lYΗ��b��ש(�O�A>,��u��w�}�6Q4p�=���������qF�����R��Xge�j9 �w��Vwh�ЗG�-0BV��~(��<���&���]g|�l5Ǹ�^��9��j��yÛ>p�����,I2�T��XBF'Q��#Sh>ABӠ0�;�f�w|{�XM�D�յ��W����$��ۭ�	���^����=q�kde*�`�G�}6X����<�e�jww�j[V�Z-�������c����ӄ�����x��K��@,�$�p�	EG)���h��\@�);7����}�$�m>�P�$�&�̰r*�G��"�o@)OŞ��X��t�Ȉ+/�X*h�B�4=jv�8h4PU��4���>˳��n�F��$U��޽������&�P7n���~dT��`mmo96D9tp�0��͈������-hThq2�Wp���z���{R+5���ٍ�zN$#�ڵfs��g9&ʓ!J���vh�4-�T��O%,��/H"�<�I�2dE=^�D��cW�`�,���6��A�h�㹱�Ů��0����e��,�-,���n��� R���ު���Eq]ك����>bv��`e�n��EI�\fXr�b,qML�F�M`�R�p0"Krhr����:;S��m�F�}�6��FZFS�R�yUJ4%"O���ЙK�@Z!��(s�յ$�X>�� �8.bXp=�Z��<;��ŧ[o���!Rt��cJ�%~yn�IYY��d���V�)b��$���C5Yp�y �`؋�"�qqq�eXs8�e��E�>�O���`��33�����0)�V�(��*Xlj	e��Դ|>l2`tn-���`X(H2�p
���+3*��hɠ7::����ܽS�v���`�0a�t�7J�2�8d�����T�R6K�(�x�V4�2�u҉%}���7��[�߿o��R��ÿ�5,�#ә�i:�������T:x���\��pjR�لF���_X�CY�lh4.�8G��NÇ�뇇�������R�0 (�r�ΐ��k��J���⡹��
�t�x�D�ʏ�}�ov���g:�%]���|G���D�[ ���9��Q�@J)G�TJ�=�Y�:�K�aFƤ�կ��|N}W�i3/�-�7�ol2Gy������RA���R݁�q+�/~�&0D&�Ab����$j:^���8"��i6��?YaH����"��Ο������?�C�ݹs�����^oqq	>����#���8��,7Q2���,;��Y����]Z.RY덷E*��lES�4� ��$8��H�X^$;���K3.'inDc�a`TH���������rH�
���ݠw;���5?N�������|N�kt�zvnV���v�]�D�iT�_��_��:���y|���>���6����ޕkW}��Z�e�~��b�t� tɵk���(%;ۛ;���cK�_x�tr�E�'�yJ�P����<?�}�q-���aDf�S>��S0
M�_�%�̶��֎!	L��Xqƀn�B)�h�#�R�][_\Je6�V��;�����^�6C)a0�󒒄*��pt�S�J����ֈ|��7K������~���Šsp���
�J��(Y�_��|������է�4]?�L��ܚ�@�Xr��|�Bp�7����Y����x��"�$!��N�zM^h�:��	g�L�� �,b��i��F��Q��x:��B@� �O>�$$(+I@a�>I#Ab��ls+uFTAM�m�����Q�v2�/�j�Ō(�A���L�����\��|��]ZCN�� Z��r�샌lk�*�J
����~D�����J��v��)���Rd_?����۠����1��l����DR�3x�,Hp��p���pT~i9�ۧ�!�eQ�*SK*Q�T+q�H��`����o�^{���D��ɪ	�%��t�>�!�qyau%J3S��_�,�?�=���ja觺is*"�RP� ʊyUbN����җ G!�+�t�E�f;��v������]�x�TN?�קL��YB������C.����~�w~g<ҚA��`��34��D���gg��sj��I�@��h
�?�R�Ɠ����4[]��x`��4l����/(���UtCp��]
����L2l��/<s�k�쎩����9Vo�6�h )����iu'+լ�1����5j<�y��{#ۮ����vg0��E2���v���C�v�����l�6���\`u:�o�e#�k��о������ګ��I��O]�p�oFzrq"**h�F�����͈���O��ߝ���_(��ɟt�|����4& Mm	)���"�d?*ϐ��芼&�<d J@���P�NV�N[�Y�.��dc�h������:jLժ���x�%+��,�"� �ث�����#��?;;��g�A?���2����d��`)���/~v��������N��ŋ��?�T性���xN��ɂ�i�b�T૾G�l{�W*�|9W�vw�{�s�B�Y&d��x�͜� :%���.
"&��T�@��4'�OC�Kd�sp�7	�*�h�\/j�	'�����7����p�P`p3�^��s�NT{0i
F�N����ַ@%�,�6�f~����\:�"Ӆ���a�X0tɈ�p�����`���l��7Y3��'E^���vr6�t�pa-�،{�o�ߵ��oP�է�4쯻��q���^�"����6-�̩RT���0�]�%ΐRjU�$�A��@2���+��9��o�]Ȅ��5�.Jӗ����e"��I(uR@V�V>�}o4� �O�h� ��W�:�@
2�?��>�J��TŁ� �Q8���rE���J�,`)2�\��Y�=Y�L(�v��λ�(�dQ_Y�)n���q'<,���<^N��CDm�1��+^���$����N_�8���H
z�d"'t{����ũŉQ�'U�qʊA��3:�3��L�+�<9i�����Ȏ-*
<��i��S������,���Ȯ�d-ͧ�:��Dfhw����Eb���d.�U�g�Q�5����{NN3��كi��j�j��#i��.3��5��NS�%S``�A��aT����G0^GXL��Q�g,-�Yx	o��hz�Vy>Y��8'}K+����>_(K�F���%�K�݆�F7�3_ʫ��7�{c�B(����鰐���8&�V�y��{�&�u���1ޢ�\�`��s��J�o��*i�D�Ƥ�r^���%�3��T[P���5XF:u���4�:::Lrya��-�#��Y||�Dk�{���d?v���u�=~E�EJU�rI=j �4�y��,��p�a��R���(@�/-� �фB!/J�v���K ���<�fqi-��Hۜ���M���3{�tp���M$|��X^^YY]���Б�.��EE$�JN��rc�@G�m+�LUXQ�G~�N��aY)Cw�$�B*eA#' �SlF��d�RCzA|"��r�(�e�-V�b�]
z}H7�\Qq�Pg��D����˕Т�:���޹�m;�bw�h��./.,��NNN���i�[7a`��
E��x��A�|i�l4n}�a�q����˗/�d��~���wn?��k+���dJ?1]2������NG5)F�z=��
D^6
��V)�E�e��,����h�8"����I�h�ۜ� ��/,�Ί<�ZB��M���4�7i�F����iU/�ϰ
�iE�txR�>�O=�����zxtT�V���-۾q��� ҁXŏ/��D�r����W@�@
�u��m�7����-
��#�E�k��藂�f��\m����`�a���w�*NV��#�C�Q ���cH\pQd9G֙�32�G&MTX�����)a���|?��~��E�H��[�.�ti��gJ�oZͻ�����u�o����'"��`HVQ���2"���NZ��SU���?~���ٙ� �����`��J@�BY��� �u]�#u\o~a�G��S�X�?7�eۍ��juTh��7o�T��?�ٶS�v�\4�0Ա|��o��p�b50��BR�ųd5Y�<^�H^��ж�J�Z�`Ɣ�Ub$":_̯,��@pCɍ���䣓�@+���!�*�mcΚ��^Y]�F�ہ~�ݛ(\`�����7=5�8�d�Z���+���ّ���jpu�E�R���=U�����=���7�.d���4:.��1a����f�㙓W_��h0�`��O�	tY�_�rv2�����E�4�x�͕�U._t��,�|����D��ƾ79]���Z��з[$k!��!� ��O2�k�֕�e����"~=�;����� kzj�T�����P/\�E��m��Y?�����LS��J�X�J�$�=�=r��Y�� ڏ�[�+P�:�#[\Ya�lt`j�hjMf;Fv�Rd�] )��N�3_YN��=^I�����J�d�!R���_8o:6J���Ks����̄�L�M$2�]3t�r���O�/���;`ff���#��ӏ���D��77����	��3j*�A� ?#߿�������'
��no�ϼ��O�H��I_�$1��FU�!�1�*��/&��b�Y�k��siZ���.�oަ��G�F������r.6�z�J�{�ȉ�΁^-�Y�!K:��n��Fv�?���鶺y�R�7��Z�����'+2*;"����YZZ���І�c��֥+W��_Hɑ�z4�O�(B_@} ���c���]aN��5-/����U�7���Qĳ�HF/�� ��{/e�n9��z�K�tf���X���}�
�ĉ��6X�<Y��8 f=Kɓ,��Pdgc�d�y�v:���0�jivf���'
q�%+yP���2�\�@"�@�h���j����>��6����?r��`����~���g�P	<_)m��;��q��ġȽ��ZƜG�Ct�F1#�X�I��c�bj��+r,�Z��OO����$�t�qlv�'�vg�p[g��
┥11EVAy=�}�a��Ƀ���;��b��I ��c2ոQڗ_�21��WߗDI��?������I�\��~�W�U�wQ]ƣO�8-�O�I��f<H�Ð,��O���§���zr�N8��U!eD�U�w$st�/�W���k7����0�,�T��Ӕ�(��\*�Ɏ](���E��U��N�K���s��Tw��\Ы�Ɓ�=TɎ
j�W���^�s�o�&bO�(�ް���ZVQy(߿�W���,`����~�������4���N��Iǣ���x����n�����t�a�'�_�����l��B'T�_x����}�K�����,33�f��3T��窥�Sv�{�d�>ފB+����.�{�l�@�Y�Q�V�>��bvpl�#dC���hA���\���k{d�9ڈ ������>u��܍���R٨X!�eK�3���n�՛,�Zr����q	��|�Ok�Ћ��O"�����b�$+
<.t
t)��V�0711	:,^�0�����g�Qh��f~�%>����y�H�(����U�^N�^�W(��=�tj<%?~�
�a�S/�E;c�n?����l�ĻX����x��%jh�R����N��������4R(#���/߷��"��ğ�h�_w�܁���ӯ /
�[o~O�����
e&EèON��YPG�D�*�<��M/I �(Ƌ��,��,D��2�g��-9gֈT3��/K:���a u���x� IuMy�Þ�� ٣�m�4�N}7���9�=�7����O�̰B���!�jE���t�sk� +�Z.U3:][]�X�liqI��|���=�ѭ�eV	J��.U|*U9v��jK�|:�a����?�FQ�5Fl�X��Ȇ�qÃ}t����o���Ɋ���#��3�ڳO�N4z��x��d�
b�E��4���\r���7��������B5:�I���l�Q����������@2�%4,wB	�O�MeQx ҏ��ԋ��{!!��$����J3%KȮ�8%Ϯa�Q��p�d7&/����j�"�~s� b���4g�,�432���+��s9���qx\���z��C��{b�*U��
��I�}#P���G�������
�hj�����d��B�(����6� b()�sO���'�Iw����^ߢ��ᄼ,�p����RI��2E�t~��]�槠�&��8n<lD�ƞE��+���FY2D�A�luI�}w��JP3��Ԥ�8�h�=���g�j�w��-L^<gw{�>~5�����:�پ{|<<<��9��g�(���q�,��ٹ9��G��䍧�1Fq`�qH��j�ABk�NV�&�iGY���1�җ%~j�:��~�[�d��oߎ]7P��G��H��Q�/T�{1{a��fZ=KYXF����bh�K[~���t�IL�ibe	����P �~�#�MBv�(
-a~��a;\;n	�G�A��t��ڥa��n-�k��S���w6[��u���}���L��g��|y������{q��3y��.���Ք��Tyc����[E�ѮI3��Q�Ǎw^�3r��,!�,FW9B�@�*g���+o��#�`��<%yb1�1�0�0�_����N�5=�콃|��M{���:$�SY6 2��W(W���;rȎZ��?Fn��f�J�i�9��1M��%kh�9ѵm�T�u*%��D��
Ȏ�g�ac.S}�$bE�O�u%mxv�������.�d�ds+����E�"�XvF���9m�5�0�^�[|���w��Z�*dlma&W�-�N�5�aI��$揚�� ��?NX*��� ���>�f����9u��3:��R���_��[[���'����*L��!/��I[ �����Fyω`�?���3/19���T�N\�ET2��J�hP�r~�KOtLS��3����:YS��V��ɐ6��͝0J]���L��B���$C���߭}�Eꌎ�kb��o��?�<���?������}�c�t&f<�`�!�u�D�1Y�z3)�zy~
T�m�$����x��!L;e�y�ݻY��s��}��;z�6�<7��_�՟����/���nK���$��,��*
B�6q�k�
uv�Y>[Y���;��B��?��or�����х0�`�C.Z�$6I�2W�)��8�I�	r��S�����N���U��؂ٮ����ǻӵ�)��d�9	����}����(�����kJ����,y���r�?�q��~p�ƍ8���t��+<�	��)AsxEt���z�8?���x��t&�@G�!O� ��,�C�Ô<&�<�t:�8}�2�Ď�����
�4���Q��ٽ������>>������b��9O(Q?�OV����`�����Ri��� �bE���,����q6���F^UԄg����[�� N$YA��
��/(F~��'�u�7�|syq��:�����;>>�t��|�&k7��m�:/�J}�����ɓ8������v��q�14��YY�������n<�4�3|��`i��˿􋊢�����<�Ⱥf��݅˥h��ӅJx��}�l���FE��/./���(#�T�����������KYPx״    IEND�B`�PK
     �8�Zj���� �� /   images/3281a32a-bb08-42cb-a591-9481e2c9eb0d.png�PNG

   IHDR     �   ��"�   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx�\}��U�i���x�b�$g��gq	�����C��lq$!	H�{2��dܥݻߩ���^ _2����[u�����߰qb�$R�4�V��:e~,.7��C��o����L�q����	#�Σ��W�G0�Gw_?L��ʊq�{b��p� �ӏ�s�C(cA6���\t扰�rhh�����N����xN�~K�?r�C�gr��Ќ�+W�dw��u�?����z��n������܎L֊T:�ʀ�W��E��;���y�Rd��L�đ��4�
�k�5;���"c���������i��q{��CF:>��">�v3v��w���.A0�Ӈ�~����#�3i�����ĵ�H�awy���/��_�t�g�8��\�ǃ�KW᧥kO&a�Z��f�q�0fx-f^z	������+��(�y�x�8��ca�����x�d��	��X�N���<�29'~۰+7mF�̯��pﭷ`���r���^G(����O'c<Ǝ��D9s�nt�x�����̳?����\�e3�WI%�i����%>�Mi<x�m���,<��W���a���v����P8��qq�9W��s�bs"�L���BM�GN;S&������X�r�At��p�-py� �s��!���l<��|��ѣ�{�V���È���3��@-�=��G����CQQ>�a1>�n���sIȯ�� ��{OL�2�2V>w�]��u����ݸ�_W��, o�ps�Ű{\�8\\C�D�ꪐ�����=�"l|R�8}*�8x?��f���V�~��33��F�:QY^M[�a��8��x����'���+_�3؃7�y�^̧.}>o9b�hq0Q[�<��<�ݝx����܂��7?�����b�k��Y�<�8���=����<?ÄRʲ��;a�0XW�� ���/�o �.�U���(�i
ך� KeF��7[PR1_��)T��� �YP����щ�_���~�#�#gEgW'ZG��"Ge3[2ȥ�ؾ�;���pv~���@��	����x9�k,�O��Zln��f�y��b<�mݨ��+�KȀ��E�r�N?%F��]=�`l6��(��N"��m݆Dڂ�8y��#7c��fL�����ISeEB�C0;�!�XPZ]��7<[�y~�-N��6d9��wv�P巣��
�7�N�e�qX�50��[����\K�uX���pV�l�t��	"�N �� ��Åɒ�"��p��Y������V*
�k�Z��Յ�Y���6��J#�0�Tv*�)m�8����hV~�h�9�M�a�a�o�P|�|���zb�)�D��=~�H��9��6��O�r]qظ?���N`dm��A<��uP��dx�&�	i�6�s��~Aqq-A=M瓀��D8�F�oüE�1mڝ�>��xa&0�-4��n"ö�Hd�]LY3�ԣ��PRR���.�Ƅ$u(�J��A6;B�4��>��}|��!�|━��I �a�������9$@�pX�� �t��x��]�\3n�*���Z��>��~^4��`\�a�d��L��3s⏵1eʾ(���E��~.!���l�"�O�Acn��BYI)36m�N���s�y;|<���>�z�U���y!��t����4�W�|DA5���J]�e�
ЩA���;���������"Ը<��gf�R��9:�ݣBrҳX�Wlio���@O� b�?�N ��Qn&M���!����G���F57�������lE��A.���߭T�<��B/�I��ts�$�����0�0��7B���r����u�k��#����-"���	(\�m� �T���PQY�,�DE���ٴ�>J3mW[+�E%H%S��f�L�Qc�Nu聈��R�l+A�L��z�{��,�Ž����9Y&��CAt���f�ш��n��j�A��+)�R��,��뷹��rDFz0�5O�0!�ዡ���9�_�W/h�IQ��A�er��5�j��CA�����3mG"ßoF���f(��V2�A�F���,;�$���	4�$z��E啺���nEGgƑ���*���f�R�Y���� �JG%��iD'�����{v$�y�K�̬�-��$�?��,�-�e���YZ�!@@�{�襬�o\��2Iqm6�G����r�G���|��o�e����gE�4*�,z^b�Vꪓ,�M���>יJ[	����Ee���h'&:�b�GD�)o�Dv�E��$(�<FO� /Yj�l���sq:'L���Qd����+�%Mg�$�9\\C��ɉ!:kS�J���}Ɛ�й�ZQA�&��'3,��r\W�rJ�RikV�p]m���6��D���ڀ�u]M-��ǿ�9Tə�<��Y��� J���V���d�Y>ڒ�*������M�L�����A�� J;HQ�!
�a��H���[12�Z�en�(������3�g�a;3IU���r"���sa|�E^�PÝ<q"Z�"4|��	\�1:āS�QD��HN,��<י'��Q�bт�R032�i�jLVD*܋ �C�.��Fb����E�;��(���?���q��b��
c�P�s��hH��
�����0$��P�L/�G��p���hL�6*�x|�	z?�D*�T�@�4��M!'�4�!xI���i(P�T�	�#k����Y�A	=DfQ4��C�@��:jX�U=?���M��&P��aTM���J��yY��,P*Mp��F��?67�C���9���e��ͦ�}Dx��g�$l�L���!��	?��+��a�F�.�*�a2�<1�~ʱ�4�H�(l
V~�	z�l������sm��\���+���6yꎕ:�u#��	+���ǩoee�
��6�߯a��]��2?*|E�L04���<��E���	:-���fS8 k�0�:��:����9d�4t�tQ�6���H9���\�K�	VC�
xЗ�	�����-�0���L����F�f�F6"�'�K'���@���d|6�W̤PDg�e(:�Պo{�~�Z�*�:�R�ښ8�GNǦ���zNV�1S���1���{z���i�N�oV�8*OQ1*��@7õC��"Ip�a�����k2����z�DK"���b"Xyȡ�a8	(�LH=�z?~�br��7L�0��aQ2�?/B�o/�ux�p�wuPA�������nWAجB�8����.���� %����](ƑG����(EO�=�$r�Y]�>���;f�t��.`\N�"�oP	��bTVWb��N8�9�X}f��f���#���:�T�8�-zAz.2OFa"���~�4��OWy9R;�ճ�z����DW^}5~��&R8'���N<��f�=v���W��w���\��S>o�����Ko}ȃ�Ȇ$�]p�Y����&h�KzY*�x����S	:��>���J+&u&`�H��]8��c��\O��KUQtt�V���s�3_�[H��O�3#�x8픓Ѿk+Մ�v��;��d	�9w�@�԰o��n��>�c�����?�D��
F1� =�������D�dn�8��~ ��dm��S&��b��3���I�kǎ��T���=�X���_��٧���+�#�p��-bHGwn��V������A�C��ǔ--Z��jLC��������\�83KwƉ�͘NґFqQF������AQO��6m�ǸQUhmn����<�>C �e�?�%/<��͛0�л�}7m�aU>�����Fȴ�&�;{�tb����H0�E���_�24�&t�vq�6:4�ϯ�_���q�J�7q�y�L<9�u�n�B��.��������	et~Eu#��#�2�Ӥ�+����#w݌xd���
��}:~��l��+A���O�S�Bf�$q�c�����9r�*���0/>��STԌ"M�!Q��|�?\p�H�;�Xllh���{��FBC�'y �w�b~]�Bo�CF�q4i�J\ؼy-^}�Y�v�}ߖsdQWQ�G��V.������i�0� �.+|��xs�{��ҋ��%m<r�}���VS���^dba�~��]�����;|�*z�4�Fcߴi�9�p��0v�h����P�kKaxA�?���(��Yz�M�v�B�c���f}��7|�	�S;��V���x�w45`�5��~�F�x��|�x{�l����HE^~�U�~�������?�ƍ��n�W_�O�	�i��U^���~��G�-Gen�݅��N(���f<��#�斻�N��ϵ��'^��_c����R��������Ex��q���Qk�·�q�5�� �'C�\D`~��ǰ~�r�hRf2�o~��@��Ш����u2�F/���ì��-[�a�N̘~��<�7��������Gh�tR� +�g�D�^��zZw7��g�Ͽ���7)��;
?��,��}����g��{f+����V�='�)qоq��C��_��qN:��|�t��e�t&�w?�0�G�F����o_q1ޘ�>n��lX��=�_|��<�ټcF������� ![5�_u-��gV�H�s&2�o���e�� �������[�q���L3�KoK:ic��8��P{HHސ�x�����m�І�q���ҡ����-@1���Գ�];�!�>��PA��HI8�u��D����S�׾4m^�[�:�r6�D2؏��u�v:�/��!�[sJ�����6�]�uӵ�Q�l���
{�p���ڄ֝;����[/c7��։�?��ԏ�۶ҋ��È����Ӫhy�yno1���+�{�Mh�߉;n��nC}}=ʩܧ�r*�����p��0�w�I� M�k�̟|�-.��\z�����&:{K�D#ݭ߰��G*^���K��&��àa��Ko��M�]�]�p�A���Į�V�M��]��|8>,X���kӜ�i*~�y�5\t�h�r�yӍX���wnǮ�z\;�x)�-�O (ŋ���ʚ�F�@�@����w?/��iRy��}�������Dۮ*&��kTJ9�<)��O.O�3�Ͼ�1q�l�~�=j3i������̊1{���^f��R���{�;p]_͝�Ӧaxu9V/[�7�{��2eK��z�RƳ5�A�|�`!�SFomRoeu�XQ|��w8�S�n�|�s�U>l$ʊ��N���"�TTb�o�a�U�ʕ�_��	�d?o}�	�=�T�3\��'�s�^�w���u�.2��y.:���`	��19%����?�;o�������]��j�{Zvn��o�E9�������ڍ��nxi2[�4�x�=�,�u&c���3�#P~꩗�Ut
�h
���ʆ�0ܢ{�g�KH�]x��Y�񆫱� S[�ž��g�Ѽ�WRs:L2�[��ƌG\ئ�^���eYM���3�v�q��3a���fq�jxLQ4�Z�2�Sow'>�i1_C�O�T�N���r%�w�������X[�ƊS�FH�ݸ����R\}�(����_�E�J9�d�x��qQ6�ɓ��A����-H�Zr���*j��λ�]��X)��$�%�P�g0��xw����B���� ��b@���˅�n��#�#0�������<���ԎF\���1�&^H� �{�<p��XMe+'}?r���0|�j�ī֭ES[�A�
W�o�~�~7��7ߛ���>#�k�;:�J��q��������Ͻ�&=c�kѸ�������N������CFgO=Y��i���v�T�`���o��_�p(�I�lF�q;�eU��q�b�5�b�� �3�W��������EY�-��%A'Yf���n�7l�{�?��������-_��]RR�>��$2Z�bd>�$fwrq ����7 �G]�p(�*���QW�Y���X֦
� �1����ղ��W������BA����T���jw�\��m�.|�`|�5%��K�dRs'��4����wBd�[��S�m�3̒�Ɋ5�PTQ��+��hn(�sO.��W�.���E�J3G2ՋhXM*1n<�ڛ<�bDDw(GQT�%���K�CqU�y�U<r�mh޹�pE�Ś�ih��f2�]��c�*SJ�Yr`�xn�G��P�.C��N��R^d�τ#�G�~^�D�LS�������#�dg��
�����)'���a��������ڎ�d9�5jE�&C)�MqOŔ�7?.���ä�#�K����J9}��|lml�=T"�L�I�)٥����1x��pљ����
��/ri{B��˽7�����D#V�ʉm&@vT�9_��1CC8�!]�:줬�&�㡧^F��qI&�$a�YTY�[�9�fgk?n��\���4���Z�r�]���;��|��v��C�o�� .S�~�捐`�*IK�Y��f�)�t.ɯ-dù��qi�F<l^�u3v���7m���h6\J|�\����y&����~��<�Pѐ�Y�&��6�x��w�z���5����>��$4)��h�/\����GkJ)mJ�L`�w��!�@�uR]o�r_B�����?%����EK�.�>ƈX��j�]֐��ʉ�R�$��\�D�Á��5�b�E{�|��[Ƶ�Uv����*7)���8J�x�/qġ����b")B3�r��b0��C���V!��`����N#vы~D�7z�������B�n�5��o C(S�c�ʙŬuw@IX�r6t�����z��K��i,M�-(*.Q%�Rɥ*��\��K��y&�2~��we�6�3�������s���ErF"�0��&� �$鱙g��c/�َ KkO�,^��r�ϳ�gw�(Ô�����G����ɀ�Fʈ�ת�<�1*b%��T?d͒W�������|�Lz;RY��P���'U^Ҋf��$	/U��.XT��X�M.�3�~�b|=7��I_�A�0B�2��!�&��������	t�:˰����D�d����i�;e�.������De��u��ʨN���/[�KVm"�(&��I���Q.^:Lb��I�#vbA����ѧ��jS�����=d�NX�o�f�Ŝ�f+��N*m�K��P�(��7���L�����׮�gIiv^�XV.*z^bV�0��T�B�L��q����T�"�M+8P��@$F%O�$}I�A�-�ʙ'�ک+֬����H�5���?A���<����?QZY��Q������ǟ���g;����!�oAR�\��EA�U���ʤ��� ��%+��J����sZ)�*H2-БS%�Ӗ
�U�Ǫ������+�e
�/ !	?�ǭ=V�Y��'�u�����(t�+����9#/VTYM�;���⹉\��99UN��ن��.'uu��]�hdd��5R��3�Tc���<�K�UU �g8F��I��-Veo��Y�|I0��i����ɨ�s�m�"��ky]V�c6�����7�-=SQw�Ӣ%x�߭� �ͨޙU��(uŢ�)��Ur
���Y�O[�n~M0 ���Ye~�%�p|�؃��@����w�oK��HZ
��@�=CF�p��� �KSV[ጲ��0lL�Q����j����x�҄e��I��3�m+uè���Y�t���|���N��C�'M;��
��D�ϼ� 0I�A7ٛ�,���&�qQ���E��k7�����k)I(��I6lT�ͺI����"ᆋ�!Yy�S`5ʏ�B�Jb*�R��.�Ac�U;���f����Ũ3�:�'���2��ܜ _��;���<4/�8Xz)�п���/��@j&�{)�Y�\�N�ZőhV>����#��uj�C�����}���HBN�H��/W���r
�)ਚ����j#���Bi,A�� Ȩ��3$�E��:{����F=��*�z��תa��z�$Ȫ f�[���6���n �(�$ĥr!{u�ͩ�v$Z�F�lH�`𦬂����(�i���yp��S��UPA�?)���_�%����U/D[�b"�"�J��f������YM���ѽiQ�̪�V9I?
�]s�]d�oΉ#2�� �v:�X$̳p(�MI���;Tc�O�������2i\�KG.u�4_J��>���H])i�M%�!����	*K��X�p����{���}�-ϳ �.R	����VGb8T�f)�`$y/�n�N�	�,v�����+o�8#���@+�$CO��:� �#��!���C���"|s�Y�b1s

��&1��QX��.��MJ���K���u�OT�gУʢ����B��a(z�Gj�͉��
`a`��C�r����:G���ƺBA-V���pp���R"�7bA��e�i�y���Z�㉧�&�v2Z���`M� �wE�a���3�ҭ��L6ax9�)$n��LB?3�5����a懃}��b�A�&�!
�?�W��O!�j��=����)�'M6�O+
�&S�+��9�O)�*�I_���F���g	�Z��L�h,�`A���oi8��T�l�pf���>i�2��B����:KՃ�ʷc��v�ƇB�-f�[�L}2����n��㥭ږ.�+)�ͩaI� ͆�bݫ��{��h�.�Y
M|z����D/�4V�%�eQIԋ.h����/��Io
�.@]u-�b��X,�MW�3�:F#T7��j2��A]�kkŉGM�p���Q�?��`W�ft�lh�f�U���( �XK� *��&M��@/�K�4d�"h�h#�sgn[I��Ϋm[4,uJ(�s�����~ꟴ'İ�QIkK'��p�6Q������Y��R*�Ԫmj(�����#���ady�8��Ӵ��A��h�"�z�����ݭ�Rz��s� �t҇�����%���̸����Â�K�9���IcN��6��f$�N�����e000��:Obw['��ڍ�Ē/�U�Vv�	�"��X��Ǝ��;S����*ҜO>FG�^�T}�R�?T;/�N腒�Ə������0¹�v�Ο�P[����mf���KȒ2�;/(�}��$��^T���z	�����@cK��/'F`��nY>CCJ<9��q8�J���*CKK�V{�{�0�7Q1l�2Ga\r��[�����Ey���Y?�`�R+{�L`��%��Wc��C�+K��"��]	��(��?�N�Hx�j���D�)�����N_�*;�ic��i�o^�1�����[��`�n'���QZV�O��
�{z4Գ2����9��vh���������0�vӀ�#�3H9J����/�UT���j8abH����8��o�x5m*�<�d�g(��Ҳr�?��a�t^��
�B�H܂���V���~y��t)���գ�����|��1A�M��H�JsTf�`��q�7���F:\�k����8�������~�"�����5M'-*�c��Z�U�z�Ll�}&�;F� ;��P\]��}�=�Ykgə��K�%�Ij�6��ɇ�ӚR{rS���k��كC?����e��^il�j�$BC8餇pӭw��-Q�+J�r؄s���v<������T�t(J�:�)jܒ�ϊ�ќ��H(�"I�i���&��w*����h��S�������=D�h�Rz�5��[3��1ދ��nAwW��2�����+�0y�x|��w|_�H��X��k�DD_*�W^Y��h��c%���pљ��'��;�}�߯�P9���@�����FT�c����B�׮Qd�Q�{q����A��QZ"����A��7m�݂g�z;�"�0ɞ�#AJ+]ȇ�cS��jQ���g�	���J�c�����l<�=�U�+�Ńx���q�������Ϸ��8�ps���p�1���5���)�	������|�wD,�ҹ&�٥睡q��.ӵ
�
9��S�2p�^R����}�q�;��&]�MM�g߹e#�~�	���Hx�ڼ�Ef���X�S�<����@*���Nn�[i�8 3��i'�g7��o�T�&���QGO����0ς *�!��D*���
�i��.��'�3��~e*(��b/9�l���;����h��-�9��776�7_C����C:�DR�)�Rb"�Go��K�������h�F�����k.��k����Ő���^]]��h��o��z�?��D��%wg�:`��Y��u�^H9��O@��I^+�3J�3��G���v<��F�G�h��b���Ԋ��l��؁��m/ϐ�IB,ǿn��?P�1=n�z�-۷���g��gf)�
Ӑ�F16+�g<�=�ߊ��.�p|���BRL�*�|�΃���R)�"����blN�Q鸔�T"z_� ��N���s�p��x�g�-�v(tи/���o��zݨ��,ٌR2�z�tt�����އ�N�]�&P���Т��}6��x��� PJ*�ʡ��~z�s�g���砤ʉ�_� �pQ����	GI��irqq�~M*�$z�v��'�ǃ�?��X/'I��&ո����{nGg�.�y|h����Y��`���������z�X���I#L23$��ÿf^�%P�$#-Ò���<��5��^R�K�)?�/PA��*ݓd[�28|�}q�ԃ��ݡ_{�r7YV%%.$��7^u�}�u�M�R�S�+� .��:t�����xsh��AEe5�����6�=��īo�'�U���������3�?�PO'|
���������y�	b�^y��5!��� ��!���:�p����&h��bt�C�n�@Iy%�N��aJ������'����II˅��e���<�T|<��-aĩ�ø�p$���4ji䪧cK�t��u$8�W�}�mMP®Rl�و�[a􈑘^U��ZoK^~�I�{�ct:9M�.$"C8����פa��m��r=��>tlڅ1#F��g՛�SȆ��W��](+�b2�������9]���\��n�j��8��+�.[	�A<��C�� �%L�A��u4�瞦<[QSY��L���.$��{��4ꡟ����m]�%��#j1��}��ȕ�ﾝ
��D+���ZLh�f">�G�ʫjk�g��j��!��i���MaLU���-fl��U�{���
*������q��*����{`��2���f����ċ�2��1<7���s��MZ~��q,[�E��e7뽕��rz�!\q�9x���
��D���a�}�I��n�p�;�1�b�}�o��RhS��Pw���q����Ͽ��^S�(R	0�B{�a�C��u�T`��F�}(�9q��S���q�*�8��[��Ho���:=�m/��<�����>�[���(&�;`�^N	@=�@D(��H�1¥�Oy�0	�WZ���lܸD�Q��v頯`�o�M�^���z���4dLţ8z�T+򣻣]��!�Ο}� ��,�����3�z"d}����̋��|F�Q.��Y�p�����Ć��X��7m�J�+�=~�2	E��9s��s%f}��6JI���pѹgR��PZ�g(���훰d�H��'�?�d(#���/�C/����`�������eG"�Yk��K/�?���|���$0���ܓ� ������W_��!���n����b���03������BIi�^i���L������3����sR)~$ҏ[���ɝ#	���[z��ST�;[����x�k/Ng.��\���z�?K�Ϥ������ ����/ǂ���\�H1�����f�PW[�SO>l�b$��<�8������,-�Ƌ�~��]�bo ��W�_V����+.`�kV�s�9gk;�T:�\x�?����!�|��/��epT+(���V|��"<��ݴ��6� �@�h�²?V�^zx�ӎn"�Pt�R�<��iT�8��y�O���T�b銵�輳�ȭ�>�e��r%�qur�e��C��ݾ"��旬\��[���l�{��U睅�P��w`��h����5�=x�)|V����o��w���&�p�r='�Ҏ�r����s��۟x�u�%li��ah�nGi�K���(��L���M"8��i���#e���i;��_��K����w�|�&4<�TXa;��q��'h��p*�$��lݩ!�0�1�Fik��o����o���i@߳���~z������v��B/�R��W�SƩp�@9�S9���W50I,�	�ݟ~�+�q�^V6̍�T��Q�W�8p�I3��,ؾ��2��W[W���3O:ڨf�MM�4�!g�&0eF� C�ҊZ,_�	���\��)�W��j�P=9h�	F�^Q�$/B���r��B���K�̫c��+4���l�o<���x��1!H��QG`��HE�J���Va0؇�#����<��pH������U���/q��HG�w/|���i^����Zإz�'�gp��!K
h���щ){N�cϿ���y��I(>v�H���^�G�P��(Hc�u��w��#?���Q� Ue�x��Y����d�R�.�-%`�f52��#��J���H-Y�9���������q�9���x�?�8C�>mw���x�4C���F�
R�˱bS�Y�LY��|���3l�6���z=�>r��p��F2��	0LK3��{V9[>��w0YL&�.��Ly�_%^|u6��հnݶ��v�q>$�a���ኋ�@v0MO�VW��֬F�� Q��/�G�~DG�A?�G�����;z1��O�_O/ً�Аz|OY�&u�U@;�v_8���15ʦv�Sgel�q}��w8�����-?�"���ۭ:㠼���C�c��e+�4�p;m�i�4V޴�A��̼�"Є�o.퀔
��f�k�=4�ˉ������N���ҡX멘{��^���`�&�-)} �ĔR�$���[�3�nk�R�u8Mck�E�c��;i,�����j�FX�($�&q}0EC�w�}���I��.�{He��Q���Ҝ�V����2����~��Dh8%Ux�����I{<^����Q�J#<����u3��7q�bX�"�Z?.\B�nזo�P_?�<�y�����O�ɡS����
%�U��9����J���0n�1��C��ړ��=���7L7>��H���Fe.N`�̾\K_�n��>�,�[|�o+Vb��c��?�#��+���,�ZawR�VpI~�щtu����`���Y�D"���[ޅ!�k���NJ� ~/�CTIý��b��=�pm*�ѼK�C�߲��`J%����Sn3�]v�t�)C;�(m�@ Ji!Ʉ��J*�;��V��X�V��9Ȫ��:���cC�:��G��q�� A�G�؂}��)�VUhk}��='Y��8��?}�\c�ܙ3_���٫�6o�LĄ������\g�Z u�� ��wW�|��eI�����I�I�N9�p�jsy5a�W<�GX�h�b\�[�\H���h��bu��)3:\DҴ��(�$�z��r;v5btM@��c��m�Ɛn��K������Mj��9��Q���ooߌ�G�Ӈ�8䐃�l�Z���:��0d�C�����.�lFeEzLJUh���I(A��g(��[Sx�$���b�ɘ�sW���F�S&���8��Ƀ;2S6�����@O�AX2��$�U�u���
�BO��r�ی�-��q����F#�?I�&��L�S��ոw���WkBM�ANzi	�D�Hy��n��=?Gr򧓟���-A�S�wr��Ɍ��RPA
f鬴���ܓI�R��SXJ�`N_	�].������/׆�࿉�K�1Ig��ؾ�ԇ�Q7r�5�%M�ș�t&a2�"e��T��
K�V�I$̓�&eU�x���R�C�Y*⬆z��܀��;
%�"=KI\�M\i�ƹ��N�+G ���n�j�~���K��GE	Yd�T
��CF�2r�UV�!�z�����SD�qi����D�aF)��(�\�l:M&'�~M#�9��`�YBc3٩o�Ϣ���b�k���Q�H�J��/��.�I��G�A�a'0ɐ�T"���!�W�QJávg���HU����Ґ�&�ePA6��y�qASdZ(!hұ�3(��э��^,��T�	��Ր=����.�����K��2���ҒP��b���ҕ'I&�e�� �)Ԥ%+Mҹ�Go(W�3��8�w�� ���v&Z�!+Sh�2��^����u��Ӫ����n�=;��>�]�l}J���,��c����d�63�r�zY*�16/�٥|l2�-�}��^*� �ej`R~��CS��TfC��q���am}#�j�01*��D����� ��cq���C�֘Tht���k6ʥ�%�� )��Z�e��;:F@��� )�On�r�*a)L:�n���&�si���A:�>-9%���� �t��F'��	���CR����n�V���F�V�+�]�0�������3����( �6�զݶ�e��R�Qf)��?o�K�/�6tu��Og�P	�҅.,�èQ{����]N�Y�hl��������K�T���:	`��$���/�h�Z2R���'dJ��̌)cX˺�L2zN�d)�qqq1=��U�kY\l@ �l�* �::���fe\D�O���tFM#h�Ɍ��=��bd�f�N.����;��e����m�&-� �&�LDz.&���`J(S�=�	�f��/�a҄	�Z�ɾ#:�O���!����'Kr�������,�Y�ۦ՘)���e��)@������
h��GI����x6���J�9�L\��\$�4Sa��X�����ssi���K/p9�p)R�Ѥ�TH��!��"�uD�!�̽&�ç_ϥp�������{���ı��h�f%���q�2�M�	2�B<TmU9����著�)�N#;�ho��q���q�wi��+�̦�?֬�H�����&i����:�^��qw�t�l4%�l�cU�~�&��R�e8�6r׀��+�zy�y�

E���TBf�X�9 VW�!&1�ɩl���z](VJ��U���p|��A�����q\C����n��i%���Qmu%�m�J�`,ӹ�v�O�,#����iS����h�$iB�(�J���v�J��$a���9��\Dv&���ܣC�-1f��Y��E�./Ş�Fi󙰯��aF(��=B����yg��'^�X�zm?�J�y��밻qB�|����}�~���Ӛ��܊��ܓ!��ki��NV��[g^�H�?]�e:�N�lebW7CAi*q�'������[��#�Ѡ�:l�NZ��L�IR���n܌	cGs��1~t:�|�G����/ԇ뮿
���4d.�M;-%���v�>�s�)�v���W�C���E��Ҳ��^�,]�ݼN���(F�S?c*�m� U52�8�>�O\t�'�p,�d�N�η�+o�2�����^ڗ��)�;q����u)�M�\'�|�=2ZӦ��2���
]�;p�ݷ�cw���h�٤=�i������q�(M{���p�Y�z�z�B��d���'�KG�e)�-;v�[Z�t"��3�Ӌ"��A��s�~�]���Gj߄x�H�|�-���{ы��d�ƣ=Ҧ��Ԍ=FTb`��?x���v-muvv�K
Z�0�䓎� A'/M+�2��2NP���^����5���w1<)�a�B=�v>�!ո�uh�Q����i�e�
6ҭ��veʮ��7^w���;�l��s<�p�0���r�ܶ~~v[W�*��O�>0���ظv5���x��9Za�<%�m�q�ݷބ��Vi�w�������'��R�����c����5+q�y�㳯��u2��EeSKZ~��g`צ�6b6��9��G�0aG1�P�ގv\v�y���:zN��\<˦�5���܀�a#�حw�-������������b��_�ٜ�p�]���@�4���<���BGS=c�$c�e�/��6�f}����q�a��av�X�j!�
:�0��+�Ǯ��>QST������:���a��_��OE�r�y�y���7,\��,ӥS����vw����y���[�T)8'�R]W6ol��yp�QDZ���H/�)ĕ_��]�S��	���6��:�%X�bƏ�����}w��_~ŜϿ"h;0Y���܎�]�z�A��4�e�R��i��qm{C#�M��8�D��}9��e����~���=�kI�N�?����T-�QZ	�����}7���-45o�m�^���Ė���H���~v�[G�3��^�%��Ѯ����������+��2���Ӱ�����hnk��݌��O��ŋP����W�'*K���w��btPI�Wo(�o~���JR+q2�0��G��s�<+[���}|�	�E�Z$��8x
vl�c�O�/̂]nij7��q�O<�,��z�jc���ӂ��^��p�=7aż��W�� ��~|b�y i����$e�b��_��Oa������ߗ����j��5�]����oѶq̛ﾏ�.� ]m�������c��Fxh�'�pj�c)0�������I+��&����q֙��G/�'���S1o�2z�|��]r�v���P�r���wQ��~�鹁ީ��9bD5jo�u�5���_t�ı�q���aê�uX���g*��_
���p?=�8��$��Ji����|��g��t��3����e�r2�b<��,�f�JK��ko��fj�TC�r�-�bѯK���>�����V��c	>�~�5Jx w52��d����'�mZ�7ᩇ��U�@��>}:Fו�k�zu|��W��	�O�҅�lߵ��B[6�oGM��C���u�&;p��G�Jo�#�k��^AYu-d	�[�ѳ2�ĜO���k�A�������O;�(��hڲ�l��0��W^�-�э*!������tn�`�3���/8_[���S�A���q�����x��:��8&4���ᵷp٥b��[���=�m�Rhݵ����K.�%�Ոf�{B6���_�O��Uj��0nx%^}��]d	��hmځ�}ɯ��qw�v�˟�fI+jG�ƅ���>t#z�v�+���I�H�'���ж���^��<��t��Xam�5��«�q��7!�{7l~�{�5zu��q'�m�eq��۴G4���p������A6�C!��f.J+j�9��%���@c� ��n>N<f:��ő{��?�?Bۋ�h���72^���w>D���.B�g��i�`��Z<�����b��^Ɖ�6]���'�#7X77u�ǟ������.|FŰ��变1}*)�k�D�D��"� ��[�5\w�G���ϑ�j�E>C���u����oƥ�8������Y�OCOo7�I#�=��k��λ0�i��Tr��b�i��+P�Ͼ������!�R���9V���HZ(W��C�v_7E�r���,Ui-�!:��m�ia��G ��NjzHZ��\�hO�����/���J�CUr�i�F��+o���C�u��i��M�D�s���[W,Em�p���GH�]ZV3��H���Ͼ�=���ձ�����i�Q�Bh�}�浺i�l Ӣ�f��?'嘦�Ƹ���-Ź�����Q�5aҡ�؍��]6lm��K�QQ�ڌ�&�v?����sp�5�!�s�!��2^���$�a���zÇ7*/2�[BH� ����ï~�Y���M�ٽy+��$��E@F���g6��j�|���#���ɳME"��v�Jk�f�8�^���Ǩ5JM�T�|���s�N��Ͼ���/B�,�c�V��Ś ����Lw��W�V���d���%�}�l�2:淿�g�vJ�6�4lG%�����2���s-�/d�r�2b�p;וg�M�j+)������;����\Z�g�G���5��3/��ʚ:7���:n�d�]=����]�a��1�BAY��l}E�(q�=����y��hH��u��H_�0_�G:�%k�P��\t����Vc�!� �ߍHC�N-�0��1�|��O��C�_HZ�d$��"Y<�Cy�h���;���k�E���(#��k��ն6l��EQQ[�x&��2�W����eĊ5���ɨ#r+���.��W�I�Y����v: �p�Q�!s0d�q~�~�+.����;H�%t��w9�g?�չ��DZ����M¼$��ǟ{7�pѐ�ܥ��7�;+k7l�2���1��&;m������3�7����<y��f�
���e���2A�[R^�(hL��-a�0(�b��_~_p��a��P(�7-=dK��H*L
m!���/���/�䴽�/��.��V�8��j㿥t��ڑX��7�X�Vˬy�E�����jI�+K$y���p�5W��j�
"-�`X�ͼy�qni��F��nK��ZA%=����ǅg���F���>���V�~Z���Wk\m�"r��pwG�aq۱��~���]H��5xlh�`��s�G�H�C�D�����HL�����(�,÷������#G"i�y�a�&@Cc3\<Sɓȳuj�����t@�P���=Q�Z�K$n$ӗ4���s6�:_��/�4���q9���}�I���3F�iv��ə-Y�N���#"�z��Ԅ�F�Kq�C���{���Evۅ"�����������X�WFR�)�tQk�sN�8�s�~��y��3kv��V���^���+��k}��T�:��d ��nܤ�RI�kυ[�z����D�K�jº�z���`�07���P4�@y��+pj-�p�X��������<���:$8�����(�s/'"&�F)���ɤ��'R�vx�zUz���X�f;�<f�HW�G@n6�PEdD����C�
s�%��Yq?�+�(e���!�-K	��p�P��ˏ6�k�th�ށr��Ͻ���Kː�X�Pf�����K�L��ǵ���`_)�Y��V���ŖtR��W�a��2�`g�ޢ����vrƀ`�l+�6�+��^����A4�`H2���V}�["gg1�S!��J<��+���(�{��[�q_"�
�M:8��9���u��`�"�l\��'^~C'��=V��.�bq 2._@R�
I�/W��*�dRu.*�s~ZH��W�$=A)��G��+�|���zɮ���?���C��`���H�ڈ,=�N�"��hPv~FV�O�����v��t�ڜ�>5hl����6�I�[rsL�1��L�����^�)\�4�X(�4udg[�^h��*�	����� o�Tp��c�����B����h�ܤ�j�|��L3�����J)()�n�rʈ��Ȕd��65(��1�
�k�󋴡-���睈�VNŮRy��4�5�����&�FBc)�Ke��,�5f���zZF�T�����Zz��;�m��с�*IG��h@�c4��=��&���ieU⑤�譨�nҡ�G#M�øI��Eޘ;��1�y����/?�Hˈ�S���x�2o���S^[��p-ޘ�e$�$�WV�5pO�EH�$�\m��0ʵr=<o�7�rx�E(��$(�ht��~�Ѻ,W�u�[��br��r��Ϲ|����\�> ��gL`�Yc�2!o\���Y�ָߣ�c�P2eܴ�;@��l���K��,��J��c��詤�'�煵��8�LIs1��>�I��TY3�DR�4&/�����r;S����UY
���`Br�A&��eޠ�������O�h��!��ʧS�t8�;�k͊�Me���
���i�^�M+E���{��/��EN&��~b|�sN���.�����:�Ŭ���u��ZNg�?�Fש?^����uvja�xd�&2�6��uF��M'j�A�Ӿ������U�nȘ�\������`�(�W�,��%�h5Y7�M�?.�wH.ˣ���
�?ubEaR��Yfn�e~h�0Ǭ��dV�aMK��bR��&>@�A�P���F���Kf4:��ϯ�VjAތ�>�1#�L!�Xt���c��3��3��xe��D&wI��CF��ut��g�YSƸ$D ��Ò�J�l�d�{���ݘ3j�B��8���99In�J�� �":9�BH5Ȯ�L)��ZF��X���
�B4n���'r�=Vc�K��æ������L�:�?����'��arT� ����9��iͺ���V1�&T0"QT@r�a��y�g���t�ש��~��y>��W��~�_�:Uu�����4.HH(N���*J�]3�l�����HJd"
K�oq����]~�W'��^/C�#rF��f{>Ŋ�ټ��1M�H9f=��hh4�d:�\iC	�}�&�3`���n`���稠G��Ϸ7f�X2ݷ,�ғ+g�%O��ƘIS��t��_gQ��Ü0�x�h"A5�^�*m����i�� ��a���RW�D@��x0��H��b
m[l��5Ϊ�����Qj������V��V.�R��&�OTCx{�C�����0�Lp�������Rhgz�ax$���\��bθ�kڢ۔����^!O�]�-��fō��,A�*�����1��R�)����E��'�|�W�'�Qۤ��99y���2��$!�9�IEa������Q�,O:��P^�������}��y�
E��R&�ZL�UyȘ|���L��c�]��]�`H*���Ő��~��a*8�J&�w`i�1|�/_a��d��:2IC E��RhkiT�7Y~��t� ����<�i�7d-z`z�����hWjq�����qm�Eb:;�����b�_"4�]��Ei�؝�o�7K�=�gQ]S��B���tX�A����{*VB	�4�'���gi��:)���ꍈ|ԣ!�AT/�4�@[ƍ���D�����^�^ޡ��mGcY��jǦ5)�K��؄��|~w4��c<>���OA�K�2��4.��
icc3N�<��Q�����=r^{�m�-��-�������`�ӣ��A������44H�����}r��&%3�gdJ&2�JvA+��f<��}u�)s��}@�~����9�Ll!�E��kȧ�niJ�1`��`�ԓ4<�6�#)�����c��Ү�P�_��Z�ӿ,7]}��_�<*�����o����\���JV4�;e���x����YTȔ4�8�q����b�7�l�8����3���m��x���0��_�>�[�V��c/}�!X�}�)�R�kds4ƍ<y�!7?���l�;��`�p�_A1.��|���*��jK\@OQ{������j5.-nZE��62Q&�r҄18�	�[(),B4��\�e+W�U�T?��`�j�V%��I^|��p�I�a�钍J��V��)���'�K,���aoT����8�9�9/>�4Z��5��x�b�����|� uu:��X����#��[45��;n/.�\,rww Y�\�-il���_}�/O�E���)��UB1�$�3N���G�8��r���J4����̿_��/F����ɄALS�+0��>G��4~�1E.��vѧ��n؂����ʄg��qd9L����z�>]ט/%�%Ɗ0q�qx��WPTZ.�oH�sPɞ9v��b����v�8�FMA9|~����'���>��b��҆����)kЁ��`׷a�%e}����ˉSx�������ҹ/���* �Z��Ё미�u5R��X��C��ً�ϛ���^8܀U�a 8��<�D��,O��a���e����+D��JM
�r��xi�;��j�<$��5�N&��A�1��ш������Ᲊ!�u��p�s]�~��ga'3�I٩�(n��.	�Q��Agg���s�kj��?���뮚�����Vșu��"nBkC=��N%��)-CSr%y'�=�퓰z��/�1zwGfϚ�!����-*Nꎨ\F�ǁ\w6��#�VﯔK���
�x���w׍W�����5�M��V�fyN��=�Tt��ȅ�p�,D���	4��߿�y�}��]
�������!��oF(ԉ����su�������:)/A���p��M�2�C�p�fҨ��R�9�1Megk�XĤ�2�a���Y��>O���K
����P���l1H�]s!*wosVnƸ�N��W��%3O�Ɏ0M�]��S����wuu4㮛��)ڍ��`{W\C�`O�6���d�sg�EKT5*&��a�O�*!�,���W�1��Q_����$���s��Zp�M7�շޕ��W�O/�eON��M�D��c�F[�}����G�▃��%0t� ��t�rF�fC�XC���v��8�{+
|��)G�\�R��nٟ;����9첎s\iK&����+���^��s�ۀ�9��
t�n��4��Ot@�I�Ϭ^��=�c0n�pc�ɧey��X}�X�ʭ�{�l���k��Dy�2�u
�:z�s�GJS ��I1�Yw�\��v\}�X���^]���d�W�ɘ��%�kaO�34�W*F�/�ۍ�RA�����=���PVi:�c��	";u�8L�4NlNPPo/zű57�M\[8"w'���8I��q�v��=H�L���������%!fzd��U�c#gEq9L�F<�؃x���.��݉ެ��q� �'��H�s>n��d����hs`A��]<[�gk��3�wHrr<�i'��i'�Q&hi�1رw?���п���2�@i.'d�hW�/;K�UX3�WǺ�u�\�������0,�)/:���N��N�-iA%���o�й�v���f�{b����ߏ>�d�I h\�)D��t�����0*�շTI*�r��6m��;j�vC.[�
.֦j�A�li��b�Ϝv��p�3�"$ߙ�e#Id"����A��x��7PQ��h�4A�Kf_,�N��8�;A6�RR�0"F�������G��C�>Ֆ2��o�Qe.�ݬU�ˍ��IT�P�\9,�xD�C/�`/�U[�'�Do�SN��$\�:��SA]SKD�E'�'t�is���}���C�`#��SB��g�k�$<�$v�ݴQ���E�7HD��v2~�s�[�4����^j��|�E����4c��-;��㗐�'��a�v�M��_���Ee�CЄ81̜�SB,��Ⱥ.��dsWD�es����Cw܀�_{K��U�KH:u�D�G�y�:֮_���C�I��N��[��m��>O�"U*�$gÝU��n���9y�ؽm~��G99J��r�(�=��7;p��-���"�b��,�؆��v�Vd����a�_���]�b���sg���G��n��o�sv����tu����F#ah
�e���?c�έ:������'c옑�ml��i'�A�Fe�����ttw�s� �.��ù֬[���.�*�q���S�B��Ƀ�߆���M蒻��W��,	+�cI<;�5�ʻ�x�-�1ܬ������Q m�����M��gr�g�NJ$!�m�����)F�7q�┟y�Y�vX_y�S�	��Qw�v�XEN��J\���?���G�����/�Ԍ�����Q+��|^.<g��Rqt��e{g�'Zc&)&�k�R���N?��$�,Z,-*F+�S�g�}��J���8u��)bw
"��s#R�Հ\j�%���8t�^	8%ťȲ���0�e��;n�?�}�Pe�.	����Jj�IJV��?�Z;���e.���ꅿ�������I��C����x^x�:�^Y�C����;8�d7S�ۂ���SN��_��(z�qxC�PAf1�Q1�Խ�����z��lt�p�,�Aͷ\p�|*�E��r�B��;�\�#,kr������RSۑS��TĴ'(�p�̳��˯j��h���W̙#^�U;K��W�A�����ک����?��?ǉ��p����q�jxl9��y�	jh��q3��-��ګ��1D�/;�o&;\�{-��`&^��m�W�����Ç��%�#���'K�}�VtȻ��;zԱ���|%�u�6�OI_T�!7i��K����碭���%���?��erV���5(d�뚭2�q�<+�`f�8O<���C��m�N���Zq,&�v)�K�o%H4ۋQ��>Z��9�i���ư����3�@Z��ȁJ�����{�ӫ�X�����K�i���a�'r��1�S� V��%gL�k2���'�}{UI��BOX�lD�bV}�=��Jq�&��u�+AJUX�K���ҲR�ɻ^y���(�#@�~}���/�'�	e��܂j�v1n�$Ӭ�}p�)�])E�|wm{ }�>��V�C"�߮���3*��JγDu��O�7�Cog���e�1�\�'G3ݬ�P��?�\��P
�M�r�CH���]�F��O9Q�a\.yy>tŌI�(�t������.�7���e��ų�W��(b]�H�D1x@V��,oQqq�*�sΪkVn�ު.44v�LZk�A�.��rT����%�P&��
���-p�l��ExG�ġ���tq|ǯ��=p�%��9�ɠq����]�^���r�)�VZ���Ʀ��q�.8��,?_^R�]{`XE1���ݣ==�z\:L9�8_�Xv��5�^}�-�R�Y���~�X&���&뜔�|M�%�L���(�;�ZŘ�tfnD·T�D� �N-w�`X��NF1��eBa�"6�I����iv���%zY�~Y_^	�X�}��߷��Vj����"A!1���l	)}x�OPY�W�x��nm�ߺk7����<al��B�q�pSCJG7�K8a��b��-�'vA�:Ke߁�8�(���O8g�$%�Ժ�A�����z%IZ=X�lr�+����dT����u�2I�a�}*�s�{0�$G?���;�E��u�\��8a��`
<6�7����Ymc-F3���fqt����>+�\���L��Y�f���0r� �Y�J�K�>
�}Z-��y�U�8v������h�(�
��/�v����%!�"K�	S1�jQ펜<�����C�WR!h̎4:�8˗�����5��+�/�-�ݻD�l�\��G4|���.Î�YB�T�u���ښ6���7��6,^�+fN� �I�W_#	�k�"2I
$���wG�}O�v.�s��U�$;Q+2����k����Y8��~��Gנ����Kkoǥ�NW�j<pUҘ�Ne,���*��/ю,�W�v	��z=f�z"����jS&$���Un��>�Ƶ��H6�u��ĕ��,��U�q��z���|n�]�P���]�p��V�{�Qޔ8�Y�'��6�1P�蒍��üޘ�\y�X����_A"�7O�Nn�n����a�+!�e0A�ܐ���Yݱd2�U5uغc��\$Y)b�jGcK;��������_y_hh֎W&���b${<�~X��)�̨
�uZ(-�괴��*��mʛHjo�W���b !�o�v�:X�"I��1�����+"!f+ g�������Y�Io-��H�VZ�	�{U��G��Ɨ����A�5�Xu�0B�!�@�0˔6rS$�l�Я�@�,���Xz��Jvlҩ�k�);_�;�Ib��䒸r�-��"��6�ܠm�$��^��cQQ���G8d�,�2|�y�*[J%�6�w`��)!)g�8�D�h�y.����f�����YP�G�����W�UX��8s5�K�H�=��P��n���FLU��Zݢ�A��%9$t*#�)���^�İ���9-2q�՚P��U[A�3}X�Rf���f&+�B֌Sy6q�eIs�t���6I\!t�$(NB�!d$$��%��qw����8]l!=	�-�]ͼ��L���*��C�8�8,��������7��6��ꬌ<��d�x֘Zf�ٻ�Y�3I�2��2�Ę|VKg�A���D,�ve�%6�u�t�{�e�2k~q���4�1��0J�p���i�KKj���Z��ӕә2d�G��Β��]����Z$N�Y�Nw���q��RS��q�'A��Y����
��j1
�Z͊�ٓ`V����˨{�Z�g��dr, �?�c�0�*E`N���P�����h�W�J�'[�ru洆t9ٽyy:	�m�Vn��8m�áT5r2`�#�x�l:�5`o�I�0g��C62i�d@���,�	�95�\/Ow}��J;t��ͬ��9�G�1�y�4��̥~�����ĵ�-*��K��{!�Sލ����ܼ|E�&E)���9>��=������`'W%a8&&�m��)�F����r��+$3�ڤIbV����.��d1fژ9�X������1��'F�ߝ�.Wr-\�9֡���I&q;�%N!m��Y��JYQ�D�������:QJ8VM:��'�ǚ=����u�( ����%��T��:5�K&#,��)���]�f۽��v�9��g3�rr�>%�-ѫ���ޓ�[/)[��-vX.nBEL��ON~�����	r�t)�7�V�ʣG�U���cY����mR�ꐋi��TxgFB��V��6�K��3����~�TI%?�3tx2T��\iT�8s�V�bI�����":��Z���J�_��권�wR=�#ˁ|���v	��I���0{t�ҕ�U�|�w�l"/S�,�577����6�,����n��c���se���¸��J?��wg�U��P���nُ~���v�&�t������W��T�%"a��k6��a:w�}%,�� DnE�7����|NqI�z'����=�
�Nŵ4����Y""���^�
1q�KB!�#����u(RJ��r�é��ꛚq��S��oċZ�1֦��	��������jB]��{r�Pŉ�m*L�/�%����Vk"l�Y1f�`�ڵK�>,�`:e�V�mŋ�x�1M�4�j�٩�Q��lX�~���.)+��]�=b�H/,.�߉�?��]�cM,7��)n��SO��g���Na�E�nH���|���D,Yi
��<�-�"�ǃ��9M��)nDt���io9�ݪ��}�I8}�L�d��(2E��s����#��@��r�&�N�Q���u���GG����1�������8�n	������g��.�/d�VBC�@[f�p� ��q
�8��]�����	t���.�{�.KV(�R@y(�l'0vP1
sNv�
рg��#��D�=���a�:�[���ltu�UQ���\�뮿���CbU�x91r�"<����ddIHaL�z
~[��v1\��t�$1k�I�l��Ɖٝ��(�3HM$e0K�ĳ8��	J�EWT� A�	Gf�:	������i��d�/N�$H��Y���t�8l�}P�(�6uY�ĈĂ8��	hm�+�Ӣ̀�d>a�ۉ�lhC��-]8o��b�9��"T���z�P;0��͍��S�H��$5V�e���z3f<�|��IQ4�z�yn9�8�=�dԲ�.�f��e�)��.e���I�ڊ��/�5_�a�r?h���\��zt����Ï{��oFUm�;���|	��
�~�9Ĳ��!�7AY�w�v=���C�����5��1p�g[ŀ�đ8���Q�	7�����o+V�9�r���N��� �d*���+#*��Ƽ�llط#*�(>�G�Ͻ���lA²i#G����NAC����ٳ�l���s�WB�D��1�����w���%�"�	�9��Y֠A�I{W����$L�����n��ǏA��?���W�?�K�]�Y;��gLE��>���ҭ\�Z�)�v�m|��7�玹hk��3�=�"ĵ�aU[��=�6u"&U�P�����lۧa_�$�\�C���=P��ŀ�,\5c2�/�a1:l�lh��7���׋�4�����|��H)NK�׮�I'L@}�n��ޫ%�Z��6�m�B�ׁ�����������Jw�v$)'��v��ȑX&�٥Y��Q�K�}c�l��q�ų�[$qޅ��Ţ��������a�٧��^��`X��Z���#Y@¡�����.����̣�胏P�S(G��=����q�]g��t��p�s�����EE�QG�� _Q��� 6��-��%.�\��O>�C���;v�DoV��rѳ�X�i�u4���G������`D��n��D9@��.�V�[X��,�w���s.�X'��sƙ���{�F�_��&N8c�.F�U���͂\�ri)����;0�����zЧj��ر�F�Y$Ba�O>~voY'���ǟ�+�ë�g��@�^�#��歛�ȣ��e�a�\�d��Kp㵗c���p�7޸e��ˠMf'^��:n��|ڛ�#q���|��gh�/�u�sQSyP�CX�������wd�IsG�m܊~e�8�g3^}�,����F�$0�ܳQW�W�TW�.[)^ӭ�Gd��Q>�t��>�M�s�@�s����R< �rq;ۚ��E� x弆)�$�n�?�9�PZR�x���s3�ڻ�d?rH1���imCia)������p�r��D%�4O����ؿm���NT�yڶf=��&��ea{�Y���ބ+�'H/�eb���U+�T�ۨ�ÔA��Sw�@�1,N*.B�vK,��f�N��sp�"1�WT��^���}H�N�r��*|LEűY��P+�eL���%:���u6P��Z��G�~��N�����\�.�PYuXi��[����=
�܇#S�(�C��'�y�>� nێ9����(�߂����jzB	s�`}�޿�whb�C����%*n�j�.T54#��d�����⽅_�+χ-�;�KOܡI�H��5��vaJ�-�S@�
�r���S.֧_|�;n�6o���&���ٚ����ڰ���5���Я�9�9�ݙ���/�-7^�6ِ��F��gh�!�];Pu� z9Tn݅�� /ϧ�(��۴}��т�q4�݅��E;�r!\� ����ml������-Ԛd���	��`ɏ8m�d>A���E�\z�X�CUUh��Caa	���3x�}����J��_�5n��*�?j.�h:::�uHR@�ž�k4���?S�ce/��에o�"*�,/���``nfb`�5,p�v�6�b�hŮ��Zf;}�d4�9=f| �p�������l�i��Cy��� ��؄`WD�=_~��v�ڝf�=3�W�ۊ�.����[�bL�B�8v��v�]���H7_|Y�66e��6��/��7��+�@ՖM(���!���e�V��f���ㆵ�Ō�鉨�c�j.�o�y3�T1���C�GQ.�.�T�]ɽ�`�3>����"�Ca��a�ԕ[��_�/����$!�ێS����r�V��K��ҫ����H�l�?0���4����j���~��{J79�Z���IA��Y�]��rƜ�!�
�ɴe��Ҿ��}�r�r�^AÜqg���x���h�0[U���j~��TY� ʣ��Io&�s^�8�}�Jw0x��A��e�aK��I��jس���/���F��
���Y�%뒛�Q
o����[v����$a4�ߔP��۟�)���imB2��%�Н[�w����w�{qP.)��@	�Σt���ˊ�/�P��M�)M��.��⍷����CCM5�myh��]x
����<A;.j9:�٦	�3��ڛ��;Q'��+�.�0�m�~	��6'�ܾ́�x�"C}�%�d�R��9��������{�Ś�%���dC��:�oa�Ҡi�MI���"k�!Frɲ_q�%s�+�}�\Rf̙(#I������o� Y#il���UIV���/��&�^��a�;��k���g,�A8��FP^��>�&�>N�H1a^�=��bT=Y��Y�a�JM�q�;k�܌m5�q���9��P�x{�>_�{�3�H���<�%�<�V�ؿ�Z�\��l޲�Y��3�_ޚ�Οq��+3z-�A�p�&7���]M�r����`�!��O���W�`�IF4�i�4���Rr��h>A[o\�Tu8�gcu�md��,�a9�̚�<�9��<��w����X����j�r��$��7Ӝ���*�������q�՗"G>;I��)@^V�8����S��vl����z��l��.�a	�=�l�1�F^Gޟ���z��"Y��:�F>���lr
q���S��³(��Q�ܺ�&	��b��W�~��"B��Xv�d�g1�.�/k��g���<sܮ|��X����Q�p�=�skhՁjoE��5��B?��;�ڼ��9�0���ь�C��Hֆ��Y�F�]62&��f�6����(�?m4'��&���eC���a��0x����sK�/q�\�/���e}��T:��m�C��@���X�շ�� ��P\\(�	�Vn��VH�\�{��r%�+[ ��w�ǀU6��Ï={���xcGZ����tкQ^�	�&����;9P�&M2���G"��CgoS�o�_~�f�m�b�����ń��Ũ�w�����k�_K��ތ�69���j��,�L��~�v�ʃ�0��x�}4�y�z��{�$Lh�J��6Y/NqO"���,=;�����.b�ckwU�����BC!�Ib��L���1��-�������L�w�H�Q�쌡��	������ټ��^���>_ԧ�Y�\��!�v3��"�`��b0ު�hʒy��Ye)��hc�dJ��
��8�މ�fhL=7Z�� Pׄ��KQ�Ӱ*�;5�e�q��"�Q;92Tz��M#?F�$��'��B�y�L�=؆ϻ��3���?icb�ޅ��S�rW���a�o�cɏ��U��,�����$>2O���E��[.�����ID�!��bU���$
�˵���#�{��#�O������b��TM�f�������%J�׳��5�T��8�QV��9H��~�i�����M�����^Y��ۣ��v�*_QҜd2<�&CK�d�f��̶��'e��n�>��������q9��r��2RgЊƑ&`n8[sٕj�C�)�wՆm�v��d+c?�8��Hs��U %�_��`�UM������0��:��Km�xW�"m.2)�V}��`)�R�����NV���	�ϧ�ߦCaR�q� �h��(i邾���{q�!/3�\3c�������]
�Ii�dq�>PO��|cNiZ�(����D����_��%F�Y}9�i;K�,�:�+AR�����I�FG:K��V���ˈ����V��T��"�^A3ނ<�Dĵ�7�迊z��Z8B�5������%����l����m�skW'�6n&�����=�� $�I����n�G�S�f��4֑U��8���iJ��H[T}�茸"Ƌ"N�E�Ҿ^u�RX���q=-rC��r�]�>���[�ҿ���#���,i�1$�]���J�K�L(�����xu��TF{�XCá���Y����1��&�9��:u���cڔBm6D�tV�դw�B��l���q�U����0�2Nj��ș���V��^�1�<i8!���6���3f"Tg���������5,�f���r)��ߥj�-ˢӤt Gβ,��qU���օ�ڥНЖ0O��ʔӢ�x;�,�'?Ŷ��qIRF]<e1�6w����6���8��3��Z�4�ݘr�,)�+Lɸ{�P�Y���v��βPlǪ�_^�%�!`hb2�q^��2��1k�fNۑ����I��l�cC����E��qP�Cv&/�YHu�dw���IչL��a��au��)��H��H�vyj�$ӆZ9)�K0i�Θ�r�a�:g�j3J�)��(7���7�fB�#���j��f��A&�!N(��H6PZ4�Lk��smL��7ВI����g;�܋,%h�U�5���Z�MƺY�I�]�2ĝx�ȯ��#K�ӓ��.�hoDϋ����lj�pƬF���3Y`�>=�2*c&C%uD��b6�y��Oj�v�ku͙u��JF�Bs1&�i�5�HJ�c���pD�^b��1�U����!p�t���i6d����c)H;`I���)h�J�O�ʈ?)����gR���(���Ø-�!B2o��@�dKT<�˪#�b�s��RQJ�u^"�wS�yB�9��j�LbQ9��&l�)�W���3)����DۙQ\�qq�G8D�]���T���X��0%���"਀l�S��|G�%�S�O;�C�z:څ��T�d�17;W� )�c�b�����eߩ?ˋ�CJc�Km
Bf^^�hD��E��Jf����h���HM��*��l��J��$�N;�0�)ei�e���q<�����.�
{$$J�u���ݘeA(�Z�N��l�G�F�q5l�4��A1hZ2��P��K�z�[jй��+Ǣ1�H�&K2�����\�DL5I(���f�I�
�5�Iy�u�&��f\��x�ШS����j:a�sR��F��Y3I���HR��-;�MV��H����9�R�E���pqZ���O4K%
C�cķ\\��?�N��&z�()�Z�Pv#ë�>�*q�����tv�%kPZX؏#������Z`��ް��ٲ`�c�ފ|߮��p���u#;'[�.�I�׭�<^��4��)���6��7�G�����1�d�����������ψ�I��0�j5:l���y����5�<V���0^�����J�ܷ����8E:}�\)5<ié��M��D�h���fLpSyICS��>B@��z�9ӕs�h�����<T]���y9#Ie�D�^NV6����y"r����k�����d��Z����'�\!<գ$psر,иQG��d�U)ZŘ��K�iy�LP^C.>��&U���QwgΙu&J}�
�ک.$߻c�^l۵��5bQuk�f��Wz��,ДI�P^Vj���
��!�b�f-w�g0�M&SRb̬����H�q��+��8d3C�X�8t�_��@�R��[��	C~��O��(�:c��˓���rZ0��5���iȘN����'��H*�Ձϝ��A����Ci�lM�ͷ��/�mȈ��H���#z��tP1��l�
]�،�;w�KPLҤ�w��VeJ��)�L>>ˣw�|�"�ӄ��Չ%���oT�Ui�d�/��QB��e�w���5���Y�
�����o��&AqJ�rvj�*rѩX4�R����B�Rj�t�
Y�:+G.��_z]ŝ,6�����)C@�7"��\��Ga������Pj�p*W��f��/���Q�ޱ��HMe�}RФ�b7� �Z�::ku�1�	��w��Y3q��[���OT�تП�;�n��O?����ac&���q�O=� 6l؊�����mS6�Jҍ�X�CZ9�0j���S���^V�=f���������`1�j�2�,��t:_���Ǟ�7z�ک�Ԋ�U;�o��V|��;X�]̀�"*_�� ��iS�ƛ�?�oS�uʮ�f�;\9�B���7��E^^�\�0���^w��V�8ih��{�`���<v�s�I��z�W�����lyn��T,��Ե����7��XfJ�gw��.�Gb�vH=y��Z�f��8k~�n������jm�1	d�.�y����@q�c�G��^\=�|��B-�Fn�@�I�A�^C��a�����6��r
20X�7]>G���k�aQԚS#��G����������ФY6'f���rT
`��M*J{DRE�T�2��w�uW�Z8�64�V)���#��5���>_��~l�"�� �I��]pŅ��aaɼ�_�����,��6�����=��T�U<�Ȃ*X
Nɺ?�h�7k:Z���5��5YW���\�;o��|i�󋔵kM�ɂ!�т���U�vJ,�Ӥq8�ՃʶF\p�T,[�j���diCV�ڲ�!9�so�NBA���J�d���~E#m͵x����_����N*�[��I��2}�dw�ъ�hB��.N�D��	�y*~�m5��?,̣��st���sJlt��W�/��w�G��hI���NY�����K����#�2��I����片Uq+�&ٳ�D�Z!��~�;z��Z��r��h�p�0��2��x<�M���71F2Z�v�]bd�4��w݂��{U���ҘΆ�hw'~���R+�!��#�d�>��:�lC?*$�atC��H=A?�w4"b�׬� ��@y�IU(
���V��&�D��r�$�%��Y."3�A����}�	���ט�ލj�̲�̼���hm�x��.�)i��d��L���_'�j�U�^�SNJ��JY��`e錽,�(��ZwwE>V3�h�9��o����ӣZ��a�
`�y�^M����C=*��i�Q�I:��k���+)7����h�)a�aLC+J�-��6���T�l`P�'�j�i'NBᾃؾ�F�"S��*1tB��-�p�9g��۶}�r���n��z��ϱ���q��r�6�Z:74��c�����h�� ���ĳ�Q��V��'n��J�{�m����i��f�:>�S;pM�,d��5�qeI�Ѹ_z�+�Du]������[䙇��1����V�$ߙ<�l⌧%\k�-�%ݗ^�'N�4� ��s��=w*����@����4l}�1���������������`��"N:?T��>p��F�=q8<��$!BcS�f�O9i�sk*���=�4���P)��A1��;j�Vj*�aQ�ՍX�����N�����J��l�jE�D�D	1�/��v��8d~Y����R�)Vu�Y���qp%��<��+H�<����<�ȃbI9��ObL�r �{N�r��㨡�$�:	��ܨ�[.1
f	ǈT��>h�K�������W����rnN�x����?�w=�B�6Q�P�CH�g�K���Rp��N¶�[����ϚqJ���0����Ŋ+��-/+Q�}oO+�u�X�v�ޯ�> ��G@ݡ=��V�_��'>�x:~徟v�{�0�\a�U���ގ�?Z(�%Kk��腹Y8���t�yB�Iw�6nU�Vާ��J� a�m�ȥ����
���GBx��G�� Q�'^��]�-N04~��{���Q$�v�x��׋�4�E9�g�r�z��íqL~�U��ԓ�b��x�A�9O<� �}�xr��3�2_�`ʄ�Ps�
%��1��ߵ'dd�bL�2Y�!DCL��#{���K=i�ݯb*���B�;���!	�"=~��}q����M<f�B��E8x/霋�%޺��k$�K��zFe���F��,EK̏{�}�H�)��O����R_��cW.Z�Q���w�w�4�4i� �4PB�(Α��P z�sL-c�� ��g�*�FPM�z��,ÎC59t(��ف����!�t�b��z�n<�ڇ�ER!	��{�A5��b,�e֭ߤ�\9\z�/+q-�p^L��]8���_�(���3�x�e�*�Er��q�Mw!E�9y���G`�k���+/Vuu��z�A���|U1c,�ުIǍ�ȷ�b^���Zk��3r(~��\"!� 9��з@PE�XG�b7��V��Z0`�0<�����p{�:�u�r����rQ���h�Kg�ܼS{����O?U��qT���p�w�q���ǎÇTD9bh��!̜9�7�?Q�eJR�-��$H̝_��������%pz�*o����x���^Y��<�y�eU�����g!�եM����9���<�	����n<���q,�O�����a�D]��U ��bwg3bu��0Q)�l�q�pԈ!�qXu�e���O��L�I[�;�����`���rh��Tt���6t��y5<P�Gc0����4�՛q��>�o�����G�4�,��;.��\|��@�W��#�a����G_���a�4��4r�s�)�g�b`?�X�J_����m�Ǣ��������c�@�xʨ�7�t�+�n��lm�޶iN�z"V�߬2t��S<��{�ۋw�(n����������_w�dI(��؈&N�W���`WX�2a1()�xl�~y���k��&0�$Fz��c��\�R>��n�v5�L��a�l[[����E:��,�=�x}
��_�\P"$�h"������B@�x8;�T�`ѷ?i��s�Y{�<��.3Ђf���eOWn�!�١�)�[!s�-�&h����F��i,_�^	��ܸ������!�R,뻩�"H�!����%�X��
���R%76+�()����n�QB�$�����#���W����a�X}��7�w^�v�2��r/�=z�������
ʑ��,��>�?IJ��y�&l޾K��|Esd����-[��O9YpD.}�x�*��"�
y��:ك������]ҜCRUS����˯c����t���d�R"*(��y&T���o�J�Mq�
oپC���~��^{VA���Mr�,���S�m� +�6:�Iy�o䳊���
	�����ko���n���_M\K�d�2ط�&��¹��Ő!�����Q��1CG(�g��5�#p=�Oc��Ԏ=UX�v��P�.j��d�1��ⳅ��-עGb�o���NA��ٹ����ݒ��U�1����a�4�M16/F��K��I[�ؓ?\��O�tH��8/i�Ͽ��J:?ϫ�:��9��T�X����>I<�\#^��Ҥ������K~��7\�ڡ왡ږ�cUO^����,¶z:p�J/y��������Z1t�J�)).Tfk��ĕCɶ�n�����Y�*Ct^�����f�Q��0W���`�j�-�Z��loC�_����(^ NjyPE�I�>xHø�����1T����̨gk�fL<#����he$�Ԥ2+6{%,rH(1��@�2O� d(f��uu�Q�s)�����סb��ګ�v�p<r�'3ݲ�~��q��ȳ�g��A�O^NVף��E�}���N�L0I�#gc�/�qŅ�$�
�ޥN�GuT's ����	��Z� gQLZ��GH�w�� ��z��u-���܄b	�����R�1C�W�}�5u ���r��n���o��'r�9��]��}��s���ei�0�22�;\]'!�`�D$�MYux���Q5L�i!�A�l�/��r�!��J�՜������AZ����eG�Nj��M�j���l	I�:�4��Z=n�}Y79�5r���p�C֦u����.,)�7?-UiL4�8L��d�����9�B�$�;2
��5��V1�#�<R�͙[,H�K�&c�zdk<e��6���v���)�0�*�j��7��"��F�鉥����	��t���0�9Q�^d��[[Q�-�\ⶔ�&!Y<�x�DO�Z��~C�Ӫ5�VLJ[O�5Ǻ���k����1s�X�8F��N��^��08c"��3���I�IVq^j�=��n�6v`dE씍OIH�c�"I�#���};��¸Řx4y�KFoߓ��[ۆ�����$�P�.t��7�ԲVAY6�OY�J�aa�������i4�r�9�&�d-��8%0���r9,��R�\��\��L\Uߨ��P�U�j�-f�+
0s���}D>��u��|S�'R�m�9L��.F6(�Gg���tE:$���O���^B���]s+�,ִ�'C�f7�s}�-��9�*�э�-�F�P�H���oKѧ$m݂p���lOwhHۛ�քZ��G.W\�8�G�l�NY��cby��R���tK���9*ۋ�r�j�&��v����	ՙ�T������7�P�$��.�L��/��Q�]��$����+���7+@�Q�"9�r��,�CaAQF^�3$gJT��[9�,�[�y��FL�Ix�+	��j�+�O��O��C��I9C.�G���~d�I,n��Y�(+/�Q,g������dZ�361$F���3��,˴�DR�f� /&˗��1YX����S ?Ò9U�<���^�_���t�r��W]�i��-r��i��Ծ�A�ٖ9�iٸ�\xՒ !Fb� �><e7�ZF�9)2�e䩳���MXgN۵��\x�,7�
�n*t>e0R4�jsj�Ϡ�~��ߣ���խ$3&��)B��x�b464����i~�P��iِ# a
�͎l�
��DM"Lήln�+���Qr������{d��r@��{]�S���
�	��J�q�]�	���)�ʥ:�����x�J�%D~�m0s
r�Ag��ѓYV�9���P��B�\Ҹ��`�9iH���5�ݿម�ys�:S%�aR���W�\'��nS}�ʲ��8KWP.�]�}�:��Ì�s�h��Z*���U��b�Y�z�t�*0Q����t�����[�l�����}-{�@��,�� �dmxn8R�)6!F�i3��9c��/�!_�5�+^�LYG���*��e��Ǹ�&N¶�0sz�x�6ٻ�#��zz$M#��j^^~|Vc��������Nr��8O[����P'����Wtj��+(q�� 'M��F9�џ���A^a�l���]ݸ�;������Pr|�b Â���3�����Zu܀�!N�#���$��R	�Jrd�����nS��<��֜J� 0�ɩ�L$f�m!b�?���F���۪�(+��\�#&�ݭ9Ȗ=	�w�Yd����ȧ�>���[^�a�e���������X�Zc��`���`���"Z���Ĥ�1j�:�5%��ԧe.u�byi�G��PT�@-��D,�x�%��8�E���9C������e�Ś]�䒉WJb��-(a���1N���0AC�̘T��.�6���W�!�ć=��6L,�xF���
���R)��9~�'G;
+��@A^�x��\�|-��΍?�h-��MrU�ٻ�8�R���c���m�UȞr��v�Db�G=\.B�&�(��d{"Sg�ODޡ�������M����Nx����'*�LA��N|�d�W˭d�Q0�[�&�ҒbDĻ3e�>�÷�q�0v,��'�/���,�:���G�x�����8�y!J��Ng�Ҩ�[�q[y��F��X�Ғ��3V�B�%��+�j�#��5;��Rc�@qSg�~*���7ݺ���8/�X"�����k��WK�X;���2����&J�JvcBB@6lZ"HT�@���D9���V\r�y�n�o�PGZQ�'�p������ {`B[0��#;��˨�P-�M��U���۟|#!�Wٴ�xH�P!�C�H,�� [2����օ������Ę1������s����Ӌ�瞍�\1X�Z�m�W�:�ɨ�qT��ǏG宭���K����w�˧�tXbx趛��@k@��%rv9�:Gg(�GSGA,�%���[*��	��KB'���X����P\X�]�M�uhD����w���C��������O�UAed�-�������n�@4�\v���\��8m�N�g�g2m(�LW��$Ba�'�AX�N��	�H6����6�ڕ+T4�����n%&i��\���N�u��_P �1k6���R�A���"�:�t��������CoN	5Ə�C�v(/;��ضc;,���Yv�G�b�s�5�	�7��Fc[J��CT�Kw&����w�|#^{��V��"ݸ|΅rPC�RO����rւDrK�9|�p4�a���9�d�*�K�̘�_�}&EI奎���ă�/E%�v����lD6�s�EMm#=Dyi�y�K�p����{��@���W�C�-��\��-E�<:��<v?�Ǔ(�q(A�.�~�)���0[[�yȪj�PZ1Pcl�޷���L?m�x���?�^�S؃�N�8S�S+��=��z!�R�k���8m�	
���Y�{�^�~��-[��N��/=�P���ʺu��)eeI�4�a�6;|�V���V|��|t��c���J�#�p7p`��R�ݘ�G�	M>��<r�mؽ��%e���͢o�B0Q.���q`��[T�ş~���R���UU׌�ݕ8q�͛������Y`��Y�y�Z����bÎ���Ǆ8sXNAx���{'*��������'a��5zV'L<NP��ފP8�������-�3<X]�%K�c����m�����O�/C[{L�Й5�(�ܭ��BAo��kNm0%�:����3�=�8ڛ�p��S���^�v+z��(N�!����H����j�6A�6i马<��6c��#1j� ��/?�!9G}����ET��~�����ހ����x%���BbQP��|���'�;��%�F���c�r�U�?|�&���Oæm���;0��)h:���ƞ<|��smb���ixA!�?׬��6E[�Ǐ᠜�x��7tVŬs���I�i�JM��A�Wu@�B�5Kcw������x����9�tIH��oh��]�@{��{�}���b0�uq�8���Ko���.��{=]5x�����UJ��/�N�3F�����/T�*�٨���
n޺%�$'����t:]T�GEa>v�ڎP(��bźM8P߄��C�W"��<�׋�5�^��}p�UנCP��:9\+Q���2?M��e�n�g�s/)�r�o0��倷c�o?�_O<(��Y�4(9�w�VY��b���z1����g��#<��~Y�%�}�6�i�0�(T��p��q`�A�'��KQ�S�e��I��W�~��~+B54T�U9�a9+��.���e����E���/!R��{����y�\4�9�K
a�pۥ�Q�*s��� :V���v��n�6�9�"O�2gÍ{�x>t��gY�@.:e�8���T���^�G��`?��U��#�)�H��f��@9
�!R{7^4CB�b	C�8XY���=��~\�R�b�N T}O�)�	z��s/��{n��d/{#A��_y]�50��g�����'�EQq-9�c���R
��0�̩wTㄣ�� ,jX�ki�Q�A*w[(l��e2����0-*�-���)�޺�G��o�Xm#�	v��j���nډ���樀�93T�:9��,E��t�Eb��q�9S%��iu5�4�8�� ֪m�0��)b����=��߮r���?�O4H��)��E6�Kb���45F�^9�����w�[#nV�ą_+.S,��א.�:4�LL��/�0k���g~%=~����ك�6jB&(���?��x�Yz�0�r6�����p�M�kY�I�f�!p*���������ͧ_遰X���J�).��?-�ygL�IS��lT]���J�vR���e�`sy�3Igx���ظ�N>Q��U�L�֨ү;�S�E�}��m��oU	?�6v�a�ت����C�N��=��-{�X���gê���o���6�ҙNO	
�r���3ȓ����7���J������_�+k�}%��l��x�b���i	N�<[7lPM����5ʜ��ѯKR�M&n٠�Q宄檼�Ͼ�n��*�����u4�aANEepe�$�ۢ� vO�,���:�C���${�T`�ϋCRvg#�a��%e��.�ҟ?Ei����jژ ���A#�W�č�9,��g#�r�ٚ`G��^S1c~��h��=f�X��q��3�#h�8߇=mZ'b�m� �%˖���Ię�e�p�'A����ǟ�7��>%��zMr�zUP)�0��t��^BQ�
c�.K�6Cݞ���l��D��0�;�	+l�j��`v*y1���A�LV�`Z�	#���Ur�}}�≗���[�*׆�I)tBu�5k6a��oT�3��	k�7�z�	�?Y�%�rnG�R�m��_����(��X�6L�d�WvL�Q���/�D��a�0d����o<�1�$�|���8o�ɚ�hj +ǭ�.7����<Ur+(>�>}ɔUgp�V��ⴓ�G�>�����w��T֛��A6�XKZzaa�^P�5B���?��k/��Π>_��)q�M�����ԼTћ��	ɶ|� L�zrm�Ab7N@�q��Y�ה#F��y�w?�E6�,�ɪ����z8)��{�L�;3�+�# ����(�����g�DcIԘ��Kb�1j�wĂ *E����e{ߙ����>�$��K>FEv�y���s�Q��1{�D>nټ���bhe&IXG
��x(G(��?H�)���Z<��砐jb������y�0턩ڹ!ݟ5g��?�p(����˺*�SyI,V���q���hK�^�c$"yu�2����)��$B*�$�2%���;��˂��+܅�۶I>��)=?�Ȫ�}�p敇@;p46����HC@Ⴒ
���b8 j�X�H��;ҰCR�0��^U��m���֞8?ae�صo?��Q#�rm�~kg���'��Y�b��QCH����$8�V�gJɺ�7>�T�X��Pt�;OK��%�(�8���Y:�E�p��(Ē��WR��?^�	c�k��׈�\�ۏ�uߡ5,鬜c�Xa\�YRd�4��R�����(-*�HϪlw��p�\hjkG�D,ܲu�b<As��'�y�7��ś��.)��ƙM��+b����:�Lb,v�A�͆ 5`x�I9�6�����)uXV��EJ�����g�u�I)����%w�믽-iP��&mJD�p�_�2X\
뫟|�GIn�R�A�gaI������ȧA~�1�2������0a#�@���e���0t�e�m����d.�����Eda�2fS�R�Ei!���J���ޒ5
t�8m7�1�~�}��8#CH,i������4�3|تd(F������'�[���;p3i����5��|��~N�j����N��D�\�/���h�C���u#H�"�i��c�86ٷ�
ʲI��VVZ~�#����VÁ�1!�&X�Q]6�+�`F�"^R(PI.�OR�Z��v��?c��B�)h�/��cю)gV��f-�Z�,'�P{4u共��~\<!��<��P�����=�r`��Պ'f֞��P��Q�F<�:��ˏ��j���,ϰ��{�Z��&�
#\��$�h��� ㈉�4��d��"��yq{�$�g�2Y6.6#��xy'��|o�M�89�4��ܮ|/��h��S����v��,t�T.]W�l5��5k�A5C�٤wq�*��GbJ-�͢�C�Wt�=���Z=��r
Y`��L��A9�Ë��D��a|�[e;�֤!Ea,5 ��ְU�M��A 1YBo���;3���v?%6t�����s�
�1��T�D	�H��ʪ�K&%N�T>m�(�R��j�~�!���0p��*�k0o���z`�r�|i��l>����7 �?�d��ť/EB/^���0�N%洝ʶ-�M�-i-ܙ]�����u�?��횖8��c�p��~��N7���e9���<;���p����s�tW|=�棪��Q�V�%��x%gM+�� 9�~]Jgt�&}���u�����oqO�bєˏ�A�;tnМ��g�s�-Ns��Ý��Z�������J����0�bU���V�^Ze�f��)�gp���m��bh],����K�\?	�I��2y�<H�xG�!FmQv.?�1|��/9�o��zES^�&g�G��)i�І���if�Q>���A����� ��#�+B>�!A1-��9�r�d6�pv?� g|e:=�Ԇ�?�r9T�Qq��l���͏��`��հ�4��0����p"� ERW(����[��9�w�ԝ�<l-'��.�괰@n�e�"Z��G<�"���6e��K%� L��1��nȮ^��)Q��$?���0����":|8�U�KsK��4�z�p3х�g���L��#Z=76��Hq�M:J��G&YeF���o��3�ꆖ�~�<5Y�� [a���@�	%B���d�!�GRɆ�%�rY��lGR��8�qis�Wg6��ğd�\#�5Iw��D�<%1,D��1�4y��3~�bJ+�C�b��gTT'����4]G�Q��\��N|�X(�����%X����%�卶^BF9�</�2+�/;y))(��N܋� ��s�F �sYܖZ�#�DY�jvD�J�H$1��g�Y�L�j~��^@:r_�����LkK��8"�ߔg��%�s��_~�4P��,����#aQ"F���p�B�g�l���<y�I3y#�`�����@^F�<_T�+��.��x#e��OvK7R��J�|�M'L�q↘VJ��##X���4�u㺛�d:&��ӱ����ҘBu;�g�vZ4��y1pc/���N#&�j�GaQ�|�sn��4lb'-��dD4:��Ϊa�ԧ۬Lf�nx��$�m�T�ZSjXN�2'&��B̜q`h�KMf佳E�C\g�h8��`�W����E	��*��^6#�sy�'�>���_������<=�,t��C6��?��?��"J]g�g#����T���|VI0�P��;Hxb���[�,Ť�L"���zr��-�RT�!br��#Z�Oe�yDL���E��.T3ĺTVT"�Պ�#�bˮݰ{|*@:9F>z��)\6G_��3ZE�|Z�`ջ�H���
��慟uh�I�(��-�|���#�y�¤��u+�_�`Ii���HM��Q
���AIc�J*����H�F�yv��W�3	�y����ސ\+f#`a5�Ӆ9�f�N/ɪbm�m��P�HO ޟ@B����1R�~D#!�}Ʃ�rJ6c�|��K���%���+ɳ����H6S%$�)\���sϻ��!�iα oǚu�v�f��J%�i��d�<+cj�aN;d�8��DTŴut��_��7 D��;ЬZ﬊��vuコ����#�􄵍�p/<�s�6�ǒ�_�:�jtC��%�.F!�w7�ر�p��KQD�pv�x�39��湣�x��UqQi�����ɳ�}�(�蝳'�Ҵ�!w�V�ӅK�Le霣���;1դ�����Y�щu�j����������i��+�5��KԱ�w?�P!�<��������X�2%z��r�U�����J*�ɪ����f|��{�"��M��<�w=͸�+�[��),R���^{SuM3��d���[y2%�9f�0�<m*���i=�jU��%K�B}C���ޣ�'��zwzX��̚9ՠ̦�c�7V���p
|�)Jĺj�9U���=ND.�M�_��X����4c���'��!����VN��P�Ks�_�M{K.��l�=�u�������S����׬����4�>p΀�ɢ`�mM8q�$TH�O&nb�zCY��c~��x����	����~���7�I����O?��P���˪2L>a^y��t$Q�ѡ�ˤ�Z5ec�l=�;o]���Úy�ȹ-Zg�4f$�e?7nۭN�j7M��tw���e�\��M'��#������p�-���?�&ܒS3�P�ʜA�K��].J��2̙9]�tXH�85�b��{:0}��(`�{�:�]�RFUޜ�������֛oD��K���*�Z���n;~���Ϣb�@�Ө�I�x��=c�n��&�14Kd˖?V*�fL7�A7���B
�Ęyt
ZSl��X$�I#�q�)�U�,���"I)��+�����=���1�@�4�%E{������t���~q��HX��D�N9f������:�kv����:r���܀A先�7�-�8��[ֲ��]�G�t�m�N�xX���Ţ��,�m��������*�[l�[y�����J�[���C(�����&T1k�T1+a�CC�yN[�%7�a��萿�Mn#�&؊� Sy�[n�
/��>rv�x��*�HƜ�˪J�p��c�jFW(�"��EE��%�����U8��&ʕB�$�q*�P�g��Z�jզYסāU<�֞>�����g���2�(G$����ܐ민L	P�}r �-���������.<����/�Ԩ��|6+�ڲh�;������ B��Ȓ�|�}�]������R���Vƪ^R��k��8e�q�./U�ޖ�.TTU���R�������Z����*4b�FSr��B:��M@T�(���a+����MM��[p�=��cƫ�m���!t�6�r��m�*�αhl��}�B�m$��C?v���ҮXI���O�~����w߾ �p�N���~JK�-�Z���A������QU�"�tbx9�9�Љ�ϝ�D��m=(��Ҵ�,��#����!U�Ȟ0�ފ��.��(��%���ooґ�L�Ee��vt隧$�h��|����މ�F�8��Dd�>o�lI�%��,�X�/Qb���]��#�{�ܫ7��Nq���dĜ����0�٧��s��X��klܸA�x�5עB���z�G���O5�-�u�ii��݋��N����>^�]�(+
���g��:�R��Yx��O�4 �@Wg+�r�8����9�%ؾ�6lP�̈���;�;l��6�$i��.FV.N\"�_^->����R��5K?g��P�ؠ�U�%bP��\RV�V�}N/4 �w����|�E<������و�z8�	�����-,�q��
İ��w�uW��o}$^�%���1�)ǙB�6DuE�zqx�N�n}Ƥ�G���o[�E��,�v�ԂC��/���\B�؇�����8=Y�8n񢭸�����K5̴��ڨx����B.�A:DftB|l�E��Ue��8px�!�{�]x��t����v���`ώm4�Z��@~�q�\�V��8m�<����U�S�h��x���Q�"	��z������+t�Q�2q�>D�p�����e�'�H#��\"�1�G��7K���NO����DEu�kCk�<��#��������Ñnd�=�����R��(X,c�����r�
%��*b��SQV����
L#)[]��"P^����J�Ԫ�����hlm�{/�&1�4L�9[kGMG��{~����2�>�^�z�ǎ��IJ؉��X��J���{0p�v�.�3U;&�5�I���umF�^.B[k��t���� �F����{-�yCV�%9�������"�ٵ/��I<�ؓ�i�����3���cG�����ո�����C�I�8d;N<�X�;{�¾+lN�2�D�ݲGg�L�����Ηu�(��7���h����~�_��Sq��}{ϝ�ş�xZ������}�4�ߎ!#����k��?n5ā���ʹ�˥'w��S�b�n� ��a�5g|b�̲�k�m�S��K��a����?j����נ��֮P}��;�J�2y�0�=�$��i��w�yx�����N�K�7_4�\db����[��F��a�Di]Ī� ��w�,�B�
xq�lD}K��(I8�����vk'k-�Ko/A}}�Z�>���#�YS�U���S��x���(.��|�3���X�Ғj,�v~ؼQ1&*�l5��3fa�ȡr�{qͅ3���_���L���r�/kk�FU������e۳�Q"�x�N9u�J�	c��\��� '���9g�	�X��F>|�n��b͚��1b�hL�r<J�vq�m�������ZM��N<����5��/���
�M��=M�㲹硾�g�2[6?�D+T�?h�F%��j<�қ��A���W����=c���]�z1����9(��x��e:�%Q�~���"��x ����{�~���i����뷉�q"jM!�t(c�\������6m�-�Ƙ�8Ңo���+.�����b�w�=��)9�Nj����h�cgc����e,���9q�п1��+;c:L�����.dű����qvbin���b��%]q�n��$�|�/p�g�H	1�f�����2�~��^ɥ�$�vW��.�Q�E9\i�oQ>������%�;�W.R%�F�˨؞���UC��/�]�Bq@�A�:�>q���R�񣪕d���a����G��A��(OG՘��G�����>�u6��-�s�,Ƹ�O�{�z������E�nGV"&��������FŠrXb!޵�5e�}��iŠ�BP���/Vn��%'��;n��c9�"~����T*����H ���~\�sfO�����*�*�����c�W�AI'Μ!�R�C=��_���9W:gtY�lކի�ko��d�!IرH����^��p�z/���D�2/��*.��_
�����>C]"
�Z���W�U2��$/S]��ZB�t&�m���NlܺS�jH;��`Nr�e߬�qcFk��)!';©<K)��<
m���<\'ZG�D()�<�X��j��E�z�$���'dU�h��Q�h��3"�w���u��������޺]#�sN�f��;\N�l[;����忽�٧h�l�ص�Di�HȄ͛6c��!����Zb�f�J�"ؼe��}}�Fo,6�4���J}��L35E��I����K�w�ۓ:[�)��vP�˰R"R�9R6xX��ẙ9 )G��%��whv�ާ^���]hn鄣����bDM�:��匶)ź�ZC���c������R����M����ч�ӝ�Bg�y X�M'�R����pL	�n?��5�%�������W����ԡ��R(H$�Ө�,�>���;z��Y�9ؿ����S��O:Q��I�LZ>�y!��[��?��=I�%ُXo�hr8.PZ����x�b���ڍ�R�3�_^|%CP����rz{B�1RU��")�QC$up�0�O93��$�8[^xK) 9���a"mC{wX�k6o�c.8_"�>Y?�ѹR�ʸܩ
�6�c�dD���MĪ�ѽ�$���1r�@X�&�6(�b�y�d�J	���QxF[��������mª5�����)��^d�޵���*&�1�(��ϋL�u���r�LN	��q�n%�~ĒI�-��/^�<�ȟ5g%���"0��Ĕ��T��ڲ�	�].�Y.����Ah;w��J�@�hD�G�P٥	J��n�0�<��DYA�l���K�a����NPp��mW[N�R��nI+X��f�P�jb6X�'e+?k�\��权H�CgT'����')yW�4)���v�2(�Pk4gEo�����)k�/ta�#b XP�P�1z�n�Bt2��b���{8r��&�%a���`;4�W#sT%�kj���@��إl�}��ǩJ���P��gt��
�ab��Z��p�,�F6I��r�6oف�F�6[{�� y���j�
uh����¦�>�w��IQ(^��c���<�H��r�ڝv%�ټk���Xe�ZU�f�)> �R�I��)Q&�I�#3j,H��(�i^4e�	hZ��f���[��Tٯ5�5M�Rz(�p�HҦ�!Ma�+>���^y.㙞8�]±%d�:�U��@ޗ-]�K�C5�4֚�l%L�g��>uB|_�ɘ�n�;�s2dC#	8�/ȑ#F�d�?寜�g%�8�V��ДG	�����!���/�/���d�,gr�����@E5�9�9�5)اCe�ތ��]�v�<�@�����Ѫ1��v3
%l���TpGǴ-�H�t�"	+�$���fٌ\�K��jC��J�GȖ�c���q���S�$�����x�K1$Y	�X �3
�?���)���4���Y�X��F7�j�?ȸDak��#�Щki��_����T���mf�*��>�ţ�65 !�!�A�6��H^������N��a1��l�ҁ>��h2�$�;)����&!i�~~2O.d��a�M[�*|��$�����#I��x�2�E$.�cʐ�c�.��Fr{�x$�X��7�^��!0#{$B�[�)9\.��]����ĳ�$��m:���'�=r�rP9����;��[��1�[֜vf�����#fS^F(�#tL-������I�%Qe�,����N��[e?�:L��gדHMӔF�����#�'�3�
�nubH�5P�YF�tfiv3Z@&R�Y�B���d������c����!8;��X`m�:(Shu)]���&`�DW=���������%e%*}��ݭ]8���u�I�BKr��b��J�3�d�Lr���DsN��݋�SO�w�V	�.б ���yd����1c`n�3hRa�e�J�րyW͓��P��x,g�uPiNֶ��G�x���P׷�>
�%�Ѱ:jF�'�4M�-E��S�ј!��޽[¼��8d�����l
��u��{����a��i�u)K��b���hi�'�� =�=�'�OJ����5TWWjxkYZR�d�*�l3�#��D24ZY�"�R�ٱk�^�<i�oXD�w�]r�s����s��O,�������IQ�,|��V�Pr�Q��-�Ɣ�'�˯�꡴X$�K, �=�HIh�S~�"2�3m�Js���芡D�1!���aÑ�k��H+��#ZB��m����s�~UD�G��(��R����㤘V�-�{0l�0��'�=��j�[��QVY����̝�g_~[ۥė������C�*��
g��90ж���ET%Gp1
\^�\4�L+9^?hP�NsN%�2p����[�P�E�uu���݈�|f��%�qț�S^������=uRh�m&C'�3�!0�9j�v��}���u�|�`1���K��\А�e\��D�H���1n�$�/G@�9a�L"	쯾�"Uw��f)U1�{�2d1��ݳ�^2���Pѵt�,�Ǧ@����"�R�(�_�v��o���O�W�� �H��6<����_s���Й�P��!�Hy)&%)�عfn�헸����-*�@�_w�!�w�o�A?����.���)�38��Q$F���.8���c��Ȋ�I3&OFP�3��$eN&2z�h�؆^��g-��0�D|��Z�$����Kl��hcq�ǌ�T��ɋɏ�5T�lb}S�1T�T���}(�M�F%/T�I��G���-��Ͼ���T3#�_y�֨	X�z�Hd)1hVY�T�Os��\�H��'M����d1%4�t�I·�<���w�&�=��.�7�=qz}jn0�0��0$�G��.QBZ��(�C��9瞡Pr�U&����~I���0qĜ�z�L8��ǎ��C-��dM���͖�����HO7�%e���(*R$�a����O,�M����]�?��im�hok����~��[6�hP[wL7��&��ݏy�ߛ$}H���s��¯Vja��B�3�W��;���S`Z��$am�W"���V1�.�:�X�ݴIR1���$l��]����]*)I�#�ˈ�\�a�d�e�{&�}�
?1-~%��ȅ;���qx�nY//vl߮��J��zv�{����X�)�ʪM[e=p��rM��样�SAUeg-�߯�vrߺ{��<��S��曮�{o���K!���z�(��ԓ&���|b$�Ӻ���3�y�N�z�8�k'�^�x��Oi�o�t�Z|�߀P�Drr	�*�;�G�abH���w6�Yp�-z�������!)E�8�J���u�����b&�J8E���K$���8m�����O������X��F^���ąg]�<�-,��g��#�� ��K>ۻ�"�X��=;��wbѲ�ؽ;���G��S���F+����+q��jm��������1��<�{,�r���X+�3s=]	��g�W�����\�Z84_,[�l��{�ᑇ�ƒϿ�7_.U�9M��9�#*�!�u��"lؼ����T'a�N<��ho8�Z!k��T��g�����p�3� ���o��}�SkS�L���OŖ�?H�W.���J�\�I0��I$�z��X9x!L�q"�N:�>���U�>^|�)l[�zN�z��lD���d�Pb�$���e8k�Ltv��_݀�[b��KH=��_�H��Mk�k��7������x5������Xp��ȈQ������ɋm��k�ͷ\�hc�b$���k�>8K44���65@>Ijw����xo|�	֯ۀ1�5/>�8�wƌ���$K��7O8��	?7lچ�ۊ22��<x�/��_@�v�<e����p� 
%�{��W���+�%&�Ǟx��q�J9L7W̿�v�Q������g�	�_R�/���k'H���o����?�k�aȠ!�ͯ��K���<'����?c6�/zWR�F5��KB�^\.�_LK/��OD��`ǎ��/�kkw�"�a����5+�3`��7�BQU)���#݁�������w�D��3�狖�Q;}�t�۶A��v*�⥗^R'�e��K��=x����d����܈��}���q�r�>m�/�r9��v�)�O|_4cBa�0����x���	�i���#�j�*XT"�s�b�|���x��Q5p�F_������.I���2~B��;k2n��j=;��N4<dP��g��9����Z�(.+�#�>��=�4��h��NR�cΐԍq,�XX5a�eX�a3l�4I�C	O����o���|�,�]�cj��8�Ș��xPk�F���b,��V�WT�;��B:J���]���M�0yT.=�qI�b8T[���נj� T�/fNƼ�OEw����S�E��!�X��`��($% ��T}ۂ��,\�����a�<�ۛ����k�6���	o�
i[������(�YZY�g��&������|��߮�˭X��K��A���X��ke���/�S��O���߮ڂ����ڄBIM�x��o��[\Wy��_��hJU�
K*ݝG���.�o���v�øp�#����������J��.�a����(E��ԑ���ɻ}�~y-�=�ض�;SZ�y�ގ��Q�k��34u%�ޢe(/���ǚRԜم-���8���F!%޸���q����OS̎��PX5O>�2�%5�hM��� � �W>\��f�*���XӇnI�w�U��v��q3"��y�Or�0�sJ����ʹ�b��oQ]^��dOXK"��o>׶𪍵����v����%���'n�w[w�A�%�_�Ʈ��Uw�qLR��?�Eb�r���Cgt\�,�7����v�`Ň  ��h��Ok4��z�Ӆ��%:w⠠�)i�2�",Y�	�D1���z�RI#z$�������s�v�Y�A��΂u~l�fb���#��Ko��Ii�j7oR�a��-:��_��[���oP>h�1�Is�19<�,��m;��������\�O,;��q1r�1�NXt��57���T�Ϣd�0�q���(Ö��e$��D<N��n��K�ǞTF�F]�c����P?&��N����c���E�H
l�(�!w��GGP�R<�Û�HB�X�'Ń�⁇���O?���Мݭq�-|H��G����=�M
lٴy+
��%�M`{�^�ܵ����>ߪ���rk�hŢ/�Ĝ3f��F8��Ӧ��$?	K�������׍a#�'�`i-�T�ں��Q��
����y�x罏To��Ѧ�x���V6��������u���qV���je�ZZ�ڎU��y�G���_yW_}%�H���S�mZ$�(--��"���0�uv
���)y剪�+����B�*r&��ؿ���3�#�����#Ym��M��Y��ߩẺ:����p�'����ۻt�"΢��O?�/-
�O��?8�.,r����ӧ!�(���Ĝ��(lرF;�'ԁ�|M$�Ӿ�S��K�����չ��GZ�~��Յ�b?ꚱw�A�#�#k~�'4�ۋ�ڜ|�D���+�� ݟx��?o���w����P�7|+<
좰nUYS��/�9��ɔ�B�������>��>:)�?���+�c�.E��v�)!���H*{_"�����-;d�0�^F����U 9�˯���.8��=�}�v��.445b鲕(���r]$�&=�%���=Y�Ï�t�xL;a�*���]{���{�X���56�����?|��F0d0^z�u\w�E��
����������ŗ��Ҋ
�W�XW�����$][��f�I�z�P�D6��u!�܊ϗ|���O��o���с7e�!ՁD����^\v�\��[Q"�I'h_݆߭���c�o�K�Uyk/V��Il���%3F���"a�޺zԿ)!�����>��T��]�mI�Ɨ⌙����&�(Ʌ->,��[����EkniĖ�_ig���T� NQ��1䴏o���k�x:��d�[r�A,4Q�]=a���oT���v��?�����#�KW�R�mm߫����Ҕ,��<��x٪�3<�	>[�-܄}�汚�K)1�$�a��u�âB&EW�n:�J^�?ˡ���O�C@� �U�0�����_����(��d���d���㳲mi��0���1mL�%�<Ex�aqM���T#���P"3��&����R˖ED��t�E�D�l����u	�����W�v.�S���eF;Q��tH����UZ��lM@�vm��������o4�eZ�y��m��PFwNeӣ�$|�I(�3Jew-��T�����3k�ʽ�H����}}��N��_>�-��AJ֬<^��P�g�kh�ԏƊ�[����R�f���4G�]�F�_:�=A}1�o��j��y-&k�#Ƈ@I����(�0m���4C��doZ:�x��OĪ5��ma�>s6H-sIՂU��\F�ſ�QIu>S�|�Ӥ��ΏW��[�^1�7ʋ���JGaeQ8�e�X��`�e�ֱh�c�����tjW���U�K��`N�mSZ�z���O7�� xLذ��I��083l�B�8Vᕞ.?�3�%�e�,V&��`����e7)B������^�߲Ӑp#㲩��R�TA��,�+��X	IHA�qq�N�z��
ꐵ�U7%R)��&8��A��@�a lY�>��w�]�d��@rZ�����#�S��ޤ\(c����D^0Xq��LfN�6AI���6��PK���!AF��*ؔ1Ɯ-]_�C8;CT�+��`d$�N&�����sd�F1��hReRVyIB�$���Y�Y�� �2f) DHS��g'�b]�8��p���� pɿs��'.�%uO2��:���hҎZ:k�2bNzR*aɝ�^ïW�d���pjN//Q"O�䔴�F�4X��J	}m��=�;A�u�(1�A����$ɗr&�7 N(XZ�sD�]B���u&�P�@?�C?��Q#H�8Y?�U�̥�)�H{ҢR�^��( ��󯐐J�G��0ރ�`�S/�R;���G.~��/��4��UΓ��4��+̤��j��j��'!���eӃ�Ōʥ�x9�5F����ݔ�E�I��H��j�/�ae�\d��?��v�1՘'���L��F3Ҳ�y!8�OC���'�BeH�M$����	��Y������*3VF;5��5¨Ԟ7|�F�����h8�3X���/Q4�P#�&�ُ2Y��)�1�T�(K��<!�ri�r���`j��"g�!:��qG�?b&��u;�D�O�,K~�m�kY}&�N)�*Ő�4�����f#/��gԘ�w f�DDcK�>��nӴ�5$��ږ�ᯠ��Y�<ˆA$��<��DP�3F��L�����l��!"X�]���(C�rj\-y"���>�X���ESVs
�gtz��1��g�9�ݟ�j��(� ���h���f�l����Y��X�"@������b���A�+��#�����_��fP5�sG�����f��p��<o�_���RDRsHS�!J?���ܨ&��辊1�8�11*���p�+�7ќ�@EI�HL� S2�팴Fɍ��O�<�C�]��vBy�@ �hN�9ְ��.�$3��"�H�O��.��P~�i����%傑Xь9�V�*�K��L)MZqΩ�7x9�A�M*w�b����{�I��մD��:}��S����`�D4���nW�>�&Ǆ�BI����Z��MQ� ǜT*?���cz����S��`/S��W�=GiѱjZ��v��,k�P�V>_�׈�Rj���X4*�G���]��� ��o�vv����$ �hOI�K�G~���� �}�L���Y.`:e\|�~��9-�-���}�(//3�ih�G>���r	��k��5��p�h ?/���A�X5X�)�ŉ��k��t�L��t�u-n���nuX����"w&S2vG�q�+*�2Љ�t���Q�^�,b=��yʅ���(�7އ5k7]#���2���sU͍��q҉�{]z^�%$g�M枽��.)�H'N�i$McA�Etkwgj*+p�g��ڴej�R �m��h��o����(.9��O���#��a����� %�՚Ndr��90�G�&~��sf��cǎ�5�:�zH �ҫ��1"Y4�WRZ���s
�Ů��E��.,�v�"'�D��:"q��	�-Y�W�C�0�C�f���$���_�g(8z�����BJ�����3g`��pZ���G��%�Vb�m�4X>;k�W�ܜ0i�{�ܱCbډ���T+k1;T�8"���-TY: �!��آ�!=�����m7!KꅏDz��gQU= Ͽ��d��_D�ߴXO+���r��'y�]),�QVQ��?�Î=��#g�v=Hq)t��@[s~5�
��
���"#פ��v٨7(/W��e�y��C��/�������Uo��7�D.�c��~9(�d&�j:�xq�8!��̙s�g�N��>|���*+�j�F�۹_9-�+ק�����Aq��gjg�������f�4Ͽ���x�,Y0X��#���9����REp��6u"$�!�ū�(iG!z%}����U"��)�bG��)ǩ�!��E��ҦK/<O���������?��w߁���(�0VJ���#�Ř2�8��A���r&�h� �!AOW;��Vy�B�r'X�L�Ӕ�b�~���E�NT�F�F�$���c1�iH���t#�P3��Ϟ#��+�EQ�!����蝿��G�����|
��zymqy5<J�o�<����Gծ������:�Gn*�xͥ7|��47�f���vܹ����c��Y���ڔ�O��Q�#7��n����L�[�h7���_�m�8�I�8@����!��-�4���D:ԍ眊���LG�sy�;�~�4�M��qռ�őO��N;@b[��&����@sG��^�Uq����%EuY 'O���z�e苳6��ה�t��o���>�
)
y*�ln��d�����u7�G��I��ٔ\L��]�j>�k����B�|�ߋ��Q�� \GK��
�u����J����&�Zq�)P#�>�ƦV-8�R�<@M�!{)Y�s��P��H�G�'7��
��:��������3��pl_���Z�b`��衃�p2���6]#�<�ʦ?���q��CA�R�,�d�"ϣ�)��
�iL�4R��>�K�ǎ���mM�;x �%^�}b��Y���Y�]x�H��{~�`QY��(a�̈́���z<�� i10A�(��`�}�x֢I�$��<90x%Y+E�7]u9�x�5���R�gvGV5O�r�%"�4a�[�%=���?����eC��0������{�z� �?k3R�\2�������l��u�����)C���D{G;~u�\���W%���:�vd�ψ����q��qDAsCF�U����u��*�3�4�+瞍�߭����S���ttBN�\�̙y��m2.��z��JUԙ�g�4	��~"�x�E��S$nNj��Cmu���?A��	>�C�	�p��
u�*�e8��g��ڋ����D�=�	%*�JJ4�p�_|:�N�ֆ�g+�����[� �Do�]H��x��?�;�E�Y���1~�=�řyā�����@��'{�	܄R�:0v�h�W'ʊ�� JR�E>�ah�xN�u½}��ګ��[��f�d�ȃJO��U�l^�����>��[�+J�.��SNR����N� �#�b�K��y睇��Ò~��m��#�"&�%y uZ/<�l,����Sǁ>���	��[o�Ӥ[��L.NRޥG�IR��B�͸p�,]�Va���2jHK�G�ނ_]+���/X��pTCsrK����	f��0m�d�۰	{7+�=#��!�݉Y'M�p�R������(����*T�����
/��F`�DZӄ��9��Sz�7���@g?v�܍B���%����;��~{'^{�cĨ�(Ǝ\L勉r�E砷�.O��?ٵ�ho��VeB����N1~��þ�f�� ��B��=CL����rH��Kp��^[���2
���w���>R�Z%�>s:J��-�L������p�:}6��եA����.�F�����bEŘ1s��~�7��o��;�*�$*�����;1�)X�~���^�5�$E���v]V+�n�n�وG�8a��P�����}���E�٥@��Օ�.�.~���hlm���TY��ǌ����O��5�,2���bPu!.:�j�<�㏟�[��(�Z���D�g̚�ӦMA��x�޻��g���Pg��t��J������%g�+Fɋ9���b4N>i�v�
$]�����ُ�?�
i�I����fa�1��+)�܅?��)�n8�eʀ~�%���C���s���ܪ�"cH���v<�����f(v6����_�l�aQ"^G���k����ݻ�e�b�1l��"�2a��&\v���z台�ܕ���:n�NrXk��}ظi���ղPg�q��KiY�93N��Uk��REx��.�W_y9�[��Vaђ�X�a�Vo��:i�w��T�1���ر{�
�	���x^<^֨��ڿߑH�[������䒳$zr�s�1�����?�I�C1���%��wie�ϰw�A�{�%R�w���#`���c'(��'��;;/�?	��K�cY��������h�T�+¤qc1t@��&��p�E೥�4������n�ıƳ%�|�*���x�Z�'���K/�a�����g��w>��@�ȳ��]|�9�joG1�$%�۾s'�n�YאNF�ƀ�
�/����%)1&Mf�Q7)m\F\c[>z�u%��K��B!�6��QIE���r���"8�E*�<q�1(,p!NR�a�1���P�@������=�rL�ȁ��)���3�7�  � ��^�w��mYÊKN�qם�k�u���"lٵ��bT�6Z::��Ã���I�<~2:��$���P���<,�+���3���K�������w�q~{��rK��/?h`���%2��?+*-(,���
�aُ�#��]Bw�i��>��,DK�"��AP���u&f�y�bl)�~��["�,��;�o�W�`���N��_� ��@�e��a����I�R:r,n��v4�6���`��W��E�,U3�(���F�ݏj�{��Z��W<�#���K"���O�y�5�
w�\"�W��>n��;�������x��ϴ�H��n�]��.2~�o|�
,�0^X��GK����c$��>��[�MN�����U���p��p��$�2H�LZ�7ˇ#9SGK�����o~���k&q����]�x��$7l��;�1b�/�Q,�[ÿi���g9�U���l�O�w��7������l�
�=Bg@H?8y�x�[�A�p��2_ˉ�b��_X����otuF$�*|��%����*���pP����C��7�����#��)�u�G���42��U����_|��~1M65!��'�8�.\�-@��e�r(�Z��h�X�u�v��l���ҶW\x��@B椄��zP6�!=g��n��i�o�-FN��"��w��$�y��(%,�F�����O�A*|�B���^3?\���=*��+ٰ��"�{����1��?jσ��a��,Ƨ�7���r<���
�&j�b�)1�K����93�I8��Yg�8��Q��v���������6s&�����^�ߴǎ�X����<�	ͽn�|N�qfξ5r���9(��K΢�+o���.�Dg~���;��f����ͧ���*&�k��c����+�?S��rLsS�8�Lv��,���JTkd�)٠C��Z��^���ZS&ߙ�񆞖�vve���+�ߞ~�R�,y��\D�x��>�\��>�g�:C=^m<P��H	5��{���G��ze��(��f���D@ӎ?V	�(�X����$(�j6&�I;���'?[.w��nI��o����b ~޾SO����V�;9qR*I�1�V:o>�b���BNI����w����K���)ah�d�n�A��'���;n�V'CgN!���v+��K)r�S�Psr6��Sf���C}��5�4�F.���P/��&X(��$�I6�+)���{�09�>e�{3��;�����4�u�s���"�v�jFKW��27�ġ$l*�S���뼈���T\W}���]���nڻWR�$RV����l�������I��j��Ix�z?����Ȕ;��iu����
t��L��������d,
�ӑҮ����2�$N��Z/�5(y�E??%�3�H��ӱx��)���Nr[��ȿ�S�������/CT��i�K`ፇz��J5~�T?
Ѭk�5�z�+��1�� H�b�Z�����[G���rD��8
�/�@!χ�m_�5p$u�I�oB��0� �.��V�2jc��mGiI!�2��ϔ�K��8`��R��r^02"�?;o>��=�z�����I.�ϐ)��N�������S��tiݎ�	y{%z��`㘽�)�X�]֗�$��zJd_,
p�h��mQO,���&i%�����E4���w�5q����.F���$�r�܈��K0�������W�eO�^�
�Ew�C��
��C��A�z�r�7}�>�9_��:��N�u�h;�xr�D��(+�#�ȪS���h���h�h_D��\��5��'$㒍��E��/�R:J��p�]��t��{v핵�a.%K���G��$�著��차�HD�8�gI���>PT�����A�f�k"��8�m��:y,BbtT#�d�+z�mb'"�)U�"3����O��p����T�$G~		�9#��h�Ϝ�	@���jN*?�b5x�8e�'a=gH��)�a�(w(� }�x倄� ����3$)��Lڝ��2��Q&�y�����i���{i=�fE�vIT`u��JT
��&�].3���xY�j�����"��i��,^�j��w�)a�䠘�@�_G�i 8R��+���x��X�ek��5����TF���J�	�^t��S�4�Jҙ<@��
���gT.Be�H������9k��@I�)(�¦�}w"_Y���W�1�A1Py�>�O���`�BR$�0(I�A���5D�;��s�����R���?�O�i��(�;98�"N6�d[7*�A��RR�N%nN25ыm0��a�W�\{v�ȈO<�<�'��86P k�Y�ci�=`$����CUR\����������i�#�bUUJ�M���TtoP�M��$�a��F��p<��gP���=.9{bgu�L�y.FT��¼�r��v���#�����և�2��t�ǎĮ�n�%���H6A��Q����Qph�-l:+)���Q]�aÇ��@B���w��bD�R���!�")�ʊ�6�X�W��^V^Y b�F/��8��h���5%T� ��M�$�<�_,nB6�zc@ʬ�1����J���� TR�!���9�*vU�äv���U=h6�� L��&%EE���zIb�>��P5�(u7<�,��!�P1S��B�MP�'�X�	ͻzbp;�NV٘���(zoEE%�%v����� V���Q�٧R���̹���ޖ�Ht�L�Dm)ńD��R�4¡����,�@�7O	��Z+!wFP"�P�x��< � р3����� �G�MR�¿90F(;�����^|��r��ʼ��34?�:|$����5b�`kR�x@<�a���y�*y�!��%!���rY����\{�E�4;/��R�I�#���t��PqK�5VF�o�wb��J��BT�,�8���d��ನ\ �0��W��]=�8�HW����PD���Yl���j�G�L���J��$�Niq��ӧ��U[j�UO�)�`i�+)��� �F�����,Y�D�&��b��i����ߞ�s7X�%��q	���_3�*${��Qs�@<���fg�au*�zĘ�h����J
��(F���&w�FP^U����H�F<���@��.�0q"v�Iz!Q'{㱾�8��zx7λ�
8d]ñ���!�AԳ�`KF{PYV�{�%ަ7�T�O~&)�QR㾬F�V�l��H+"�ML�x\�,TO,� .Z�U�H%�G�Dr�1j�j�fTI��O�s�ϧ��0��S�&���"I�D�����x5r-mU^"!X�!��l��~-�������|��R��b����T�$i�b��iX��{��!�4�]6�Z䰌�\�v�v�Ũ)�P_�,q�����&�1�|��TTC(e ��v�
��CT�7+����[��p��_5G�ĸQv���K�C�T^T�ו���)��5m�<?�,E䅴k;9.�B�D5��=�4���k((��%k��n��
t5�S��Z������<$6.��'�9�I�-��0�gB۱sN>��-N � ׄ�_fe?[:�ʡ�����K���o��DD�L�N�vg0f� 5�lc6����`��|��1q�xt4��ߎn���)�素���1:���q'GiD�/�N�H!'%����ͫq��s�l�*E'Ÿ���<�p�aJRcw��G��LEe��ΊG��:0qd��b�d'i�$��q����ȁ��=K>_�L`V�mp@�;N��n]z�4lݼR.s���UP�g.��j�75!P���������p�2PQ�D��7����|w��'��{$5u�����=;�� .�t����$��mܾ��q:�n���s��/!@U7J@�z1�܇��f�#����c���t�����hG�zP(���+~��?��8�IB�4��O�u������������8�=����/�E�9��/���� �%��B�.�ط}={���ٙ�!/	#�Ɯ���_pBb08Av'�JV4��*���������ڹx��$*�ߢa����@YY1���$��y�
�A����e߭���W��%s��G_|�D�C1�^&�㶢�;���˿_-�|���Se�l�cb��������W��6.�jG��u�߂�b0�rK겫��`�F
�>Y�W^6��6<��?�ٗ�c/�A1�s�?[�!9�-Ln޲U����ɥ��/p��W�S����W��b��� ��4��%\�B�"��b~�b�v>�"��I���sIX\��Y�=�W���ghkk��֋��]��6���%��h�"�H�F��ޖm;0e�@����r?~��c(*(c${'����n�.�n%q&|��H����˿U� ��]͸���������H*�S��ÐA�5˾.�z�v 8�C���TkE|��b����`Ӷ�J���s���b��mJ�����V��4�Y��,X��W�Tֺ�� �V���/���+��b�	p̈��'��	c��J�3F�K�ev��q*,b�.�d.~�������JK���_c��`quI4���-p������G"� ^y�-\q��i�*<��8����y#�B<|іg��z�Q~˘�:
l��"�p�Q�r�y�F<��=*���Ԩ��A4��C��.m-��y
�V.<�n���w��7���K�G���{+���#:؈r���f�� Q�|i X�[�����c�XTZ�[�/��1��Ĉ����3��ʤ��ķ�aEe���"���شk�N��УDaq����Z��YZ"��,�'�iܘSQB�q8�j��t�<��V.[��)�O��MZG �և�~$yV�!�K�My��?���fM�`�]R�8�����PҐ�T^�X���	���HJG�2q���
<��s���ף���?��;I[x�)��&�'��Hk�\����Ȥ4�u��䋯U��R�SsC=���ɝ��v�ܰv���&���.�����2:��@���x���}��p�BmY�=rhB-��N@C�����e�//�,���7��u�^���L�<�5CB{��w�Ҽ����-�����3�c;3���C��'H��]���ҖR7��B��n)\��8�ͺ������y�	��~ZJ�3��_y���9Uux�ϡ�H��PHs96���`���Q�8�Z�}k�`��������aunehP�a"��y軇�쀫9�m�+`�h����c>V~�.~}��JJ���I�]��y��6ハ>eÐ�𿲐e� �x�9�=�'�vac���-T���߼�z<�O>�j�5�#��j��{�7q��G#Gõm�J4�����ø���4��\�Zܻo[  ��IDATo4t�j�.8��jSN*<���8��30�}�{Ϙʵ/�r�͛��z���XE8�K�Y�|�#��a
�~��~�I������*,���F"��[�����b>v�#qb6�`c"���������#_�o���x9�S�=��ی_��!�?n��e���S#�榪�k����7�@Cߋ������ƷÝ�VIJ�|��݁Ǟ~�x1�r<Ŭ텸kz��q�?�yg/Bǆ/p��oƍ��~�tS-��U���[��P��:g�GL$�6s&n���tݵ�R�ټ�f�z{{�:��砚aH�>�V��ȳXN���!�Y�p�cIW��~ȁ(O`���D�eδ+��z���̼�۾B/�½f��X�:��W�t�#O����ģ�0}�ģ��۟�s 0��	˗��[g��a�q�Q����U3�H}��:9ũ�������W_���nz�V�Q����Hk6m����WBF#׺����y�X��;�`�G5���D��i��UUր�����0*ZL�I3	�'(�$��q"��x��v*&���6^R��|Yw��nk��۴�3�#O�)��_w?�+/�c�C��܌�V�_n2�j|���ǐ�hJ��iі������
���;�k�y��$�*�u��4�\�:�IV�QK�5��ʈ��ց��	���X��+�亪�a��k����}�9�(�F�'èw�Z�pϽ�*�u�a6�՗Ǩ�A��0�hj���y���ܖ�v��/��?��\u����_c��6	��E�/������e՜Ďie4./&�x�|�%�R�[Ôbm�H�P�t|��7n6�?�Az5hiP�@��i�˯��c�<��'B���~W \�x�������6ËZ��r��P��o렲�(����>b(s��+W�!���lP둧�ex6�\)i]v˫��*i|~�����o���)�Ps�GE����g��X����٪S^1�g�ƛZл�x%5_�$.��4L}�Sc��Κ��ͯ���hT;W(~3��B�X�*�Z��;pم�a����&,f|���f�Ê��14�i/��0�J���J����@��#y��|�[��|�]<������ahh���5�v�y���ɾtǀ�ʥ�J/���a{���f�2k��8O7ֹ���0�+j�I�pm��x"au�v������p��gr��j���/k�}�6�w��T�=����QZt�y��M^|�~������X97���e��y>�b"�j�.� ���T2���Ɖ���d
-^�"���2�����[RTZ�`�M��=SK�U��=kL�J�y��&�F2<LH?����=��6|%�8T	�/�\����b,WIL�$=C;QLE]�S�,M
;s3.G���@t���<�h
�1���wo���u��[�`� 4vp����V�x�m|]�eM�Vƫ�����>�?Tikfr�&���Urt���[��<���=�����7>\e$�6;$��uw�@��.��G4��^�&��<(=[��V�����
���a�Z%Ao�0����ܞ!���&B������rL��ȕ���v��3��sW���I�򧿙����+'U���ٗ�O��P��#RQ��|���7����L�l�J��h�#E!!p8JN9��@'�1L���o�����P!觃"��YT�L$S�Ұ���mZ�^?�.~�?��H�t�Gok0��D2 �8tp���/J�+��j�&\|�?�<�Y���x屸5"z����?��̶J8�P7�(���Y���o#���6��҉D�lycrc�qq���[���/����SD��EB<��s�K���K#�$|
I��༔����H�XѹH���S,�xO{��g3p�l�2(ٺ��yvL�:����;�7!qbn���om��Ha�]61j���4ol܈�h��'��%d�[�H{�9�P���Q�ӟ;��x|�d#����Mq�>�=�0O\���{��h�N�Xz/�@%�<D&�b�>�4`b����N��a��|[�1pi"Y�|�*w�U�1��p ��M�yJy�Ck��S�1���������`bҙ���1[o���=E��|Œ�S�*vU��>��|�$��t��s��KѦ��A�����L�h��&3>n�T+�ڔ+�
��$ڤө!^����Dee�2�	�Z��N!��$�&)8=!����g�tf�G*��X�5$�	� 66���/��,��GT����2Ӫ&E�'���%'�%�_�?k����5��+TY�?�D����m��G�b�7�e��c/��a�q�L���j��1�%K��2�x�"�Vǘ����歆Yg�;>�"(�lԁ�����y�1���a�*d�)��}�+�)]W�3
��m���e�f��#g5�X���5g��:�bw�YZ�f�s�W���@�62o�^&j�����]��D���
�����0�!�i�� �3�J<;.�-|���m��.K��3*3�(��o˩�}��-]X��j���A_��򞌤����44S�[��P��蠫���
�_pf������k�	��h6k�b*��p�����z��������o�>��r^�hF{nnE�唝��b����e��ٜgk�ҽc��劎�)!V�֠d5N�+�s��e��WnG�D�~o���|n_i/�f�w""Q'�JP[�XzӼ/`��O��(pJƅo8)
	������e�֚0��)�{��2��͍/1��N�J��Û����A�|�W#W��p�]�����\�\�cgQ�Y�G�9�Ncϊތ�����T�<VQC���\��+�.��+�n��z�����(}i	[��>O#:u����c��91w�n�D*�(k�ì��F�Kd6�cPW�ؘ�:4�NBcM(jT<��!��˩�Z���SH���(��l6e)P�I�������h�@<<))���V�z��+����=���b�1|nCS;8�ocJ�#1�o}	A�,y�/�	ǌ�C��\ֺ�.�I4(&9� 'æ�)S����,D<���rV���	��RF�Wfk��7�,�P`"�p<e�����G��P�{W�CB���*܃q�1Ѩ����;E����X�'U�//�/��8���_q�V���-֩t�aɘ�d�t&�VSnF�ߘ��f�oOco���f*2��t ",Hs-襃��)cCw���34~!͂C�ˠIOu�Jy=9>��B�k2�>�� F�,��}���ʱ��n�H�DX䥁�,C����I�*�Yck�v�659����j�smb6�Q;�����x�x�	�C&Q캺��P�KbC�.�H�GÎY�va�y3콪��0:܇a�(}cCD�5f��Bˌm+o�yӄ�w�eFP����zI����jԑ�1һĴ'=��" ҟ��J���C8x�=��	�!��Q|���k��li OsU���Uj�W�³8�ݎ�w��g���5k�Wf|r��wr���C���{�.�k��]�{}b��!>���BY7b�da�V	(����;[����u)�������Ӳ[t�~��ʋ &Ņ��������ys�X�A�yjo}��O�������Ƶ�!c��An+��[���QG��3f������5$=����e'/�Ƣ��8V�E�یCݏ}"��k�y���w���-p�Ė�#lq��\:���Z}�1�}���K��F���OP��`�[4����>$�.�(TKN����3%��R���z�����=/��Q{�����Dl�bt��y�!% 3�V��D�=��is�󎚝�Ŵ�Z�:���q�I�BCu�%y�?kh��g
���-7aa� �u�:����R]E9�;�랜L'PWӈA)2���_���)s��l����f45i����چ����X�|5�kkQU��E�����>>]��1}��^Y�s�������V9b߽p�)'����ɑ�x��4|?�ůP����͖������7��P�2T����w��B�gXե��~L�1=�8��0i�a�3����:5E� )���}���ʺR<��gZ��y�\�u��6g'���ʟv�5�h-?1�3O\�yӧ�C$\f|�������9Ǳ��8wRy6I���G��_�lI�]�����L�N�6n��QYY�2˧8khIq	W������3Q���q&l㕈V�����cݟe��(A�����J����7�����P#k�ǢA(Z��� �>�DvoG����C�?�c��ⷷ�ͨ�E�j��Wˌ0�Oc���}���C�F��� ��ik���ko�O�M�-���k!�,ƇFp�����0ֹ�1��q)BkΠ�+.�=<��yΜM�kv&g�W�!,<`?L�a����2�=Ui\���u2x�1z~�/hp�	�VF�p�v�;;�jEr��FzҌ��pA���������ko�ظH���3�[�T�.<�t#"��NZ/�O�H�z��o�_��-�&m��߯C�8�q����K��;1�u�Oe\�lD`�C�����W�b`d�D�e4��0B���A,:�zd^�QzwAX��-��Q�PQ��>
������z�R�����k]c�SZ����10��K�$q����+L�W?����?��~*�=o��%W�FW="���~f�j+12:�u����1�C�7��Ϗ��TI˗����-�ч�i��ؼ�g����\�G�����w.�{�Q��Z�Wٺ�.(���0�6�d����2J�	�1����}�8�c���8%�sBX��h�
|���==[PYc��i�4 ݈��Y�������FD+�fҲjټ��4zߦ��c�����@�?�G��=@c�y����+��/��W�\����y`��e����Z�{�噬�Q�*0"�m:����W��-��|b��c�Ia��{i����ߡ�����Ƭ9����Ai�����\	�J�+V~@�����sf�����׫�J)�-�,ߔ�(����M��q;3뵸)Lo�ӾߥA������rq���h����f�믽�۶Y�Z��B#U����6>^S�	��g_zۚR�~!�yxu��~�ш�H��&����l�OS|��iz<��e��՝�X��8�@�n��ي|�m��B(g���$p!�cϼ@x�Ё���)r��ښ����*�d�r,1���Fl�괖������K�!X	#A��J�����F�m[�)ƭZ{]z���p�7|�
�~�=(����]|��H7����S�h��Eg�F�B�՛�Jz����E�p���#�����To�֙TG�*�g�R�����	c(���&ėR��G�x��e�U~����&��N��4"ܣxM��E���RX71؇���}�q�C� �9L3�ռp߽�Bto�d�R��9O =�|'��M9=�^��g|�1I�P��rJ�e�8��0{f+�{��ܶ3���m��3Dke#*cQ'x���{ �
��-m ��0���qã�����4�k6Ha� ����O�so,���>㤵��C�g骋�g�R0�Θ��߇>>GUC�U�*h|�oހ�o�!~����#��A��&�p���i��m�u�nD�c��x�]X��D�.�N��1�|�9|��k���k��.~�u\�槸�u܇ז��Ь�f�a��;����}����o�`��0�+!<����[�gIX�_�؂�V.Ƕ-��F�%�p8d���`��(�vt�T��jWW�%�h1�;f!^z�MD*j,?�l�4~ɢ� ����E?]�ܤ���!NH��-8c��xc�'�����K��������^D�M�>��[��+]�p�Q�In.PFk]E/r>�d�����N*E8~
��Q1�Xދ�>X�Q��Y\��u�p�ֲ}��O�CO,F��M�F��3o'��� '�Y�$/���܍�-u8����ف9��o��/b<����)��?�}kG������[b۶�6/3o�N�c��x����#8��xo�*��Y%&��N:��:�Lm��K��;|��j�sfN��Y������5��O����Pg�,�w�����H�_z����2$3.S*��p���Kh9��v��G`�ko�x�R��^���hk��x�i�,�ǽwab2�X����pʜ��Z��S[���b庯��~匉��o�=��3RU���1�����LE(��NӦ�Eǚq�؆� z	/}�1��h8O�wO� �\\3k|����;�Z�Ǯ�|��T�Jo������8�{�y��Ӕ�(�� f��]y�|�� ]l5��o~�3B����8����xi�Ȧ�:7�#O=�HxUiZ���x�wp��Z[yp��&Vn���9 �<�#�b�����D�5UH�x�̘��~r6�[M��A=Cי4J���-D�#$��sq���3t��Z�a�>��ghЋ�����s/3;���,_��9Gz�M�^s�%�����a�U�:{�ȝw`����B�����ۿo�����U_�F�a�����w��B�=�����h`@�ڗ_t��=*���3/��	s� w�;�:�zÏ��g_^F���ћ)N���p��nDO�V�Kli�1���D��V�1,<�#9j1�`"����6ɪ̷����u�;�$�o6��ӧ�w>D����c�=�Pz�^��3h�o�՟��+ɧi�_�����?���QkK=^y������#A��Qy�
�v��>m1�dbV:��Cq$7X2LV[G�p.�,��N8�p����;�?���j�$/�|�j~���;'��DS}Vl��
y��8r��i�ǡDrus3~����;�0����y��=���P�D�����`E��c�Д'!���u;��g�no�j-ڛ;Fq罏��x���,%��	X�Cs��*cF��=4�%K��f���-�dL+�~�E�.Z`�7�C,�ҏ���0��OC�B���x����:���܍چF�	��&�����(�.ŜiMF&4�,,_�A���	Q��OL�����F�!4�L1�	z�M��xt��E��c?��}p,e��A:����Q���}��|=��
D�q��ٗ��6S�Z-��e�&4�v�Y'��T_e�P�v�?��w�T�1L��`�ˍb~�T��{p�a�̟��j���\�(�`�tq:��|ϼ���N�l����Z<��K��͹�vL����^G6���B�:�����~2��t�y����A�7���4�Zo?�\�&X�%�J��dHR�����N�},��*֛��~�틙u�����λ�.�R0Le�`oà�i���_��XD.�}%�?�Dk�t��{��~�J��~0>\��}Ą�<��"�i�^�`�w����ڭ��1���������j�v��F�mm���8����V����n�M_N�O��cO<�
=�^��>Y�]Y[¼�	4V�M��:)���L#J��/�➇�˰#�4��4W�،?��o��.�����1k&�aQ.@��	Ɯ���w=�<B���x�B���?�v�7q��r���0f��&��+�@y3~�?7�;bz��������꯱��fZ�=Vnl7���:	yн��Y=�~�St�Z���A>;���b� �� �;�͈�.��LmiÝ��#<�r�����y���������@-S2U�%����=�'S���R��1�R0:zM����5�*�� ECP0z]j���g���к�in��/PY��hӨV�������c�}v��W���?�:�wU������+�u��4aR�zI�{�'&ѩ.Ȍ���^z��6Yxy�2��I���
�59�����AT�+�����W^x&b�r~~ԪV:�yz�4�W�qF�h$����?YT�N�w8m�jv����@�P�f��)LZ�:g#4ȯ���rx��8'+��M`ZsV�ـ���Ѩu�7����bѰ5�}��*T7�J�1nK�Yzo� �1�˗�;5�Y.�	�+5n��sУ�;fJ��g!^|�k-D���"�j�[MzB�c�J��R��/���5�3�v��,���I�/H��0�7�D0_m�d×*��a�6
c#D�v���Stf�$�4�s�3Ѝ��qxS�%CD��Z9m0���e�X"�:��P/��9/l2K#RcI��	�&2��#UW�^���OW�����b�����-r�J���ћ��|�z�5(f� �<�w��002؋7[�U+19�AJ�)A��Mc@��J��ЊfU���s��l�y�47��?a9u��j�������i��%�p����K��/m,;��3�1^5�i�[c�"�!�-'RYş)a��٠�����7F�H4���>kHRk�ˊ>�'Y�k�6��	����R]����T�\F �)���sY�hC��k>@@�3�-�v��U���n*�L}6��1pU��E#��3��wT�T �	�85��D����I�+jsn�:�*���Q�BZ^S��d�5H��I�?e������Pv^�#��<��{�O�jb�٪�vAD�7ݕ�u���Y����:4��(��1�Q"�H���$�XE�5j�J������%I$������c;��a���-×����c�0{�㸊���&�B!�K$����J�$��%��?c����p��O��W�T�N��B��rX�g�f�C4��ҁH���X��DfQ"���)%{c�$͛�S�r(J�M�5��g(�����p_�����B�����#SV���� B�������"^U�}J%��]=#6�ю`�܊���BU_��(�Be�-y�|.�U#�Ǜ3^���:��LN�p�}&�����d�;D�rU:#��z{��Tی�|�*�aJR�n��I|�ܴV�H���\��CɨӖ�H*�m�:NE�&-�Dr̔�4}��C�r�7���[b*�$����ցR�nH�6?��f����(AOXVY�"=�ȃ$J����(����\�	�pe�s@,��h��IC�5�$�b�A��q�F�G�$V��;|!�=[Q�<��C�F��G��X<j�T��O�6W�(�ГG�+4���2g�D}Z�,�8� �66`0ىHM5�z{��h�Rb�
0��Fj2e�o�ݝNd>Sb}r�J�m�b^<��q����Y��$Z�Oq�j����G���!=��Mk�3�)���p�*ߎM������e%oV��������)���ށ�3���7?4���1|����A�./���s�|�6C>��`�\7hڱeD�.^ZQ�k������_"�1�,�/��M�g#�g!/i
��4}J�K۝H'Ƭ�����>���F�G�ӑ����RD[��;{:G����0�д�gHZ>�1��yD+�Hd��4�!#�VZ�!�VL2$�=���Ћ��!"�����؇�v�7�B��is�y�f����zv���4�V��vD��|�B�a|�C[e�);�As�rĒ�4�":�ysfcʗ[�)OH8�P��#��r�!Kx��w���#g��������S��1���[h১���{8������+����2��>¥C	iz�C�������F��$#��?��5(��.��VT�x���uv�5���W{ϣ��ʣ��"/�!�e���8�ŨU]�|� ������_�������:Ӯ�R�5U�]=�
$)�P���~
��/g
#��ц��� :=��Dm|���X��p���z�	��A�1�N�[���{L$b�4a���w���D����dFQ��x7��B��k����&I�����k�\/��8pl��<�U�b= ��p͕a�v����(�iz)j�������[�F�f�"2�J�ea5�y��Ito�QxWnJ�*�mz���X�mzk/�rA-Օ��k�4/Ġ1�:���pi�N�H�T���1��Z�@��uD�A�y�"���bتy�Xp;F�P<=ч�3-��N�y-��{�D?�8�tIF��'��?�4�Y+�jE��n|����'��qz�L�go��u��x�[��K�������D�*�ws�Ax��e�m�!:	y3ԇ� ֮E�(!~�w�h�VC��w��e��}:n�ۿP�Pia`U�}\�k/;�DbA����	Ջ#4*��X��7bN[����t���}�?�:�q��WXJ�%�E���N�٦��0���w�Q/�^�����?:����&>�7�K��Y� ��`?�?�$�?�����_�W�M<�W���;���h��5����K 'kts��0v�?��iEW���w����WЍի�`�E�5��g���]L(�LL��2\���9����!��$w���K�x	%u0��S�*�U_��v��i�ԭ��4Uct��Jo�ކpe�5�(�x��q�A�"L�př��Χ�E���'j"��ւ}1cj��9z���Ɍ�����}�c�s��4�	�fO���c�H�g|��˜p���r�2�|��Ʈ<�e���hk5��iյ��zg�FL�`N�Z�}w�g���@�e���	={�n����~�v�ϚI���uW_�G�}��(�Ì�z�o#���D��/�J�����{��Gp%/���.=�<���<��9�UG�Z[�쇔�5���Ͽbk��PL��G��l#��>�(T0������x��;�l�٢��&���_��.Z�Kd�pc�m|ם6��k.�[o�����3�D�8f�� �!������54�W��'�W`��Ga��+q�qG`��v�z���Ģ'`�gXapE]-z��Ot�<6ئ��.�o�&����:<������p4�{̞�ٺL�1�/�Q]�y+|4F��gx��p��`헫�_���I��1"Y1aUb�]vB[s=*ba�O�ɧ���)Q����^��(���ڋ��;o�%��N���Y�0���1ޱ�V|jc9� ��S���?�����p���a�⧟Ay4�i��8�ګ��Ո��yν�R#�R�%�X������N��t���}�%�ʘ)$.:��:{�) x���B���غ���яS�85匛z������AIg򓀅��埣����
��f����?B�q���&s�"tm��:��l\o��$4>�t
��w.<tz�7��O@�f{Wji��A_������Q���!�4�Y[��)�T��s/���Ɩ-[q���SO7��;-n�y�PS��mAcc#y� G;��l����c~C5��F�����3�p,mHG�I�����q��K|�����ϼ�
�dG�;N9�=��s��tۿ^ge�/x�7v����d�O|���,}��|"=�j)�>w�AB���v��c�M���,^�t����D��j��Ye��g��@'�lۼ���6`h"�G�����\��>����=���q�������6x��&��8���^0*Q
(���|�x��-�b��q�׶?5-('��l�c���-|�OV�%�[���4�%�����Oq�ӱ`�9f�G	�3�ǵ�J�ܸ����"��\)'��Ž��Gq������إ!�sEV3=���!ZU����OcKG���	m��F��;665Xxx�Imv&=A䙒�R��w���#�s_����#�H�q�C�q�O~��5_��E����e�����ޯ&�GF���Ĥi|e��{���"L�E0�i��m�m!`f��梊|�OW��{D�B�>�����be�w�\y�y�^�
�\~.�o��/A�Q:�a���A���cʗ�e+�j���܁�������f��DL4j��Q�/�V�Y�ѭ�p��{����ٴv�Y�T����G� �����#�������P�O���9�e]vR�����5	�c`/���X�$4��9��d��,^~�-q�A�n�Lrn�/7ԁ�H�2�#��3v�8�a�)�Q䳄	K�^�*N^t"��V�0f�M�%2ʃ�u�:45OųO�`�_�����KS���]��G�,�s���}�r4��S���I�����<�V��k�,CC˴���2���xd1~r��бm��:j���!��n��[;:�����D/�K>�*i���F���S�ޕ�c������#d�%�T��ɉ�8����%��gJj��l��o����aƳ:�p'�4���0���{�i�xQ&K3C���Q����>�����c�q�[���1�I������dY�H#��B+���r���̋����܈�[7 ��#�u�,�:�}��U_��/6X�0�CS����7m��C���J�C��:���J)���yF�-��p͝s&;5�X�<ú�{�5����5uȊg����e[�������ϐ+)ʀ��!Lᙗ^��#Ɣ�Z���T����uJB4`+׬�Ko��He��i�OQ�-�3��P�ﭷ�'��;1�i�Z~i����ʚF�鯷a#�Qo�f���A�|u5|��p�5W`jU%�x/��N���vgx����+���e�<�jqs�Gh�dH~����?�!6oڄ�͛Q�CH���ǒ�ǽ�ǆ���GJ���E�q���[p�?�J�C/GO_��t�������ޠy�m�ۑD����O���I��.��mڸ%���W_Ǣ�dl�1���eΆ��=���<�6E����b�.{����/:�[�Gjjn�g���|r4���}	Q.��C�7(8����S�2TU��|���:�V�`@�O����{�y����~������$ʫ��²����ZS�DB]�!�CN��g����PY��L�jP��L�
��|$�_�}N>A�y�n����I�7����F�g�R�V�R?K��
E�>�{�3�"<R^c�J���ϗ�Qڴ��	�U[<n+]Fy9��5u�!46Eģ�������{�m0�Ҭ�.�w����C�إ�r_�f�i?_�%G08<�{�Ym�Jf
>����Eq���e�Go�@�?�0=x�
"��6n�qs%ȥ!�	`g�Ec�e�
l����c���F	�5 �8�ƻ�*�YCS�35j	Ȝ3�)��iЂ���ށK/��9��Pچ�4.��6a6�Y<n$>�J�= V���I7$y��~�mvЁ�M��˭�j���Ƭ�f�z�j���㷰�V����byˤ�;������S�Ik�R������C��1>��k�(����sp�#O`��sM�3�2N����?�W�j[��x5�p��c��/��_��_ร�v��чv:.͎}��稡�Q"w��Y<#F�\p&��D?5-S��7b��w��T����p}6Շh@�<��M�i�.�*I>��k���[�^j��3ʬa*e�@�E"��_��1k��"Ԋ�_�z��Z����p���T�7�O�?:��B=ieHyoq8�͍rZ6��������lh�Z�sVI��}?��'�Y�'gm\Y�Ƒ�*d��6hQ�l�Ў��g�0���e	Ǽ�&G4�Z&V�|�L"��qdW���h�r6����L���K�%X5jit�}�he=r.��t����hs#�c	�¥X�f���}ҥA1m�x��^oiH��Ryک�m�7�����!S�4��[iW����j�+3�%�h��3E��D%�@8ND��'_np4Ex�z�sz���(��Mu@*Y�)+�nT�� �t�x��O�"�w��wATq���LE欐���Tmܦ���ҷ�^ǲ^|�b��_�-s��cƨ���
�Ç��)����x}+�~�%+W�{ӝN����5�o- ��ڤs�IJ���T�6a�-V�v�(��7w���4Mj#�>��Z,:�&Y��fq4L��]��r>;�;��ct<6IZ�X�\��b���O��J��	��.�vts��lC��]��)c�jp&�]�ФIK��ä��c+"P��[aL$���(	�U�9BT�Ҵ�#�Q�wuwB�MjQʈ�Ϲ��A�c(7���0�ִ�(���)%.���N&H9 �JW���`�ʂk-���l��]�YŨ7Dׯ�¦B�]8}�����ao
���˰�F�%9����t�e|p9���"Ѽ�_UI�3�l�P�(��9q#�����Vl�*:�y���������9jz�A,��0Sb�b{���z8��]熈Jh|�eQ����LIXJ���LD�0�@z^M�\f,=A�{�`�v!��<`&�L֊��F�������Lp�w�����Z O�#����SSޡ�w�A�Uu�Sxq4�2�:����%9!*��@��-�hs+�)L:�:h2R����|��]f9	��Ș���%7�f����yh��o��6�rHs�G���]��3��2c�ޙ|�!�Q�S��-����j��r�~���|�b���.��򥭱���^��Ƙ��bє���T	�=�DkJ��2+���<��E	x�|�,q�'�z-� ��cTe�{O�y&�0I�2��Ah5P��QLO��|�����7�;b�%�������~����,�-	�����GK���(��z��_3���S	��k�������׸�Fҕ�zq�Ċ����[°Dbc���$S��Hg��=F�+�A������T�� )�ē�)k�Y���'�%Q�,R�o�_t�
�] ���[W�%C�J0�r�E��D�k*-��U�E2t���p�!��
�����+XK�2�`�&Z�K[OV�6A�/ϋY��LL�6Rfy	��J��D�G�	��-��1ck�@f���x\颪[�<:�[���F�Ρp.�}�t�����y����^����Z����J� E[#�|�X�`W�m�@��P���q�-w�Ky�!@RBzǡu8B<%���M�ʜ��*x���)�o���9/;�4���rIhJ'�GF����|0�,� %��b�2*��rc@ݖ��dx�3�~!�4�Xh�D�*}v��v&z�� |�}�YØ��D*���fkF�����nk-��r�����ُvY2<99n(A�/�6!��3Cu��_��khӻ����5>>��	a̘=�Ш�(e;���q=^g�J���xr����8��C;)�+��@����v��$f�������c����s�Xb<*:���ݒ�
O��2O�K�P=��.�8-sҜ��<��W�rTS�z7�$V�T���
��ܬ��:�B��M{E���qx�#��~��	�'�#�-�w)�XQUm�o��9�y��ө������NC2�2f#ux��b�s��� g�{���Kи�K!G1o�,�ҫ�<2<���-X�v#=g��B5\�1n��4.	��$�T1�yAA�4gk6������m%�%y0큦[j��8��hX���'J�j�Fc㶓jC^�$�c8d�ːO�"���o/d�@,Va+���+��`��+�e�޹���rȌ�c�=wA\}0By��Q9vv�`��mWT;�s�%� &1��1;c4�͝���.��U6�r?��T1�.�`)���%�5��$�M�a��w��=��c����)X���X�q��_��\�RW�;p���?��G($��������w��7��a,������7�WE�o�`f[�]�@A$�lݶ���?�(ע�Ǩ���(+.�[PH]H����7��ܯr����J�嗿AyM�!�΂5H<F�$����v�8a�F�%*ǉT��J����`Ū5(/��*[6��1�Kbf*�'8t��8���_����ƭ������_�bQ���I�Wx�ŗ�3�0֞B	K��Zq	��wv�ګ/�g(Z�]���*�Sl��ųϿl:�@QJf*�adż����Lᅕ�nr��?�	��HO=���#�T�� �J�Z����X]��Gj����Y%���	�|�)���˼����Q*6͎�����G�VPL�ҼL2T���٧���{��ube�J��*Kr�2<�W]|6���MM
uDf5����'�g_z͆�R<�2��O��Q��ƧG��p�A�`���4��B>���3h���/�Xޠ��DFUc�N�T0������`^X��&��ϞaݛBe��>w>�8*jj�S���wrJ�ȉ�-Jt�?I*F�2�gh�6��S}���b����D��`��Yd�.�)j��Sm<;����bL�j1�����s��gA9.3v;��A�*����؅�V�-Io'�����n����=�__���41m��t"���8��et�-S�1<2������Q��mlj�Z�c]�j����όS��E���W^���������ӡ��ԏ_����ֿ!Z�d�:B�K8�^���}v��4�����M�r�{��ù'��_�Ϸ��3�M�`���H�Ao��r�O1>�ϻ�5B���qG��{�??��q��	�7Vx5h���Fn����sNüY��$oi�$���<�1:��6���k��K�%�$}Ǯ��b�}�E�8r��e�2�mo7��":����	��[*�(��JS����%o��������`�ޤ�m���{߱�6�F>�Z9a]��_�ҋ�����5����:�p\t�2}�A��P�2���n�C����$�� .;����SM������A;y�#�B8�CxaG	>$��ϫsO�>�����J*�v��T�3���?Y^�q��e��PFU<������ğo�-�g�V�����ɱ!�w�"�PoN�yj�͖�q��t��xu��Mn��;�=�po�=� L��Hc�v�#��\EW�VLm�72XM��l���o��<�9h�=m��/M�^Bl=c������4�w�s*��
P�PbW+�kz�q��K�6�E?Q�V(�<��$���_�AGO�u�*W$�\�%%zx�.��Es�5u�Ñr#C��R_�sN;�>�$Qd���ғ2Q��CDsC�%+*ch�2����<%	wm�w.8���^�9�B&q�j@�����Y��*S.��jz2��p%�+
8t�}��g+����K�5��@�w�Y�!�S�p�i�TTVb��½q��k�����Oh����F��s�=v3�5��gWQ���шir\�؇�?�N'��<,�X4��\f�{ݎ;��K:�Zg̴�'IB(���,d.�A���s�����hE2E�.�C�:�Ӆk.� 3h0�Z�0���&��UR^#���=
�D_��ڐ��vy%����y�;�4��}����Cg{���XtҷQWCX??28dJeZh]hMt�&�h����0|A����+L�U�I�����^AX;n���ռ��<-��",�$H���]����7-�T39).�*u��{��eԋ��k�P�4^���a�.:v!{�EK�8$�+C���|���5S0���4���}�V�?w:���OV��;�,�-]�Br��J�1,���ɍ��͝غn5*bDx���F4{Ӎ�����h�-�.dr��|���*�po߶.>qX	L�>_����l�!�%�����
"s���O��1h��^Ǫ�����_FMu�et�~H${��N�iHư���:�H�i���[4J"6
��w��d�F����;����2G��k�����S�ϥr�U��<�#1��_�?_��6�y����Q�{�]w����"�9b^x�-Od��n|��9=Acp�CBKcӺӮ�ӭ�a����#r�1�0MV"��NX����zAT>r�o��1�m*$�;m�p��Wa��.47U���
��j|��ST��k.�oo���mtp)~"c��?�����u;á�ڦ���P����{�9��yҪ���tɗ.����z'�$�?��R46�4���ϸ�g2�g�c�R�]p��h���ӯq�M� ^�bNT%�9Dv�Ѩ./���oeN<�4n�RT����KcRƋ9Æ;?X�5+��1����������^�}x踍�=��[�ƅ4�;ͣd(��;��K.��Q2�u�����������҆�ν
]�yLk*��O��#�##��ƕ�]��5u�=����\��y����0��7ނ`�Q����?�n�ޕ�}�,����'�����M��B5=ɘDx��k�<=�(��W\nM\����}�5,�j&Mȍ�v��ӿ}�'o~0t�ʵ��]_����j�)B��D�?�c�A�C�"�?�Lz!�|
�~*~���LG�]0��ӛn��CX��>r�SX�n�����x�Bn����c'���B��B9.z��:�q�C�ܝq�O��l���3mS������9&��K�����)K��sښ�RW������T���I�2�����jZ�Tc��9<�AOĒ�B�z2F�(���;0�_�l��v���02>��	w�܇��;7���N�0�߅��|�۷���G7��@i_��5�7�_nMoW�M�b��:oτU5R\'	��vb��V�������_!^�0�qm�@K��м���mV��_��(+�0ԧ�8�K�*q`~���Q�<�V�pm_�`%��q��ǃ�ӌ�U�JIX���ٳ쟱�z|ĉhh�E��v@�1[���܊�;De[142�{�5��i�^u�ظ�K�:�p����{�j��D�+�|���n�^�33dr8C���y��T��+476r[�n#n�����"J+��՛��ܙ���;q��k��܉�˥���ꅆ�{O��t��eϽp�.DuC=Қ��gh�~w�?������/�������.C0VmF#�˙��4�l��7��h��ɜ	��C5�0�;�t�bA�oXk#Ci'�׸�ԩ�H�uY��9]�B�ͳ�Ƴ�Z,���k���zB�8~ᡸ��K��>{�fDǱ���U?D���)|ӱ���D]x��ǰ��~�K�V�Ï>�:6q������.�����ܿb�9��R��AWWf�0�S�&T��S�n��o(j��J����f��j�}=���5���UV�QL&����vz�?��� #��s�'����� �d�HZ$�+����_'�6l2~�$=���yk��F����%�r���o!�gjm�a4����,w��Q�H5�2n0���G��q����`C�$�o�.;ME.A4�܎圔�ʘ�:��?���!��:h� �@���3/����9��i�xT)Q;n�-��,7S���h�6�$PE�4J�۰O�悦��q��bR��X��t���?G�RS���MsD��!z�ql�C�*��qV[�?�����C���1�C,V�?��!E���&
��1��;�3R��J�Cw�*�D�U��i����݊�i-\�2D�*y&���ci�Z�	m�d�n��C�p��Q��������(��W�"4��o���i�B\�|n�N���\��6YV�| ��n�-��ȮV�H��xᕥ���Si|'i$��O(oIx"�\%�ip��o"��-��p���$<���<hm4d��^��*i2gG�T�	C�t6�W�[�*������S�����`�+�c��Z%��w��נ�A��(�`*WDR���b�;i�;�����5�����;�GM\a�&�'x?�y�]���R�Dܔ�)Ի��~��k�k��������_(,��b5y�ar�:�3$Vj��%1��Ǜ�;M8f���(&n���
�������U.�`D9;zà�gCJÄ��=��Kkä�$�R�#�?�������r�6��+#�2�M������{��fJ0�����)�	0֢�S~���ohȈYrf���|�-"��'B�GE�АJ"3>�?�j�zL�~
���N2�l�F�e�,�1��5�/����&}��#�X��f�۩��r>˲�$9�M�٤��i3��ދ��z�2�s��>#��Tm";b*[j��ԯ����#��M[�'�˥����E$�K��Ƨ��W�&jHS��c���E����ҀÛ�䬚�4d�.x���.�=2l�X�]H�<�[�(���T�s7l|(�#QeA�Mi]�#�4�8�7܎l��#��1��a��-�j������v<��*d��|"�������rb��嫪�`Ú���@�z%�w�Tռ�
5�/I��X"U���9�!q��|Y��7"�s;c�.��\U ��F�	42d�T�$�=����ڽu���RbzxR�1��4�[�'/�zz��]�Z?MCKVl볼�ZBܟ��>T�+�HƬMD�2�s2Κ�3��zjl�Q�Z��\T�t�ӛQ)�xW�{\f91P�A��U����� �_���dD%G"�l:1%��h��I�h�3�㙗r��oi����v�i>�[����e�_�LR�C���hBҧv{5�9�/��@�%��颗0�
�ɤ5�H�:���aU�B�tE�VU��-�=�)������8?n��&? �S%�mĪQ�H����s��c�v�I���0����8Ms�����51�렃�E�66:b�$�#�� �u�y^�Q������h�\`U�<�0��2�.�	#��p��:{5+e�i��(���] \+XG��?8:$i^�hM5�C�ڬ���u��O%���Y49Ǣi�����J]|�9��V��Њ�`��2OYQ5%��gh������v\l�y�G��������Y;�_��Dр��9�$�v�rG��-%.�]�`��21a��L��	�#	z�V5�@�T�!%7����z�����@X뷐��s�$!�H}�D��P�%I��I۬�@�r��YmX?�!�{���/-�2���[ّ~��9Mbn���4��8y� ��*Pr.���d-RR���F��9 Zΰ�x�ˉB*c��b�(X���ԅI$G��PG��D��Ms�,�����7�"�C4��{���x���Ռ����0��X�&]vf��w�g�P����2:��J��D��[2<�U�aoZ���,2}݊�
3���1[�i��$1BƧ�m8c=)�7����P Y���A�JɈ���QfdCELi�7���*�X5�Hv��{Z��[YS���68Z�<�>56DX�c9b�@�F�˷��F���:�4���/6"��R5�tP�^��i�&
�O��x�� ���K1 @O�C���؈��^;�������h�:¿r���&a�|�$�1ҩS�`��t�Ob<��8ӧ�N�YW[i$&��d]�JX�ˠX҄m"b��aJxx���o ��C��Xk� ��t����.^��A��q��\+7�''MQ�mѳhTk�I�q�J)�dbq4f�E:���ۺ������ϼ�D:lg!iRp$(n�DO������b=*�cIc'�p�0��9s[��������w��bT|M1D���i^ bykv+:s8B����թ��;VX_<��U�P[^f�z3��%��(�Ć4<'#�i�z���x|�b�C��2Kt�&EN}�~{���ncsFڪb����矉���	c���D��sjC���q�)'r�S��Q��XÓ��pA�|D/�]�Ua�8�9�U�D�3�h��q|?��c*'
UÞ�������6o݆��0|
�!+a��f�@���x��J�L���vTڲv��hni���Ɠ�8�k��ҷ�ilj�(�W��iT<D	NEID8�Rá�9^%*�����ǞG1$�6i)Q}����L<:� ��11n}�j�JRɴ��w�K?b��4��4|�0��P�V\�5��\&��Ն5�	��d��D�#04=��}���_�9Ry�,���1G�XE9��#=��Pm�q�aF�-����02�㌴�Ʃ�ѩ��Dy5��1�>�e�c�Y����ϢSO�4.��m�v�z�{MAʤ�h��r�/V��P/��5#�ƣ�N!�8�0�~��sC*���R�seB9
���#� Mv�2F�Vr$�G�������|�����t&z��聢v�5-����$$"s-觫7�X�'4��c��9�7m".���z8���}���1�C7�����������k��bw`���-+"�b�����0��0L���?��\����c_�3w>�w��zl�o�M��j������@KK�wy�-��n-�&d�\r�O<�(�nj�x����,��(��ȃ�նuj�3u_|��/��^�oi)�;K�p�&{}:'���!��H/>9!�m܂��
1�g�x>������%H��K�F��u���9ϼ��xb�Q����op��S��ю{�݊g�{]	�iP}��;Nx�!��ذqk^�X��zy��9���G(޲k�G2�}'��A�Fi�xP����ft*u�Gۛ;z��BV�w�g�z>��s�ɜeQ�{�E�K,�%kk�Ƭ�6k�֛r�]�n����݂�/9/��H���Z�I�
�'��h�ve���rqAS�1м���6�`7�s�қ�"��/9�`���d��<aY{�2��۰����8� ֵ�7b��q*��{4*pز�^B�,���>v̒�o����e�٘Ǣ��WU�z;p��gc��ߡ��%�x�?�Jě�K�U�X"�6�\�!���|��釋?���BP���x�w�g�5�W^V�k�\/azD�y��%x{�3������ �?� /��4�[v`�*�0���z%���V[��H��[g�t$>Z�	�eI ��eN;�H���*׷����ܬ������%�࣯p�?�`gc#N8�P|��Oؙ���AEY�|��HE��k���㫏�Q>�y�X��6o�Y.pyN�۾�i՟H��ls�1�blU	:�B�K��Wނ�bh��˪C9w�� n��z��ڀ3�;߯]�M[��W��%:�F{����_V*��I��C���y�;�L�d!'�.�.z�*�A?F�{�4
$��h���	���d�0�va��Kqꉇ�i�F\=k>���6}rxp��b��O�vh����;�ŋ��\	E\��G��+.AOC#j�>r�MvE�A�.=�Ӯ��c�ee��G� ��/���NC��#ų�q�1�&��9����_�S��ƃş}��)C(��+aC(â��'��ߗ����7��G�[uv�]m��ų��ր5�����q���o��_\x�����*L^�C��WɊ�GKֲ��6�+H����_u8�Q��C ����2#F��oq��[�E��!ho�K�<�����XQ���|�����r=�������K�,��̓�����$��dW�"N����ÏTB!g6��K+�����E����ƉG,��VC�h"��g��vm����K＋A�,���IB�f���>�
�O=�M(
�ڰ�ʋ�
������K��v�f|�l��QP��1	�z�<|�u��#�݌��>HP��(�Y�m�^��1	�<� ���;ZεM���$Բa��	:�C7_+h$���}���m�C�b��Qx�g%�wK���P��1_�7�p;�M�A�۟±��g1�cAi*�*�g�w��b�t�,��5��[nĖ5�jo�/��G�����J��<rB�no!�w7n��D��p�!����d�/�����a�Ckj0����)�V�:��r��㯾�g'p���}�D���ؾ�O47v��������!n\b�� 
��'��\��+��ā{�9'/gي]�uR	��Ak���C�r)r��E�$9��5��Y�ē�����'j�Ӡ��]�5�8 ���}��a�u�ưB�O�T���?�'"�n�Ǳ�qcF����M�Q��aԈQ��gQ(��	-ͽЎ0{%�>��`ޝ�޴��\�%N��Aڝ�����?���G����r�(��x��/�����[��>1X��~}bx�G'2K+���M[�ܺj�Ⱥ�r���ݳI���[���y6v���A�(+��Ukj�DO8!F�W��ԁl&1m�� �`���G�~�ߔ�/)��OP��-0��t��_E�l�R�b��l��~Y�
յ尦��cï�A+�*+%N�PO<Ƈ�(�ژgUîj|l���u��7��E3NEF�_�W�h726�����K�0�j"�Р͉�g���o��k�>[��d)�Yʆ�hD� ��=�l�r16C�T;��:���_}��MVժ�{ɸNm]ve��a��F|��G��:F��Vc��_X,��	7�����|�n�G�=�p�b<�+�P����
���"�#2}`��o�UJ��rֺv�iz@P�S��#��}x��'f���e�!	ռbR�ٮ�yw܏瞸��DI�(x�� �89v��sO?�itZv��ڈBs�|��XQ�8/��Pu�5q$�\�b����o���������7	ds*�dG'�g{�}�+G�`�U����{l��[�T����.Y;v��!F�O��K�I>��[���$)Q��Ɉ�V$L�3��V��O�R��Q���Jr����X��U.p����!l���'$��8���[q���5KMn^lG���lmڈ�+���jҜ�͏�g�{���2h����_q����$d-��`9Q v8���yI.K���2�"�Ψ�vN+��cp�3/��CDͰ*AaA�2t��+�%_-U��l�=�/pj�F�U��a~�]L�oFa�T~�iOF/�u��uK�@m2�KHe7�M�,~1�	�$���?����S�6��#�ղ!M�}#0���\���\��)cP���fg���{�y�qp���A�\DI�9Y���/�.����� �1?�lP�ɻ~�ӏ: ��K��p�<�]B�n�����2����QɌ	b~?�a-a۱x�2Y�CQ�sk�CB.밚�X���|��$�QU5h�|vc�@<��/�a���v�l�p%�DcZ������@�\vBE*�4	��$x*�Ưl�@8�����]�����c�z�Z���7��^�P98���
s��U5n
���.�<wJ
��z���B�k���'PP5T��%>����\��U����G�J9��5��棉�2�'�n�����%�**R���c��Ysymf��Ko��n�F9m�4�$��$����;�[`��a��*1eb���T
4���״�f�4�Ʋ�^��{�Df�/��U��T�)q�\�M[�+�*��,{��-Q�@c���ӯ�Gmu����6��]�dVX������fP�ÀU,7���#�r��&��;���mbH����0e��a<gr��k�Al�Ig��tN��CBƯz�r���t��B�"���rP}��@�2a�BQ9�m��O�r���9k�����Ͼ_!��3��`R� rxT�ڢ#�����Nt��Qy��8|A�Z_������eJ`T�_�W��Ps��F�r0��r:������V�[CH�g��>g6KJ��ln�Q&���JNH�!�O���ԁ��V>J:Co�����:��P�*&@��X�/~�C'K�?�Q�
�^\�TCj:�W+�V�6U��k���|�H�W����B�p�)��1S���8�&�[�iI�ϼ���s���}f"�ȍT�"e	�k�5{�D�Nj�y�а��z�y�[6?r�lb������o�;?���=��L���_]��V�[s�:ImI���RY���A0�:;Dy��px�����f��x-7&}�8���"��8�d�y�(���@q!�}�e��rd��	���8/�XW��͠�7Y��Ӂ.�ļ��ص	����.�*��݅����T��j����H�f���1	��{@#ń��]�!e1��ߢ�z��@�X����:lf�� 7�W��42y��ϰ8��S�!c�d�r��D��ŞM�d����\Rf�Ĩ�X�Q���;5d`��b���f�1�'�!7��9wa��yd�͜�NYhos.&�1mkS�#�P{*�Y1�Μ&Ȓ�b�w� Iai�ѣ��J5gџ�ӫ+{!�95�Ғ���i_����~2�sT���=D
&��0K�h��U`6�,q����h;s�0���I��������tyI@�KǴ����6�貆d�j�A�ï�90x[��/�L��~������F3V�0PʦN; o����,�=X�,%g������٘���ye�"8����&-�;�~�d?u��a�Ϧ]����`1)��`��$D� �P������v�C��y)��9��s������l�w`; �-\%���Y=�9&pM4����*F�j8��aLStrH0;���xs��|V�ct4?o@�2����>��f-)�����SAJw��qCI�Bh�n�t�/dapRd>��"9}.�j��ش��XՓ��{F��)6%�k��)�(�0��i������񈼞,����'#�G^�ڙh�Lг�"����o��l�6
y�=�ѕ��lMv��ǵm�ӵ��rl�&�1�f���w`U��}:�FC(�Mn�İ��~UNc�M.4{Xj���g ��h�%�����1�b���A��ԉ0.�fQ�x$/ۺ��A��T\�K�����S� �-�;��|�_	�������sK���i��g�D��L\S6%e)j}^NCK�U!�٘B�[:�F~mw&?�ٖ=D0�1t���!g�/:��#/i@|�ׄ{�c�D��A೦��<�Qƨ��b*OɮˤŬܶ&������AR��U9P�5ʨ\���ukY5k�+�:®9�T�����h�A8%T�a%�"�_ָ��R�����tH7�w�3�����1�|�]�4x�u��˳�2��Y�Qq�j2�r�6=��B�uJ$d�4f��4����)z��2&%|2�SF�U�Ť%��uT��4%��'�&*�j����R�{q2�A��=q��3�P�O�p�@<:Ɉ��9=PVeqb�Xl ���$+l��d�����s�z���?�2#!��IQ2i�-n]ؤv)҈d��`;��#mǡyX�k�'Y#UyaTP�d���F�K��a�s?��b9�Fb�Cy�@	��>�Lg��P6*z����6/�1��������(��2�,�&������1k��m�b�AY/�6z�(����z���.�� {��'����ϷK����#13zj�(���զ�!��A2;e�":m��R���vT����$�3cxU��Is�F(�VFC3��A�h����j�ߗ�Q]]-�a7Z[��,��ؑ�!��a��@	�Fl�Ps��S���TS&
a@ �Q#̡{��TS><3��3*�I���ELIs$�E�����6��`@����Ǎ����5ZZ��
EEt&�$�K}SL)�'&ap.iL}��)C��V��{�q��gj(��%>+?/[f��1����O^�L����6�c�8ÇԢ��A6�ɻ��rX�b܁��X�!E� T��iYّK�Pۅ3/�S~�Ҳr���ڛ�RU(L�J#Dcd�# �CA�^p��ړ�إ�ͅW�ƶ��a=��i��^ҩsQ�4�,?\�),�)��x#-����ѪE��q�!�c�葈r�@�K rJ<\SK���J��Phy�^4cxxznr�Y�ʋ�c ��!fˎ�-xlט�}�E��A�pw.�x����"�Ooc�.�R�،忮�XΑW�N�?q$��f�6|b�V��-3�-�Z}��Z����!��z�wb�8l�ڞ���	<Do)q>G���ᔋI$�r��4`1w����#��P�_/�数G5n��:#�|{95�~�{@~V����g��!�P��lV��ؗ����D�R��z��K��t�8�CQ�s�;�˾�WVb��ߩ'��w?�^�*�Y�IӲ -��1���N��쥥���lǈ�F�u�,��wljhV�o�_�������ܣ��)G���vMx�3���<�`?�`<�������Wn��J�m��g���+Ʀ]s$QAi��9`߉X����h����Dfq�<P�k���G��3i�x�Jt{�̑S1��/�]R�Ҥ6�)�1HT��Ӟ�U�_-���}%�roo�V���r1�y�m��2B�����Q��ű6̜~2F֖)2-V���A۵�>���/�H�����-"{�����R�aݟk1~���q1���}���c���y��4�c���LY�������;�r�ل��:%�m�yga�GK`�wR`֖����.�v�Uxp���-i�WO�﯈X�3O=��#p��$�7���C+�p��S����p�}
�5���|$�"���3N/�)��G�Do8�d(��
���ş/Մk��%󞜂٠��w������Ҧ�nUbI;�k�aP<e��1�\�$^��WNC�>9�D�:P� *
+u���S���x�d�Y�c�s�j�O9�A��L6t��8��CQ�kCY*A,$�_�*�g	�p��}PWߠ��+���Z�P�̲3Ԅ���ۅ���QS(���KB����H��\�S�������m�yW^v�;Z���5u�ˁ��2l޼YT�/������K+��yyY=��ٽ���7�T.3������ء�藽����p�cO���D���a+"�zz�#=#jʐK��'�B���
Ƈ%i����A���v�Ԧ�wrF�Ŧ�L
'�z���!M�8:$d���3 �<,@	���þ��s9�Ճ3�?N����-(- �s�1�.X͛~����+�;�A0�"�*Q�p��8{�ihoځ�G.�[�� 99��.`���W]�{Y�����$�\�::2n�v�\x�e��}�s'd~������;ճh͓E�h�lQ]:s�����������F:�wH���^$F�Cx>#?�j����Y��暹ʖ����GF����̺��.���<�p�(-�F.n�5��{�;���w#-g�v�h���hmlBUq�:�l	]�q�ɰ���J���-��ա���p;.�y.��=�5eB��Aq����:|�(�;��')1SEE��ƃ�A�wu"&a���z���m�����0"�醫/EH�C>�5#zU�;�M�r�&�8}x������QU(��γ��jn�՗^(зC��@3�_��.���$c�l��DOo�RէT�У*Q	A��x�l��(�$PVT*�+��[�ḓO�򟿂��u�\���>�5{Ū�w�orā�1���dX�׊�D�!�)��4��^�u�a�p�wH�
�����pMi!��۵[ �C׏*��v6a���PW�eY���P.�w�nA@�8���+��p��P�N�{Q5�h��a�	){�P�����C0������/�+-�^��b�P.�q,��>�,�������-�#(,(D����f<t�\<���0�;$�ؓ��ô�GcRu������)V��Jˍ���D��0~$�Z�Y�6��)��)g���9	&	��ሲ|��B�mm��Qcм}+���ܷ�_x�Z��6�����w��]�ހ~���b�'N�_}�-���B��L�1���~�9�b<��kpx�$�J�/�^��R8r�\�>�k�~��=����M��/��7��R���Ͻ��E�r�̚��7�vANy&�Gx���.�P�)�&"��� ��o��LֱZ�JFèL4��� �S�x	�p֬�Ѿ�WB&�;�Ϛ	�)�}'���}^x���yb��3�Wq內�Uَ�.�Ǖ�t���[�^�����u�H���O⒫�TV"km7�][���<��f61���3�שq�_:�a|��ny�9*'���uw/V�X&]<DefL?UD�t�y8~\�R��2r1X�>|���ز���/xO,YT+%Gy�j�R�0X��������be�U��^�1(ErJ��⭅�����p�?.��1m�͎�%�z�z�:�@��뮜�3qY��{�{�~;�ש�,$�!�2	�%�ӎ;���@� B�8\�p�7Y���)�M .��#�>�X���f��p)n�{�2���v���������0��e�Ϩar��0 0���
�����!�s�Qb48���z��gM�+���iS�����h���z�r��P/��0�3NBI֊��bT����MM�P��y+g^4C�L�x?F�3ϻEb��$��a쇣�O=R� �aÇi��:��c��,)@gG/ʇ����~�V��a<�?y�;�Mv��a��s�p�7�%p�ZL�K�̠�jn��	4�`R�5��~�$A�P������VAL�3an��s/���-��������7����"{]6z��8m�Q����ų�8~<61���(���CO�\|����Ϝ�b�*le�D]K�L���	��ss���0��w��/ԲvW[���/��B\qͽ�u	Em�̵������M�\����ܩ���0���4����4��.�n1^s�:E%>}����b����ܥm�}=������s���k����}��$k���t8N={�|Jj�*����U7އ�3_{J&H8\^Z���]&���?�j؜Y�?��~���
m�g|@RdV��|�y<��honĝ��Ͼ���������gIH�-c"μ�
���:X�0�tؓ�=�^x�qX�on���V�����j]G#�nx��v\���6[v
f�F����L8FNǪ�7৕k�by �����i��c1moA-a�=i<V�� �ܣ#Յ��hllqy��G�b��p����DD��s�y�n�F΢�)�(� �@�z�x�<��N����At%�{ʦ�I+.�i	)n��2�dQ��J��yg���ʋ,?�-�+�FaE�y��?1�a��DV��7��;oF���j�ur���.Ñ�vv�'2a���!��A$-N����o	ܜ�"/�&=�oKh�%���Ws4=�-,����y���0�$����}�G�I��[�Q?~/BQcr�y� e�f��_v�m�"��Șȭ��k6o���W�DW�����.�;�3�YC�U�U9d^|g�lo�]K�$,�mk3�޵8�詚��HB�G�yxɭB�g��蕵���49l��,g���aʾ�/и��P�~|�L{L���s7z��q��W�Q���1	�T�ε[v`��Q(�Y�)�w��MbX���TUh9��	��_���Lb{��v&~ch�0����䙉ʥe%&g��K�[�D/�b��w`0%�΄4A3� ��;��+\t�����y�f=G)	���Ə��9'����R�c09�p��������G�����}L�NOR��d�j�T���;�\��fN�0|��8|��E��ǣ$X���rl��2��h����ar�Tyo0M*A��p�I��+2K(���#Q���Ҧ�*��v������b�J�{�Espʺ�X�`��'�	�[�6��ڒf�����/��0/�!���YZ�ړ��O*W���x���j���� ����5��'�n��|f	��Р��<���~��.;b���PW�@;�셴}����X�t}�}ho놫ʯ9*��.t����މ�ؠ</�Y�>Yw
�i[#�2�X�&���4S��?��^r|��r�2���N���eXދ�Nf�c���e3����-�d�>��қ�OkVy������W�ʋ�4f������$�h�b+J��G_�%O�b��߄|UΊ��v�;u��,��-}����l��F�o�KH����%�I9��Z�w�B���j���g2�[8�C����/��}$#5[c/Z�:�p1,J,N�/�נd���29d?��y����)q6QMDS��_\.c&��|�JS��"gp�����;�\NQ�Og>X�d��j7�>��A���)��8�v��$&%�)$�����"�)e�r[sRc�ߖ-[1m���,GU�2����P�SU��o���"�K��9�N�V�!��[!F}��iY-pZ�j$B��o��
Oa@Bd�ʙ���,��M�f,�a3�@R6j���9�h�lt^�CU�8��镐4������%غ�N�©�Dو�aZ2O������r�����ήe%KP�M��'�LW�f�g�T���/pO�J��\�Gj����G�D<�_ɚy<V�
��>�I"���r��;Ki���j�����]IwRTM��N4<.��4>���Zy��3Zڳ�mJ��r=_Mu���7�~��}r0�������.m&�ƍ�-v���u�y�kU��EUm�Lr ��o�֭�K�lK�yt1d��t]gg�!f�5��3*C@c�g�*�u
�h��(��tŪ��A=��py�JDd9M*d��䴏c�IEYBU*��dn�M���O.zX������$Y�R���<�n�j����I�A���Ŗ���b�P�����l��w j��٪�"� $���� }1�3�$J�d"f����s����٥�����M���,�m�!ve�&+�C� �~A)C�ʴ;����1������1�I2g�y}C H�1��5��=]�2 B�4��X�56`w�.(�D�l(�S�Hޱ�Ч3|�~YOδ�Q\1�䠟��uii	�bEIHÄ'�;��:�RAa,�aM���ƼM�[�ϊ�|v��Pƃ��u�n(�y�N��Զ�j���l��S��F��!Țƨ�$�w�Tf��MY%�����B^|�$+�QEb�<!�F%b	�<AE�oQ(��%���{k��W���.��)(0��'$���]�].��}O��~�c&}����>�
�75k%*Mb�TV��$q9l4R��v�HH	�j�!�%�TT��1���bw�@69 	�d��Pk#eBL.=����R�9ZAfs=.�da(Y��H��Z6ͦ���"��e$����$�M*0ZV��V"���WoH��Cڬ6��T���!K��ݗ�9ɼ].�S����5M]��ȑ��pZKF�x�hƁ1N�x�m�vC�N�?�)^�"�p����4����/S,��K�Z���'r��>Y،6�T	\��y��y�W��UQ��`!�ڣ����j��l�4��)1�	�>�e���v>�P�+��ÑվJ6�5� �0�Fޚ�`J%4���nMi˸�	�(�ވ�d�ݫ��ɥh���
�X��*�#��A�ṔSI{K��ѩ$�b���s;��#��`Sv\�tw����ֆ�Z)�ͭ�q���0z��MS���r���\'Q�G�a��{����!��eAEM�6��׃(�)F�*���Հ8�,n��W�DlknC(�Vb�w�`hm�s�8B�?���I� R&D#I�XI�{�Yx�W�+���a��dc;x�(1�vt���
i/R��'r�Y����$���)h�Y�?��}f9�>1_�8���NA����L��dM[ZZ��T����8l��h��	}m��i��N�I��qԌ��;u��w@����IcƬ��mJ⌓�ۋ�j�0�Ug��7_=G�[J�W%��P��I:���ug�|��va��6	C�ؽ�7]�r�Zww���}�eS�cd,ʖ|��G*����d��b6�`Y��w%�s�}Zڪ�MmnnV�.�@���:A�W�dS<^B���2{qо�R�5�6�@��q�	A
���Wc̘1���)1���Q<b�\t�6K)#�\�!U��j�������69�Lk6�Ȉ!m�e �Dca����>q�4ly��4�ɡ06���KϞ��8�n�6��?�������Ȓ�bX���{�ݒ��N�0#GEww�r\x}�0�<2�1,��"TW>ٌ߮�ɯ�ڌ�����V``�v		|*� W�h�a#�<)�)?pܑa�?�)�S��	bʱϘ�r9�Z�]�~�:��
Y��Є)C
���U�1�,|��/�ZI��p��=�ʲ�>+ߝ�jt���KTj�����Ι��Y��#a^nK
eA7&���D ��xa�V;墧S�O�����ϲ�($Z�IPVǜ.	!�C������(�ʁ��Ҭݭ��a�<���#�',�^ySBM��v�L1G�qάt=	�)����+P��Sj��ˡ�r0֏SN���֩�� �bQ%T�8�Z��ذ��R7��9+u<��Ԡ�nΝ~:�X�^���I!u��.:�L	3�e-���u/�����P"ݽ�|Fݟ��S�_|�R�Wi�WD�>�<;�*�ʌn	�@��MN����H8[ļ�n�7_|�>i�6T���5�M���"l��O�_D�9�l��wLs�$�1t8��s>��3�
"9���p���"��H蚂��c�â%�	/�� ĵ���15˃����s8�zɩðq�Fz$v5l��3���?Be����nڅ��ESm�	D�e�r�,��S�a�V��.�c������'b]�%%��jW3�:o:�v5�����_b*1l��AlK��G_|s��u�p��#���k�YmZ����?�FK���BY�\,n0<�}�f�A�01%��K/������%%����a�X^L#�*�{,Q�0ޒ�˖�~lh�Kč����xfO��J�B�P[\�c������X(����iYzo"�>�GM=��.̻�,,\��w6��'r�q��{�F9P���E�
GƦ^%���g���w݊��`dM�n���[�L2i�8L;L��.��,������pzj���32a��E����L<�Գ�J���<v�~��8���/�P.,g!��8��\�_�m�~{���W��kgc���&m�!bt�aBŷ��Z,Z�&�O�a�D������Λ�O��~�������{L֪C&��r���;���_�]P������؍1#��u��?qǜ����QAL 21���O7�9�w�{�@����Y%���E̐}�2���NmM��ƌ�AW{�:��������!iM�?�W_:�r���W��k���%:�PS6D��,��._^z�u8|�L�1MX��G���#�FF�>�8���wz�ikz�C��#����{�<MbH��.:p�����?/��ٯ�oS� .h!H
��AD��2���-���/�a�͐N��f+�y4i,��b\l8�Ô3����%�qȹ��2�4�Rl�\��@���ƠH Pc���G�zF&���b6Ƕ��X���R�Do�;�٠ V%��lASS
�ʱ��:t�	�qs ��O,a�������L�.�l,���>>�bR`)v���v��|��P�Ru7��ۼX���8b�A�65��:��g����U_/�#��X~֋(���|�}�y
y��.��v��^Ay���34��8����QQ=���v�1��9�r��_0㔓䢬�-7\��ͻ��ݏ��S���Uo�<g�h�NX$��F,{9[;�] �ı#���	2�䂳Ѳ�]����!�߷4���jxR[�M��n���{����GR���_��g��x=5{��Jx��bL�ej0��4��8���0����։�ؖy���3#��y�6���d֎_~[���	O�K2�!�l��6A y�!�퐟+v��}�ku�y+���\>|��4��r�ٿ,�V���O����\�?W~�QeV�x��:�W�m����v8�i-x��TV#���%�2�i.��kL?�48d]w�# 0i4�B������T���}O%:)R�R?�"�q/�cu����P�c���bX��Uڸ�^� <w�~ߤ<0�����j�^iy�������J�t�o�p�c�/����ڌH�Y9d8���.]CFq:,�@<Gw�^�#�M;.	�v�ߤ9�E�RiQ(d�zï�g�����fY�ܲ#�N�����ӏ��`<
� a/��G��cxM�����X�ɗ��fՇg����R,Y��;
�nx0�mo�1�FC	H�����rr@�1�2��m}���E�K�,��*�,���L�P�ᇕ���;0a�P��>Է6�C��4;W��l����k*Pg4��.���K�ƕ_(�m7�w5`��Y�%��b�����o�<U��H�\�,i�x1�DA���&�iݱ%�2��~�F����b�~�2u���H=�}<m��/~�駝�
X=m��¿gc���_�f�IX���Y�)�>H�苯1���Q��	STB=D���iǠ�5�6��"G�>z�R��4;X�N/~^󧎰��x12�hشI{;�����X؎ϗ��K#U���f�4��P���"�t�M"��Z���4��b�����j�����5?��(�]P����s.<O�i?����
�%�H�����^Aa��0UZVW8�'����[�<^��0�w*/+9D}�
�]���:`w4L��bvĲ�B���j(��:��:l�s��Vtut�{(U]�/��9&&��͞�lL.�G�Ӓ/����ӮI&�9�Y������㯿AL���:jVFw�PVR=���%�\t�R:�Li����C[Y��=~��}0�b;=��ل�j	^x�m�s�튮�b��97ӟB@P�U���O<�����#dSʨ�f��&���)���*\|޹���g�fU6!"����+�i[�^x�萤*��4_VR3�z�I̻�J�sFC#VT�1�:A�-�X��<�^̳��)'�9�]��� /�dj�K�����t��jX��>�s�}d��D�r1^��;�}ExK��Y���FDf��B7���9߭�]% ǎ�կ�%PRld�W��;V��>��,G�uJ5���^(�#�><��[8��㕍�P,~�c�n���c��-���F���ҋb( 묬l��6nCg� &O#��@ii� �^��>���7�$4����Y��#��*�fu����0rXJ���<*|�д;ۺ�#D)�3��bM�f��"��HA��A��7�Ҡ�]mjLȚ�ھݡ���d�ݩc�9EeL���Sh�n�L�8YB�]����5���G,�OP�!8��p&�t���N��4��=�.W61����R��<�:���thД���ޤL�6��y_|�}A��ɥ#C���D������Z y<�*�����πA���a��N��)A�}��ա�[&[#�����&E�����(�rWR����{����B5V�eZ�$�[���i:[�������� M���Ձ�o�Ζv��M�Z�͂�
�i�6�i(��|v^8M�C�::)�-~�o˥O�{2��s�ή���耗�ј�Q4)׶��
����0f$�nى{�Ę��u�4,�F	U�8�opT�t���%JW�l���O.��e�ِ/�Θ�|�ɍWps�S$�
 1��3��w>��^a�����ɺp�������6���]�e� �E�\6��,�Ig�6Mr�X�����33�Nf(6�Xăy���Ƅ�)O�<�,M���	�^�u�VH�QjΈ���W(���	O��!/��Ub�z��>��dR�X�O�2�TȈS�V2�f�(Λ���g)�&���7��~�Sbθ��F�K���i�?� �ӱv��s
X�*[�ug��?��D:�]tv�_If���?�����*SV�~�5�W6.���!��ap�BgoLF�:�'p���I��I��65��$�
���<~�a��NX�7��e�F�O��D}G�1��
K��G��*Y۔��`6�E1�˯�rt����a	���u���iרu��r@����0��)��"3�,��J�s`����g<�6���&.��j]	^@Y�����1�?uu۵D2���[�m-{9�.�F�(P�2�|�Ϡ7�dq�lq�Mj�uh�b7�JM�"p.�b��2�fS��jѸ9�"Ҭ�<K������l~ RY�Ām�s�e�6exr�0<geʤt�T}~xR�JY�wB���_ɚ���*��O��6;�e�z�ւ=�DU&kJ�Ǭz9Vx�lA�A�,���y
U�K�]��g5?��0T�u]�{@�������S"��euU3���Ua�,ZRW�9yQ��*;���:�1^�����M�P#hOJ&������iTttژ1>C��9��z�����@�-׶��bX��Y�h���ZG�"��l���t�un�����})�y/��|^ :>�Ʋ�ckS��"��Ăi�����a�k�R:k1������	�rd����d����Ã��&s�r��|)��ANs�06��tkӆu�!4.�C�L���$��r8,��a�?���4P�g]Wn�/�Xs��=�y@�v��YeG�4��ޕ�9S&ox2z����I�7�,��RD���1��|&�C�c���r�26�1���"T3��h�܃�����j�j�e�_F#F�Y~�1̸X)�y�JC<��쬱��*����_�2�G�� ��=c�s�A��ܞ�ϓ�!5R�wq���Q�c�Yi$���M�u��)tU2zw4B�wR��<���[شڴ���?25̃���eK��y��I�����VZ�٠d�2����E6����9.�)���e)\{�l�Ġ��R�9�+���J�xdY"���sa� �³��!�㸰,�6Bq�I�1�:��l��zMLJ��^>�BH�V�ȀzY�p�m:	�SBc=�$��ò���8AƈyN9-���R���A�?��D�;���J�U��j��ƢZp�Sʂ'��(yI��(���SȲg� b�Avn�"������\l���9�3<_T6�n��SNH�U��LQvyV��|�Kk6ɴ�����B�_D.N"��q�Tʸ0d<#τ��Z��l ]�sյj�d���1��nUf6v�:��aR�hU���9�΀+�I�gp�IE���^^�Bi�*u:�DL�&�T��t�+��ߣLW�r�8�ap�R>��� 9c��˦�:1bp
��]���JF�s�cqA{�x���3yHo�'0i4H(�~U���I%��Y����C_�&�)���3ر�΄�_{�S~������Ĺ�ք�{��¦,m���gY�A͹���abѐ�����4�\�,�+I��?:�����p�r_)t�P���Z{�|nC����KE�<���mNG������s߄#��%t�z�J0M�`�woljV�Ik�-���CeV`jL6?~�m+J*���!� �M�R��V+U�B;�P/&O��hz(f�m����/��֦|�H��xrQsf�z��M�0�F5��b,��a�+T]�<�:����Ye��9ډ1#k0e�aH��H�B�z";�nS3I��nv�of���v�0Y�� �q���kq�I���^�h*��W�Ǻ�;�s�T��I)��$ĉ�g�&"1�8���P"��q'Ə���xmx��P6lR<�T�d�(6)���ܹ��:W.LVG�y�yfAN/����J��;90��+����l̠sw'�8����T�"�=��\��͛�ê_�,�CD��DD�Ia�1�p7?GO=�~m����#"F�Ͽ�5Xh��ё͉;��Cc��,��I�[������k�#%1�Gb�/���1�J��RH�Qa������W_|��(%�l�@������Y\��ě����j1��� j�+12mq1�r�����u�t��w�ܠ��4r� ��<��eH�yjb�&;)�9�&ӱ~\z���T4I�^���>A��X��W�)�L�I%�������ц�>�#���鳣/���\6�{�|T���,�D��l\�R�$�2m���-^��g�t����j��{��a���b�>�_&˳��;��L��1���e������i�����z�aT�-�lL��;K4jhnގg<[�C�uJ�+��E�+�����uƙ' L\��� ��~����Y��R6\�'�Z�<�g9�l�ӏ>�]��*��Y�>��������GD%cC��+�n$v�ŕ�g���dS�l�9����#'��'����F�/��ٔ�x�Y_�p�;	���H��,��Ρ�̫�����p�W�hG�E����FZ�ɣ���`���@P�0�OA�QÆ�@c[��"G�0jN1�l�noż�"�E'V���?Ы�F�r�n��Z<��T�WrW:4�� ��x������y� 3@�+�;�0q�x�ni�ŵW]��x��
#T"�$�$�|e>�x�4T�ɻ��*[TH��#�(��������u�qK�NN�)��c)A�Ua�>{+K�sڻ�Q)�*,��=�q�iZ��2�H\�;�j�IJ�d�-�����P�n����nt��[<{mn��Y����u9��A7�;p��1����u�1����ކʪ}��5e��Q�c�ʵ�\��s�S0�Y%�� �C�?=�ʳ�<���bA��p߼[q�-��|�0�)�ZʤeWΒ�b��GyI)ښ���staTH��Y�����{Q.�U���(�!��.�ɲq�/���ݝ`krh &�݆�|�o�#GO��vk��,V����޳̻Q�?j�3^�ĺ;;�I��.�C^V���i�Y�IQ�j���ĳ��/Ϟ@Uu��,mxP[Q��������a����+��ip���F���V<p��(��i������p1IG�ԃ�kD�kww?*)&lgw��MQ��S��G��H�U�pi��rica� ���PY��Q�l>�ݓ�6ӏ?�}�����V�+�e���[1�3��8�J���P;��� *V������2J��!錨���){c�xj�1S	eS�݁�N��t幘�����8|D��Ҝ�)��X����*�C��Q!_Q��6KD�p��S���_�vs\��������!�khk�*�����J�X�+�.9Dnq�-�q����yA��*�z���v�ۯ��إ��e5���zWG�V�\L�nۈ��Q��Y��!T�)�����#�ʥ���M��q���
�3�	$-)���C��~��Z��3F�.�T$��N����� %Ϊ8	�$�I���K�@5���ϼ����i[�8�l�����
yF+��%�rص����׹W�>_�}av�RĘ�{��=����wf4�%&|� ����UlUq&�����u�AȂ�zz:1�� ��8;(�Eqi�\��yy���DdOi��y��j��n�a��C��sf]��1
�c�����pU�����I�{�uW��Ǟ�͉���k�ZE�zq�	�Ț;��N>o<�:Z[wc��!�k�H	���(��3�����!�ذ+5:У���<rv	�2f�?>��հ��ç��C_o��F<��h��FA��s��u�V�}�M�h�ia̎~D��*)1e:�JH�ϹW������JEkj�����K�N������ڕ+�i�f	���᐀e1�99Pŕl�҈���2YImM�Q#�r�����U�<���P�]��嗜/�e�&����C�(����q#�j�����9/��И�u2��T�8Zn�èQ�2}���\�_��T�a�ӔFnxE1��r��~�@C�,vd
�?z�<IմYt�����U��؄�`�w,(���֦t��yQB��8-��A:��c�!�(���/�`��M�$��c��� ^�c�Rf��a��$b��5��d����.xE�ry9`
�o/��!ͷ�8�$|��r��^-o�����@�x���j��;z
-�mʆ>^µ�O>Ve:[�q�E�♗��RFs"����K
��Q6dz�y��yei���L����X��!�N�KQ�k�0��tp.�+f]�m;1j��x��f�z����~��f`w�V1�\|��X�ŷ�s�6�0%g���O[��;����"�����\8�hX�?�4��p�Α�#�,��S$�H��5{���/���M���.�s�v&�:���{7�wk���R<��*?Q3l4�{�}1,[�B[����7�J�Ǒ�p��{7n��AK�5�L��d�.���e�~�m,_�Zg<��c�Źg�}'�A��{�w=����(���cGa�{����v�LmcNk��:X���>{��qWΞ��>� g�J�q��C*2���8e�%(��D2�F[_����~߈��}r�^2w>��n�NӦ�q\z�lx�(�Lj����s���8肀5�<vϭ��{����]�ş}kd�dhǍ�PBB�@	f�>]Ѡ�9�lo��n��
\��ٲ��z_�@�%_��3N>�0^{C�J���z�$>����){	��lp��_�����B�y�*^�������m8���x��9�
8�(�=U.Uss���X���;v��(��.�H{�<�����*��.�ЮD�x�DdPE���rr�J��`��m�R�7����O��;o� ?MP����/�U�?&��b�J���K����� �d�H�d�r�yX>���^�C���Pb4���Uvr2aO�� �1����
�s�9|��2��4�)	�UU�q("�:f�M����x�ꑸ����x
�+(݆҄�6�}�D.�Y,�k;��;K���uH

�)� ҹ�CG��=�8IwMD㲆���_.���Xir�j���])Fm�SY���f�`!n�����WYn$YŨ��рO�~�c�GsV�&��\�J�`2�MŘ�Z���/���
.q8����Q��_2S|ݠ��tG�6�X��>1�#5�2q�4�b�<Z���<��Ë�p���R�Q`����SϽ�*��`�VRY�;z�:
��Ꞅ!�Zzp��O��/78"�I� Zb20.�9tH5:�}��;ll�wQP��=�����_��1r$
��vu`��4v��OLP���Ir�5q"N<�R��t���������FJ�F� yA���v��۱�8��W݁*1~)�ʙg����[���o`�1C%�6�g{oX�3&Nc��F����ĉ��A�b��=��������O�F9>�C����X�u�T²��h5c'b֌Yr���;/�V&�⩧^�/-���u[�a{5�*�&u>�b)N>�D��$�����^i[e�+x��>ĳQ����O���W.��D�ž����݃H�V}�I�mŚ].	z�+p��/���ި!E@Ά+6�����������3l�ׁ�@�ZY���'��waG[��0��
�/�����⺹�a�$�����V���D-��)q��o?oi��cx8�e3�b��z�v(�n�=��7c�	�z[6]y���WT�f:� ��p��#9����T�>U�2Y�4�X(���/9*-���.G��*,����@FJ��A���Td��{ =���d�����Y	ƶ�li�D���-u8hl�zbo�O�،��ˀ��Q�)�aW\�eZz��a#��͹��JJp�#��9U�g�8k��'J9q�lT�ġ�e���dBf444��,�n���2��;5W�Ib��3I�򷍂f�Z%�>�?�ܰs�������DS�N5��*y��迉��[%������`Bg[��"%{�\�H�\�Z��B��ʜ��D%L���H�l�f��p'������b����^(y�Q����QYH��{<�r�]LcP.5sѬ�(Y�na͟��ߘ��w6M�;䰐*"(���z�w��2�O������dJ���>�Ee�[�/G����TJ�fc.�cۼq��v���lm��癏1��(OIX�4g���)�p�I���[���jUM�s*��S+�LԋQ�*E����+qm.�����	���@8�/m��I�s�!4�cȨ�X��2���,��ಲ?@�&�T��i�2/r��uWW�z3j�6nܡ�d�x�a�RF�w��v�V�F�Iֈ|>=}hpP-�K�]�� :�-)�5��He!YOD���>�?�J�$�O�b��wuvcԨQr�Z�f����Ґ
��I���d�ʋ���Bb�XM�`U��N��q��{z�9|	i,�s)8�m�d��Ȧ�ذ�O��V%���T}������^w���,]AA,(6� ��P{�h4&&�4K��]�"����{W�^��f����s��7��vw�y���s�9f��g3"��a������;��:�/�|��úq�V{,T�b�<��mC�@F$ek~@�߬�C�>��>����!�۾�ɕ�{���q=*|�$�/{?�ȲY��[t���OP}��`*Tx�u���;7��bdB��5U}L�˗?�a�����ҵe[ɔYfL�e*�G@1Q�8]�ƣ
Y�j��Q��S�$���i�+\��L����ڱ��
cN�߰#�A.�
Ի�H�"���!��ţ��5>� �&E�XB��&��k��NO��jm�:1tO��]b�]r3=��ym��*J��P-��r��P�Ԁ��ł\p�<;ud�HD�.!�ve��q~�7�D�XXyc���S	59œ���,�H�@zH�x<���V	s�W�Ԧ�K����N���k�Ѝ��+�w&cU1��>#����B�F*�^L�x0&Q�f,���6�h��^V�\Jo��c��uyU�����l������.�h���/��e�R7����bm�l�rRʎ�uT�&y���<�:���8h�s�&'��'�6�o��$�*���<D�0�S��B��,BR��L��%꺐�$����Q�"�x��,���E>�@Ie�Q��,�iC�H�J	?R�(Zk��X6.�%{�r�v	��v�n�=��X� �E����FC�!�	���!m���uS!�-�U^T8r��9l�4�k�O��;"7UX���j�!�1X*��aϣf�r2�$$���A���^�yuj�\6Mv���H��T&�c5�T�ON�8��f�i���jW<.^w�L�2�RP���BFW�3+k�FY���ߘ�6� ��LY�^�;�#�4bC�4"�!�g��^[/�!���n�0�E�2|S��!����"�r)�>D��-��9�g���`���̋ѰY�(����6{X͒0e�h%��ϰ�G2$9��\��c�Ah^�TV4#�UŘҲ�il��^B3_����eZ�	>����~�E{�8!�hC� ��*�k]����'����A�S��Ì �beM&����MC,�?=bH X����AS���~�xӠ��XI$��	�)�!���Ԭ �e���C��s5���;���K��f�Q�MpHT�6�񭭰66����N�&���<�>;"�1�>ʃ�hZ2��Y�d�-)G�G�90�`y���$�"��I�Ԃu�dJf�.�K�x�TF���3f:zYJ�J��1<�x@�ܯ�� 1ث�5~z��j����Q��/��zAF�9�
� �'6ech�P-Gw.?a�1sb)H����,�O?U ���~���0��-�1e�xɤf�	�!��B}�p@.#��ASF��ݙ1deJ���ߓ�,>�IwhSZA����C8`��ᔰ�����g��Q��J�@���2Q�6n��s@�wU�5HǇ��|���=Hp���1��3c��IJ�FX�R*{3��y�vw!�T����������r�B<��Mh�f5��*	�D��"'�ס#�;vv���ǿ{UU�r��Ġ�Q'���"բy�r�ĨrQP�F�:ƌ{�ՏV��v�r���N�%a��M&4����
^6����Cik�AO8����$��(&#8p�}��2/�n��W=T��E�|E%E�0a8��/�_v=�������f6��3��1x�k`�gDU��YR�3"aPd����M�şn�G�W��[G*�:wb��'iSc8��;TRA0�rmyx�H�9�\lz�)��r�$#�<l���>���)�����5"����b\c����>���n04؅��*�F�V�PGW��#�:7�ә1y��.�8��C�b�*Ğ"q�یP�0���<�������Qc%dR2�t1�}��K<%��V�s��ڈC��OҪ��2�"�jkC�����KM6"�]^��}�a�&�6n���2P��	@~�1y���=)|���hji� ���aw�Ac���K�lh6��l��͛%>� N�q:�^��l"	R)@lGeU%?t��&À[b��]���ve��_�m��L�ߜ��{��#A/q�feGl��6Llo�I�~�}��7:N��K��'�8��k���B���3r�rڗ�&nԩ��P�f�<��Asi��Z�^�X���P�p�9X��U�|�	t�a9��9r@JZ�f�m�m�nl��|[�o��&�8����1g�=�͆Ny�j+kaI�q��h��K�!��/{|)|���İx����:KKi�G��Y��寽�aC��'�tdD�����s�:�P�r�q��7^#+��	5����8VyO$�E��c����z�b<�l���*%��r�YX��s��v�찉A>��1~T��N�X�����i��3����G;C�(N;n>>��l��)HƮ��3�����b��WB8>��'��3:r+��2zV��.?h�~�O��'�����$ޞ9��9M���Ј2|9<��p�֑�Wη?�n^|�&�S�~��/7��GGG�N���g�yU���1YۊV�J_����XR���W��+�e5a������'�H���y���r���\���֌���q�5�ۉ�O���|�����Z_���@��U���e����x�8Ʊ�Ïq��}P,h�O7^��]���^��c�=�d��
��~Xo��l|��h�l���NL�6͜����vlݎ�XwWE������p�Q���G���L�7��$`Ӗ�Y{ϖ�������,}a[Fk=�ȏ��/���!��bRK{����[w 0c��du����&�}�#��5�b�n��Ͽ�&�2[<@;��q��C�es���Xf/��lHo��pS�Тz�m���bNg�(�s���ՋR��R##�ʏ��@u`��.�j��Ֆ�8��{�}���_}�!�=v.���UIܟ�V�X���x�"�rP�\��|V�����ys�*��{&�7	���m7\��m�%,��A��1���#F��Ecs+"y��O�֨�Ǟ^��9m5��k�T|�z80k���Q �nI.ȫ���rwj�@wR�=�̋8aޡ���S�m�.R=�HV�b� �������P��6-l����8�ȹ(
"�Ѽ�Ke��m���h�|%ܨlh���ޏJ�G�05/@�В�0��y��q�����f>���H��L)1����Ns^Hūő�7��O��'�_����9�s���HL�!;7!!爪�lچ��}������wf�i]G/,�oq�{a��/�,���(����v�%��jq���W��}:Hhs���	,y
��wul�C����'c�8���3��,�����C�ى�vQ�����>���7��U�����lP�,!��$!��'�TтG�zN"�jAc̷y�1-_��'����;���c���],!ZF�!sJ������ ȬQ��x�pcM}3�|������ǳ,����Q�6����ڶ1��;0w�ݍ�`L�x{��iy�^9,�_}��Z�����9��Ͽ�&����T_�x����us�ǋ^�FqY$�;�}
~�R�]s̏�%JȆ���G�)�<�z'�
��%�1ƃ|�cϾ�,9ΒX��x�_p����o$l����VLm���	�Hȥپm��/>��k���W�!���;�fgRV|��je��g��G�Zg�x�≣Ȅ���U��~RN�ۧ��&����1I����C��G>A���1�����,��nY��WU-�B�
e\k��ʺ|*����n�lz��CQ�gC�VT�:�Ef��(Xc�Ӫ�!�Gbc'v�w>�Qs���?`��Zͨ����t}��Va�>�ucw��g�Uo���_��tAmm�c��9�yC$~�$�Ǫ���O΁1�QT�AOi���so��N9VA_��!&��v;�DJq�P"�>�jZG����B��d����z���۸���i�je�WA�d@gY�۟֊S�C�Cc&�ԗ���	x�����Y�m����WTˊ9JV~��A�c1d1mY5�P�ǎ���
���E2S�R&����0�F�t�mry��e�]2��9�V,#�%O.Ņ瞩y�A>;;{$D�"g��Z9��+o���%�6�.��c�C���z��;���S0it3:�yZ�[�d''!��K"���_ߤ�L��I���	�]}�oɓ���Eb��12�k�%��Aj�����*$��U�Ң�	�ʺ6�p�q���֎�ȉs�8��!�<���Í7���"�����l��U~�۫>F@��x��d�\BNm�����O�S���$�MFB�ATV7`�x��^~Y<S� k�w9�u(�a]�$�{m%.�x����8p%1<c�A�1�|�}��^��9Pę����uj�^�y眉��.nm�Wsͣ����#MjV�N�N�ř5t�
�ߴU.���5:tg��`sK�5�k��"Ƈ��%�.iw�E�k��1�>�����Mk--m���<P����_���5r�
�1�,bJ#�R���_��A�ԣ��J�;�����˂�XF��Rrc����9�nD����fb$-�v�(��*|O�����7b395qX�~(�!U=τ�,Y*��|mGN��`��)��e�x�JCĚc��(��hv}�(<��+�Ѐ�g�<�k~٬�%d�Z�F<g}cy���+W+��mer	,yz9��w�:�H$�S���ୂ�v��q��v�����:�5��q�\A�ry��B/��~+���[��!s�z�5xVz�~�
^��Ѓx�3L�6-���Y�H�����x���+9/0���Ug���<z*���Ǟ¾��JAqԒ�ڒJ��?�r��Y�d��0:��J��T���8~�rm4б�id�0���BU�B�|��>��nS�	�w^%���ʺn�nl�ۣ=k7n����PU�UxC}���M�gq�^~-��>���~/�g>��Kե����g:�dc��l֡��׬Q�vo�R!QZ˄cړ4�lN��᭬�s�_�r�]K�F��D�a����V����U�[NGB	I(����?���%�m^�Д��p��-�C�C��C��X*$s�Lf��?*�H���n�k��%��&$���2�IKX<�� .��n�KX��nBT�T�I��!�K6m�'K�V���)�v@
�L��T׌����.~:�'!����a��"Q��e������^��>\/W�k��ЉW=��*e0�y�k��h�U�ni�"p��r�x��P,[.h�#>���	�̂N2T�w�1ݠ7(蘾9T�֎�z���W��v�W���g�(O�jH@>���+e6��E�̠�nIY��}
O���N�K�\�Iy@�v�B&m�*�&d c�(c�bś��$���#S�rJ�*4��K4ٰ��nI�_�'߭V�ʹ�7@V��!�Y�
�D�y��]l*�G�W��㥕(�3�̚�!�s{*�ϔ�y}�ɧt=8��$w\�S�Vk~Z�U��Aɬ�8��#F��+�Uk�i6tm5EO��;��[�~�a2�V���)㕐V�[j����P��j/����cE,!���߯� �FP�ɦS�*y!k�1�����ez��ΠQ���B(uSvti;>]2��>."kWx;�CeY��6������1d�HƖ���Y�^3�b��;���K"����ێ	��SH�\�K�&���g������X}�c@��t���Nɒj���.O͖�OC�Vl��q�(2]Yg=9�5��l��S�r>�U���rA,.��5��3Z��A�����fu�\�����0��P4�����|Jag�0���[�������W���%̈姺���f�Jm'�e,�08M�.�M,�Ϛ�0�0S���t
���}��EU�3�����9d��Y�`[�hJ�g�
)�2�5��'�?�P�
�*���2m!�FPPg�S����3��IKyU�=���U�B)���L�gƙ����y�͟�0�#𤕷)����:XL�����Ī/����0a^�Dj�\� �*��f%�!͝\&�C�����*������y����&�1n3���Az�I�Kj6�Y��ʕ'�+e�x�~9��͔�(.�l�6����|y�J�Đ8�8ɩ�/Y�"��L�NPn�N1��W�� rE�����\�
�J8�WA�2s��cS� U�ƛ%-#�1������	U����c[��Ŭ_�r���OU����dp8Z�_d)�ڛK�8!�Dkw$I<���d�r8~�bΗ���A�,[|����l�)��-�[H	G&'U��1nY�����,�F�/���烇�݉rQv�*A���~eR�^ЍQ�^���`L����T;Iw�>&��ǐI�i������iɶ���ԝȔ�K3��r ����Z���P�-�M��0����kPi�S�JTD.��l�J�bza��AAK�T�L%Mnq���鄱�e�F�Ɯ���{UR.�R�B	��]�I�K�6��ј���u���Ք+��A:�+Ck���)���˾>��dg��SP3C�uo�c� +���i��B�HIgt�z�sF�?q���.�B�ͮ���8v5r]��؛Li��%����Cl#<�����b~&D��,��P�� ?K>�\��0�g(���R$8����eA��xH���.	����io�F���މ�>!�q
J4�;pP�tH���S��۷BC3�Q�J�2�Y�U��x����
Gb��M�sQ�PMm� 㙵�g.�D0�tV�u����N��:�,~$F6AM&y�@O�! d�*d����`?�n�.O��Cci�Ҷ����cբ�N�Wb�|8*�٤Rp�|�Ms��rV��Z�`l�3Zd��H(�¾vC�p�J���C�0�d�t��#�A�1�DB�t¡UUנ`('��BY��l<�@c��_�(F��޾ACie/]�PU(�%�m�`蓊����A��x�V�,N�n�ءc�N��^]"q�vy	%v KZ<����*d���@�І	-:���Yfn��@W�v=�d�������GU0�G���������%��kO@�l��m������������rEb���ذu��$�{�=7X� �ɰsxL{;�L�{ސq�ڶ�+?�U�Mb�L���Xz��Q���~�	���ߘ�-�_�!Ϸv�:YW9[^�1(��)���M.���>�~�� �~	QA�q������֗��"(e�"j,5228�f������а^���z���ʫAA��(�`*\��9�U�X,��_�F�XL�}_�
��x��TH6���`2rt���#�;w�s��nW�����Z,y�YA����$`��F�	��Tr_{�{p��a�^S$$s#���y]KV��
�~�C��U.t�wJ��M�!�v6��\���p=�� 9<�U*��F��>�}�UX��������K2��e
xj��ڇo�4�LW( �����t�"���-[ᯮG\����^|�T�7+�4�E�wQ�%�b��c�蚕�ӃD2������_}�xT��W��.
�i�s9=��-�s<�Ybj�8&�?�߈/��Yh#�*[g^��6�a���}��ޑ`�����Ӌ��Z<���n\��fV~Β�|��{��{M���{��$��v "���E_��ߴ�K��l�h�?=�Y�6H��#f(��(u�A,���JTK]�^����4Vf���7\)��������ߣ�ާuw���w��y��շ�C���6W;5�48�����S�U�ö�z��(���1�ʵ2���~��r@�ɑ-�t9Z��	G��Wq�P�UUb���Z�Y7-�mw݃��m&�e+����ǣ*�t����ޅ�go�
 )�Ȗ���7��vǧS)�F4_28�����-8y>�4�,�7�򰕻���N�>�폇
�	in�l�k"���s�n�;{?UT��]m����	�p�e��ĳ/��{+ڈ8t&CY���H���]ǎ_։����Ij��!�GT��Y����O���,�j�G���ݲ�s���k4�x���=
T���JV���k�ǿޭ��FU�4�$���PO'�=�4�mk'�m ���w��s�_�揿�Ny����g[�]si�5֊�Y���DH��	*Ā��$��<�Z�a9$�\\�͑ui�q�qs��g߫��d�RE/�� m{L��fN���lԆ�j��`N�����8��Yx���ĺVib���b8r	�5�ȋ�R8�,��v��g��yg���o�����{SdQ�b����v��l\�x�Cqb5r�8����cl�.���k��4q�K�3	�x���\x�n�z&��"��
Jb�;٨��}@�
9Ah r\;�C�8���g����'b+)�b�{G������W7��~�<����Vb�=�(X�����u�IB����V>�O���^���Y&���B&B�|��"w�DzcR�X�iG`:2$kt2~j�D��
#AX���C!5�K�
9e��I;�A;�1��Z��A���OU�N]2�����p�왘�^��l�&���d�Vy�nܼ�J�q��Gu1^&�ٽ��w$���AM]�x�>}��t�c��Xx�IxM�BV3�Ų&�U��)�u����j�����~yNء��fC��*���cO(�9	��r��%k�����Y��`���0q�����n֬#�ݳ�_q)���{௬�2��Ejߊ���z]s�Er��J��ssS�#&�N+�L�(��~��C��H����m�q����p��~4�|5�l���Sε��0������ވ��Z�R]u^�͟���jmpWU�u �*�5�V1.�6C��X���"�2��8�B
�A\�h��������a������a)���AX�hE�;��93y���s8�J�pԡx�ŗ1B�w�vP�T	"8l�:K�X�lk���a�IU5U���є6���Ͽ����Ւc)+�+�����ہ�Sg�����w�!�ƕ��:W��O���x�b�m$�����p�� ����J�2DUe�	��;�=��N8
�=���ե��n����h_�٬e�T���~������[�];q�Y��ѧ�jc��U�	��Hs��*�S��U�x��O�ǰ����s�8o#!��S�
���y\Z$F[]%��;}]�J�S�<��� �Ï׎qm��n��������SY��t��v��7/Ɛ����/��6�\��N~�k�ǉ��<�GŸ�{�)��ޒ8�b�N-�՝}�a��`x�ǨI3�igV��H~�����U���������f�x0�G�{��='��T��2u��x��e����g�QsҰb��y�\�_|]ַR���U��������-g����j����	���BF��������}	�S��aY�����%ԉ�fb��W���/ 2�܃����c��1]x�IX"��S�#��k����W��k��⥷?���O�C-����b���~	����j���'UC��:�$����Po'*}�H��x����Se�����k�؞���`�߯F&E�A1��(���e��vP��_m�Ï�^��E�CVB%7.8�X�׆�|��_�?��_p	j���,��w���}��h=�]}�o�$F�${���8O�3�a�����}��Q�����&�{�E�"�ʢa�nXt�blڶU��� ���e�����h����/��� ��c�����s�T��SO�8�m$
f�1��M��Yb�9a��T��ֻ��q\��&�ׯ���=qL�l� ~ټM�X�0���2tuv`���p���[[+����ܻ�,8V��$��Ib\��A*�D��[�p6oZ���x<5���J:"�ӫc�5r��u�m����8h�>���d�
b��
�ˈ!k+��_����^�두ɁX�u\��D�~��	�|�qX��J���n�@�"VW�&MƂo���Q�~���7O��#��}��ޯ2�vvj_�mN��!���?w���ߡӺٜ��O�0����t���:�����wk�����\|�;�a�����ƻPrP��S>��b�#�p���p�fXI̚9���,.R�QɾZC)��j[�`ѵ��;�DM�O.C���!�}�\y�)rAR8Z~��G��Qr#��L����9�t�{��Ե�%�+?C�����q�
≠�}f썟�3IJ�2y���������_z��F��?���ᖛ�DahA%���CO��3�T�_`��:��m��p����MB�Sи,�]���S�������G���C��J$$�>�سUկQ�a����+@Vt�Sx���q�9'˹n�w�a����kM���b࣡a�\���?�
�x�Œ�_��:q� ���$M?p�}����	2����>�C5m�?�����9�gk����%Oaٓ",�+�����\-���*z�̞�d2��ѣp���2�aFA�T.�wV}�L<��)�'��O8�o��)������BA�QT����N[�}W�M*��e��^�?��v����a]���رc���W%ٶt��o���/Ma�0V��MbuXf�{�I�"QL"#0�e�d\y�M��Pd�S��h
7�v�z�.U�s�d|��/rH}�q?e<�zz�¹q�S��]G��4J�%ӭ���+�b�~�h�K����"�a����\:"q�Ă�j,��H��kl*�L��޾<��k�o���6ԣH��v��d�B�DW�GrX���b �H����W�>�2�>�LjvaP�bD��.����o�n�\�^X
k��|��M~�`�oJh6�9�^}�'bp썲��D�iFC�J�z
��F�������\OVp���6��W�l�^���Xe���.L��'y��դ��[?��OH��S�5�2$rhG����`�>S�dT�6���V�d}rQ]:���۟����&(���1��Paշ_��3`I%����%ŵ ��xF�"w]=�r��	��!.BЌ�$�Ï7�P�0A����0�<����,�;�IU70���xb��+�=R��Y1�}�9<���q�\��)����T���{�H���|��M0{M�\T�aCY_��x���p���ᦼ�v�R����8Z�Nk�r/ɥ-)XȨ�7�P������󶛕�'��i^�D��0��wⵣ^����@US��xo��������{7c
LጠR����8b������v&k���[��^J�H��Q�X�A���?���>Y�~i[R��&9��x�]�!�I�MYT[c�)�+�E��>�g�q�+?::�T�BCU��4�E	a%��	�O�iO˿v�iS)y��p���^��� �4L���o���q�Z{�h:g�N��{L,�-`Q��^~E3�W�㲐2��U��̴j)REk�e�f�I��l7-;�(B�2p�e+yh��n/�� /�BV ��8�[�RX�n�6�V%��%x��!��Z��kל�H-ٱA��`OI~��rhr(k4�0.Vr�Py�g��
�K�,�q�-��oٲY:��Y�\(�Z��:�&����]K�I=(��;A���ς�\��F��lh��ZsHm��dY�cܘ1����͘@ki�pK��+�~/��,V��������VSmVUv�ɥwhY�#�h�K�U��Sو��z6_��_�cϝ�#��O?b��:�Bq{�f�Q,+�5imn��U����]��(��O�X�$޴ifN��9 �S9E˄*+|2���;�d��Q��ۛ�{�2�)1�Nٟ\"���r+	L�U�Ex��g5��Dfn6�1�ϒx__�1�!��Nb��A�/7���p��5����Y�8,v
�qP�e�<B��#Nq֢!��RmB�PJ����5���͋j�	ڢ6����$����j�����V�*n��%�8M_��6r���/��ʝW>���S+�^A!��0��j
�0d+�Gz�eC*�딄�.h�+���x9tӤ3H�Ysbph�hN���
j��%�|(�����8�o*��S&�)~f�3�����|^m���f�6l���ѹ칛X��֫�����Il�ڴl�jl�x��OPFcօ�Ⲹ�H\	�y���5鐏\h%�M�竀�iEMm"��,��\A���FQ7��)R�%�jj�Q���������gsV��^��������CSLdҪj�[>�W���<VA�E��lha+�EB��Mr�,�$����&#2I�t�BM�'Ȗ�%�$����4�Y$�3�(76i7��L�\��Į$�-i�N����U����@K��-�|�ֻ]^l��&F�E�۽]�E%��$�n����tj�G�%Wݍ�x(�͞�D����EM����9A"��Ea�)"�rL�Q���Z��d�?�YАx��(�d�$�C��Ї)�Z��b��_�i�L��Y�
<o�	H��UgS4
�P#Ȥ�fQ�Z
���A����f%�a�z��v��n�P�r΋�˥t��ZJ��G����0Jb U�ۤQ::?��	U?b�r?��cBª��J����Ⱥ?
�q�9�yLHx�t4N9� ��Z���,� �#3�#���j��4j�����g�1(�˻�!A�1H�;2���$�i��UR$&qy��s`����"����Il��V��m�����ٍ�l2�T�=���a3��پ�C�8�xt@�/�h8?�is��p,�c��,���A}V����-hj-W��r8�S̮��yy��@��y\���E2_RY��  �*p��{w�28c3mn���u{�k$�mi�F!�F�p��E��l.Bmu����5cE�Ţ�m45��O6��ʄl�pL���`0l��tt�O�5j9���r,r9���
5�U��ģnGY�Wj��7�D�LD3�L���֠@�=���-��@@y�dVy(LrX�J�B�p�p�#���C�P.���d�����&b�w���g���y�ʴ4�iHH�]�q��Jf�nBDb撬?˽���y�W�`���1����'���n�hP0g�C˙��KT<��ǡ;����݋�����UĄ�v�^�;ת�Yƅ�z��9�WL�m<v�f� 7͞cg/D&�W�ľ��?,{���#��ǏE��s�d�8���8R�5r�95�ѕr����&�!ә+K�C#;�}�g��B�BRp���
�F����1Y�ֶ6tF��l�%���QQ�*H�k���B^)�oP���}���O~|_P;4����y�~�m0���is{!���	���@7B#��l�2���Ѹ��7�p���r�ܪm�&/�T��;p�⿢k�1���a�	zsR$KB��'���O���w
:�j7�N��MMu�y�Ƌ�}�}"�RV97��L�{1�1m�IY1Ғn��-ο��g�R�c�g�������I8UK�2u/��C�ry� ��&��ȖXv��Ήѭ�r�b���(�E� ��%��bb��|���R1��_�7m����G��Y�≗^E}�B�r����;���R��f��^�]��iQv!���9uw��f5|��Z��	t�xR¤�>P��	9�#�Ngr���+o�%_? };��ϔi�a[A�Kl[%�Z���>���r��0)��l����9�����9��ߐ�͂85[\d��c��m���87k��h��U��$�q��#��bnft��Ѽ�&(�)��9s�l���i���]�dҤt(�����}8����������xd��5�4<b z���Ő�ޅa���9�L'3����Y�0:+-�HHV��<$:�����J9	,*�d�s�q׃�k[~��6�]<�d��1�����_d�oO�/PS�šǷ�m�6{�l����:Q��l�,���OJ~?�I��;�l ���aT57cd$���Ξ~��e�"NȒ$�V�X�8�X4����Dǒga�����"���O}��ׯ��w܊=�,���#9e�j	�‽�	j��,��Ϊw�o���b�׮ߢ���_���s����E@��+���|"<�g����Nyw��	8\^E:D��CC>T�Au�\�e1�v���l�<���ߜ�$���ǆIYs���y1�^-����c�i�л}+n��R\w�-�����=���1���$4jP�^��5��"g�Fө����%�?�p�w����SO����>��fSq�:�`L?A?���oK��r��q i�~�ˁMk_{A ���~/�Fk����e�v�3u�r��d�>�Ȳ�l�.Rf^�:��unCP⫷��5��N��Y�D[�z�;���ƙ��Eb�M��K8��̩s�Ձ5"rA�].�Ȓ�K`��Ͼ�lS#��8��#���b(�FC�s9BuC�L5bY_@mc�"
���K�	�X><����ǟIL�R���f���V���C$Kʓ�QB���x[�0��~,:�$��]��:NL��K���_�`��h�}E ,y��{����s�<��y6lآa3�{O���P���}��zl�F'94Jh����ct]=�A��W'n��
|%{�5nՊARdh�H�Ë�X��V��l%��d������#+��K/�7?��j6'Ux��U{����[��}.�,�6*\%���K���E�c���pΉGb��y�\6EU������g��ܬ��!_�XmP�I(��?b̨*��j�&��u��?�\U��45w*{Z��B,��S�-G�}���
�i;�z.9o!:;1k�I�g�)ؼu���
����&�:�����m�N6L�Ǝ*�n���˸���e�޶	�z��bIDcQ��9��e�9�c|��jt���akI{���;q�������7]q֬�Y1�	�#*��"��⾇�E��ފj��/���[n��P������_�S�t:A��HR5��6��~�;���ꐓtś�*7��э��u�_�r�Zd�|�^E#!8�����Ix�<�MK�v�[iq�w�� �}]]8�ع�7W;��T��\36Z��Ѐ���a��-:��>f4,�m�|-�q��GP����^BN��І�}���s�x�jlc��֠��Q�t���(]d�:5R�?�\[��'���0�E6t;�%'����GNb*��k��I���;�	�K�PĮ=f���>����;�nı�A1l�z	kH.렄=�;{���o!X[�q���0�"�����QMC}M5��!9d�nFJb�@�W;-0؊�F<K�291Wu��S�KϽ�"�8d6�	i<f4��F�Pps�ކ_~W�S�ðrЮ�!5	**��U��FW�f�5�	�|ℳ�Ň�P�Ђe�Wb ��u�k�2��N�
<~G`��Y�P%�jg�.�=XT��1��~�\Y�܀��P	zb��Xp�1��EP���d&���%���tK�� ��B��v0��IP������ ~���pb�=u�J����$-XS�WV~�ۻU���b$Cbr�(�����3D����Mn��IR�z�x�ض�?�W�Z�ږQ:���=��T��y�)\tکH�"�\��M��#��0�m,uu�����a㛜s�\����S��?���:1\�+���5�A1���?��K��ޫ-����n�0'\���׫רO09�61�.g�r�i8Kb$��r�_������������^խ�͕竞Lvd@	��¤��K�z���{�a�&w�՝�C����Ko��Mn�gNAZ�K<"��n� ��)9�x���.!�����V.SVO{���?㶛o���?�R%�Й��"�����uH<�G�����q�z�#z8��V,��Ϩ�o�hu���Mò�Z�.�U�c�9'�c�Z$��p�%�Lđ����ʫ+7�}p�Z2�&� �Ay��0�h"�U�����n5q��$f�����2�U�R<�9���\ޅ���1�x��٬3.o)��f��6��?��}TVU�AJ��ąt�r�W}�3���rlټ�7�u�0="P>P���}���JV%na�:�i�%s�N��k|�r`�G��#/^��~�-���}�+�wHJ�g&�lrQ]��jҾ���}W]r>��L�s
c&5��~���-�d�ysQ��<�U�C�R���<�'M��>�
_�V����d��FP�W�>v�-kc�ꖈas���U�ќ�r������P%H�B���J��c :�iN�&*K�/��c��t��|���`�8`�&$<��ų����n_@{x��T�#\��{�p�<g���Y�� �g��Z��t	�����z��*�RńnFP_ڞ�#����e/S�'��
�qHB�\�%�?�� C��I����|�Mbت���0���r�ƣ�lGH¿8��ZF��ǟ@g��'��ԉ1`����|/r	��e�nډ�/>n�K��,^��=;�"Xz�8��4�g�}dx��w��T��ko���/��&kVɣzz�в�t\�hj��1����5Y[�p�߮9�b��}8̱��^0�0�������`�G�ޢ��	�X����iLU���hv�o�c܅���cg
��V��k��G�+�b�l&�ڰ��㺭���r��Q����+&.wMr��/�y��s�컷<�l'���¿����Rzx��T�1n��!�u��>C���f�~Ӄ2>&7���*AlaeDe68d��������{�����W��;�tTxk��2b�����q1Ӊ���Y�&j?�wK%5Y�*C<��m�y�͌�U]�pP��P����Y��KZ���9�Q�4��
x�)�2�E��Z�/K-0�O���cO���7�i�$�H�iծ%�t0��wؘ����x��ux��K�Z�DBQ9G�^߯k�7ƿ3,E���e�\n~��{�
B[�d����T�ۢ���%5G��OO�X�!�NA��f͵�����ie���;c-�ڑ���r�|��f5,&�� {��R��Jy���1ޅS�4�9Y����:��R��f�!IG�g��0��>���b�(�8�A���Gxm�{�$9&�m �H�Y,�e]c#���N0ł�mw�[K��CIb���Tr]�X	OT��<�X2�CI�J����ڊ�/6Ά��^�+��rT��r��9˜�x��/Q����Ǟ}Vs�^q^d�S�@���Y�Ш�S*���f�8f+���ù_��e��R��f1��ʰ�h�~�f|��:]d^LjJ|���e�њ�d�����a�:���J��,�c�2�V
4�D�ףlW�X�W0���L�qd�����H��]�V�����1���u�.DM`l:g`4k�3Ğ������`:�:�YݕA$�:M�w���h�r%�)=D6trd�9�.o�2���H|>�toJ�G~�GC����P<�,a������(�I�#=k�|��e�����px�G"!��kw���N���P+~�8�KWTNƳ,AӀ)��2VY��X4��v�w��ƛة�F$�(B.[PV/�KkM,^#��GR�JsXɐT�~�X\6���D�3�5ȕ��)/��;�숁"��u�J�}(���;��T���F�'��4�_4�R�W3f����:=��O�|�˚Smv��k�r��њ�[���*��QxJS�H�P4�J�.Ƈ0�dH��3Y�TV"j�J�����!�˞p:7��Em`�}3�-�Y95��x��p���la�?�%���4����`U���Ǝ�;��@Em�Q�ZdM�sQ2�v���:���UQՠS��)򑦀{�q��)q�9�o��t�$��Y�@�ДL��y�w��v�$�x�"*�R�mЃ�|%�#�P��4�U���`_�c�,���Ӟ�)Je~s�8ƤV<%�2d-���Khb��Ԭ�i26L�YaLy��GЅ��ס�#V���Sq �FRY�d��$�f2)Ë��g!5�III�1�Za��cX�Ƅ�Cg�%K�Rg._�2�g��t�5=w:�P� mR��������Z�|����k��hz

z`�2�ڽ�?a2�ʇ��+�{�,�RKE�7��u+�U����
�>�rr��qx�lp�h|ϰ��'���D�f��*ɩ�G��,cb�0�W(�3)����'g34R�]�o�I�u'���5s$�\�ϋ��9EM��3[�=/��A�h�qk�h��u����>�fEwyU�3�~�|�LZ"7�0��l���#{���2O��\�𛌰DɕL�+��V<��/bX��$�v5P���<hf8S�I�|9��~6g��e�]��,�u�����2�`_�[(�YȪν��d;�V�ؚ�:}~6/�W,��T���#���w�������2ИP�F~	a��H�\�K�:5�Ŏ>#�f*���f���34�'���ţ����aq�/��Џ�MQJ*�E�_V�����t(
�������C��n~���C�?.�<�9�iUU�24��T��(?�d����Q�6)'o���CCz�8���"$J��ԩ������L����S�<�?�J�����I�#{R_�,�۬���r"W��|@RB��?����_���׵���Waxp���e��`�2��I�bW�46h�E��q�&�< ���E+��d�%[3�oe/�~��@mu���42��ؖN�F��Z��L@���(��l�b�@Jb�l2��Lս-�;�dݚ��m�k�L�dT�k���T��l8���	�I�k8B�u�Ms_N���n���$��e�ض&��"e�i4�6%q<,���re�g)���3���@7v?}����Q�쭐���=jb�<���Ԑ�{�V�4���XDּIU��N��r>�6���DG����yN��HB�P���'�{��#!��Ў!9>�هym��++=���Ѱ:���tB<� 48�G���}�ǥN*/�q�7�%�ce?Řq�c�Q'<�FF�%W#��X�v�%���e��8��p��>]{����Le;p��.����C�P�d�AU�?Y~ҽE�C8bΡj9���'�����_)���sr�y�Ԙ���h-������gy��ӎ��~9)�#�Y���\ AR���>C���Y!Ƙ�Z��{.*�^�䔒��00��˯�!P-���U(ܔFpl669�q�� C2�S9@(�DB�}JMp%ۂW-fCq�?���1q*:N! �ن-;���'�����P9��T<��brDu;��G���"=�Z2��s/�*�J��#��[DQ��c�m�I'�֦�FBhijB����;�=���BK�d��f
9
*�T����W^���h|uu���7H��Y�~�-\>�z��ߔ�;3���p��)F�F�>��e�h$�������g�dJJ[X4�+�uqk%�_���������b�Y-�g�W��|�n�٬Ȋ]��|&1���A���j�UI?�1��Yd����;%�i u�xw�ю_����\q�"�-y������r��x/<��u�=p���*�~�3������Ϝ�y�/B44 ����;��P�{o����3^z�U�ׄ��~T�u
r~8��n�A��s��o��/kY���ߍ�n�UB�DÂ"HYX�{�(�J��ʇ��;Jb�8B`�Vң{��;Z�,��=We��#{F,��h����|���xވ���&�f���_v)R��R��PW�Ñnܨ|��Fe%�{mZQ��p�dpx���pႳB	�kK�ٜA}K5F�47����t1��M��&�K1�Ħ�ӎ?F�$3�x�D0uB�,�&�5�`��yX��U������+����I��S��^SǢ6HZ7�zŢ~/{��|N�u�|<�ߗP3j�[�s,�0�1�����<�tT9$S�A9T	�:e��y����>�!$���l��e�e�F��� !D�3"Ʊ��VTA����w�����O= �3C���a�ƩwB9N��Ʉ�xעx����>
���RK�%s9���Ur\�yTW8q�I�h�)������0�٨��_s���K��e�Ci��ݠ����[���?\����ڽ+V;�rV�aLӦ��o��/Ph]*g	��(t�,1z��:�`"g&��S#�<b:&p�y���ҾR�L��0<v򯜀�P���!�(1}N�#'��������=}�:]��D��TLP�	q�,<K{B"�l� Ҙ �w�� n��b\w�mh3�pe�/���`����F�غN��M�]PRPG��|7,�7��.1B^=��EF�6��N�u�_�1��Ⱦ_�ܤ�LO1�����q���D}c�"D�Е�$�
xp�e��?����u^:���a�)�����6q��~l��L~�Zq8�-�iq�Ew*[H,N��{�4�E�kh$��j�>�ZO�Ňe���V�{�Q�w�4��U��եsԕ�%��a�K��0 ���l����	!�E�/�#��b�t]��.��)�:{q���.���*)��q�����NKR�-d��CO���$ھ�Yy�Ҳ�'̙��?r�{R4�5iv�u�D�a��i��U_���;����<B�Ɔ0��g�?;JF9وQr�bho��6��GM��^r6�Y��[����:umc!\~ѹj�yZ�M��ݲ
öz����O��g���ӝ�L^�e4���.<��[Pc%���V�X$Tb"�c�f��>1�u%���sX+6�Z���A̙��j|���D��Q׶^	�B�o�RE�b<��Ǌ�N;�~�14����RN8�7�8|ξ�?n�}�v�v�����c�D��s��v"%h�3O²o`$S�l��hE¢#7�漳��P;��PV����O  �/IDAT/r��M�{M��)��k﯂�ת��S�f#8��C�{��+�
dcv�ݽʤVm5��@�h�ix���PY׊X� �%A��łE(5$�����z�C�+^���R]�ƻ|�-]��]:�ː49<�K.�s�G*�ƴ���{T����q��Q��H�1y��j�1��.w�+�=�P��p�B���S	��}4��v��k�h���嗞��j����k.��w�.WSR����vG͞���*��[9a:�~g�|�1�io���=�hU¢�\{��x���»�̳9�\��S�d�'ae�O�˗���u�0y�D̙�?F�	2�c��ǝ� ��"@NB�
97\z�怪���Kν�׬`@��J\r�4k,��B��}6m܄�^{��'L�5W.BSkZ��W]~	�|~9<��ӋE����"�Rb�8�`����|�O��m-c0g�~b�"��ǉ�~v�@�ZU��'�#^s���$^���m"�{���t�NN��;_}!�{whG�9g��寽ב@8���_!�7E�|�J~��6���!�P���j�I�x��y��=�)��7��	�N<�h���pWx�5�-�N/z2e���L��3�F���O?��S���ާ�H��8��eႳ�+E�k�	ܻ���Շr�hΜY8��c��(Q̱��3/���}�ũX�{6�l\���Sf�[�r'~Y���Q_�o��9Ys�7�h�\��2W1�żش���Y3�3�ؽ�Q'^�j��6�e%��Kl}չ��F"ƥ.��xOָ� 8L&�� ������e���_~�V6����.F<$є�駟���|A�	q�TG쿇@�0E� B+N>�r8e=��9�����2�sJu�Q��9��3ڕ�K_a�a�Q�M�v7ብ/��k�&�) v퍓�!�>�(얛n�mw���ZED���|����p�R�p��g���Z�������8\r�q`1������l�ju��I�'Y��c�;ब����^vf�.K;�"�E@łQѨ�Kl�%EM�Xb��޻��R�)u�e{ߝ��>��s����1/�3��/��{��|1�=�TTF4�y�&�������bkO�.�q�<,�j�:��5���'+X�����J�\TWU�Txw� ���[q�i'a�F�e�����B�g
�|�C��dX>a2f�|6��y�aڰ}9>_�3fN���=K��{�w�C�!��?�r�=;�5T�a��T�" �e��Ւ=�W��O�S�i�|�Y\���X�����مj0g֩���aV�(�)��O=�Pȅ��r�?��s|�����a�|��[��������E�_�8���L�ʵu�*1Ǚ�OEJ�_<w��7��o����tk��+�J�8S���z�٧�{AEM��p#%"�mL���o�ޏ��4Ur\^4u���o�}��	;wl���������(��x�ko�M[6+����[�/V���0[�P
���~�x�%��������=���Gq�)I�<�eRr�-������*�4�̊�qa{s'^|c��d!ƍ�����^���}��"I���G���Pm�Rѳ:�r�%߹���J�-i��+ƏESW�x`�V��^��(�u�J6����j-B�˅���p��WC�)�:Z1���x䩧�K���[���P�KgW^�7��k��UM�[^�]��x����PUU��;�B��II_��k/9�����]���uH��H��W�-�]��\���X���{$F�P9I��&����	��	s����3vIǺ��@��רj|Q"�I�X���l�Vȳ\(,.F�^V��^x�ކ���Mšr�n�/��q�jz��@^qwM�t��z�U ��B������Uzf�9w�Sb�^łSf�����6�~�Z5M�b]�(Gʿ;0B���G��zI�5�f���b` �<�n�寚�VVVHZG$�5I�K1p1����:�qH����!����;��#��C�>(9ߑu���m,p���w�W0,�K"V��\?�/V��SR�$\��bN�u>\�vx�ּ阶��5#q��+P3�AT0U�aܤ	���;�����-b��PZ4�}��eǴ��X-�5�;npY����rF徾�ҋ���a_�iސ�H/fU!�!|��L��j�0���]H<�ۚV&oΕtIx��ˁ.��;�A���[bl������~u�\(��n+:%,�k������Hj��f�G>뛯�/Ѩ-H�X�8s3�吒_����:�������7�t�K~��8}�	ri��{�=��/�zM!j��3W���w_���`U�v�S�
l��e�B�1<�m��<G��7����T����;;*9��n6���&$m�@��v,Ռpw��\�D��硂:,L��_��tF��Ƭ�h])N�*��!L��V���مڱ���ډ��g��>�d�'E]4:C'()���zV�\�����5%H�gC��@����=*����*�O_w�Dz��.�1�i��AY�d&�;x��zesc4��I?#Z��|�tRĠ֥�_�A���4�����?|�">ڪ/�MD%)����8��j4(ˠ�
t9�;r�7'iߒO?C ��Wf3�ۉdފ��4�}����۶n2`Ţ�>����];�0v�8�r���Vt)n'+g8!�c�V�<�Һ~YN�{"�Ig����<Vʾ�$j	(��6�;��[w�cLM}}�ک(�Pf얱V��X��ёx��+h�| ��8�z���{������F��Ko'ےD<�T��ޭE�|�LZ;�n(�-�V�<cKk�$<v��7�$E���|���L���M�+�}�o�q�=�6�����結�9��m�-[�qܡӱ}���n��U��(Ȣgdɰ��v	ه�Y��S|'Ki���xUD��{��nm�ڵ��*�+�l�!��R)��M -[On�髳�G��@8$��x� \��x�;,_��2�������{�y{d3�r�]rpb�uP�u=Jx��uz�ً-$8/��*^�j�����Oqp��W-�d�L�֊��)'����G�5k7��I�u1�ɔ����v�<�Y�݁*Zh������E��
	��zXK�Y[Ѯ�����pVD賻�ˠ�݇F}eAəaF�َ�gt��-�Je���{w��Y��Ԋ�&��\�!�ȋgu�j�<B�w�V0��_H<�+��)B�,"��]��μ�VտѨip�pDҰ���)A@ ��;�wb��)zV"�h	�gר��K>�d���s�9���S4ZaD�*#�<����5�E��w!+gBְ����]�k�=%*2ǎ;@�#��#
�93�ZP�<{䡠@6=/S��r��>�%�����~ZēCJ@�P�v���As�3��$+�[��aZ�����$�M�E�K���	1b���zVG�X͔����C��A���s�O�h'��eɤU���0�ɽS�/��ģ���Ds���,��Lgn�[~����SĶ����bP,���K����JA,����R^(���K�����^�)��7s�ɞ�q5���<H���u�K)����K; y	��e>�rry�-�r�57,A<�SB��;���\�R}X6�'����\�I.��=9)x�k�@Q�)g@<���E��J�9���A��`D�!-��W�%�L8�S���%���6��|���6��M�/I���S[V��T��$~�R�,�P��*s������1c��/m�!����q����95;�ۣ�e��<\<0��'�%h��	޾X֔HcQ�]�*	��������۪�ƴ
%��C�#^�G}er�I�4���H��o_"�t�bŵ��NVA,���1dz�0���X�q����!*���������HT?��j�p��VY_�і��_B�r�H�e2j�fU%� =vV��,����)n�`yĹ<u|�|j+�;R���e�^�l*��	V��9�)g�_�,)k;1i���x�I�B��3^E����#N��%����$��{J�wb��UC��;T�!�. *����o�Q���+DmuD�gPE�<俐�Ш��9�mڶ{���o��X��Y�~��En���/8Nk���:iEqKD:,��X~��G�7���>�O��N�sDb�m(��G>_]�FU��x��Wq�a3q���l�?�7��1��p����㨣G�압AΉ7��B`ЕØ���	�Dʰq�]�Y�䢐��"��V��Ov5w�WY��B�C�Ca��S׃���ˍ(++��"v�1T� aj'B��Z���r�&�9���*o�,����y
q�2�F�U�솝=��b�=����q�r�zT����Gi�(M�C�-y_2CyC(���%�S`K�)i��M{ED���zQ�.rY��=�U���a���?n��Ʃ�g�����{���D4_�<�a�u �}��\̌���9�3$-��_���|&N��t�[+����g����7���=�vb�ѵh��@o\�s]!�e���ա��O�Cr/�iz ����S��b�ן{�)x�o��,#n���j�}�y�TM�9/6Z�y$B˸�h�a�H�7��C�͊�%4��k3d;eb@2�>I1g(v�B��=�%s�C�?�?oބ����)�������3SW��[�[VY� ���i�f�`"�8s	9���")�]�ȴD���;�b�)'+�%�R�S�D��R�?�R�J֡m�j,8�x|��F��a�(A��X�;�7�R�����A�t�pgH�[��[����#n���9e(B�t�&�3�Ð�S�ڡ���g�t�^jH3��#�n���;4�U$2�'�35roi���	|bT���˙,���c�Hu��c��"H�32���ℇ�ǋJ�Z��C�`L�։�u8��ִU�W�s�/��Eg�釟�M�_"�t��z���=��gw⒣`Li�Ԓw��,*y�J�Bhj���u�I��+p�,B_�.�}�	x{�'7�-�O��C+]8��rQ��|�E&E��Q�?���i`��a���T��%�����ry��dyؘ���I�œd�v|�ŏ�o�q�H����r�I�0L�Ar:�刈gQ-!,^����R9H�\�2������.Qa�C����o*�]B��s�$i΀�_K��(KA�bPz�bX/���2�1���n�Ö]b��+���%�����	`�Ֆ������F��ڱ�~�	�~%����#���a�����/9��J%�	ԍ�C�}�P����T}�EX0��}G0c�;>��+8�L���c��8�!�)Ǔ�?�"�
_��Ϩbݦ�?�#�C8�����b %�v�q���bP���W痭���sʰFR%�\�e_��3构��/�m�]�G}P�=�2	w�^'?�hŦXlTxs��o֙%�6�4�lAOB�@N?q&>��3���éMQ��a�=&`(�Duu��i�n!�<��xa�}�{M�i����p6�h�g_}��5����w��b�$�Z��=W�p5��3O>�"n��O��	p����?�@_/���at��BEbr����߂���$�iW�iS&�}��s{���۴i��B��}�H�S��P����C|�O�X��Ľ����N9]M�p����e���e�89;�{4jBF:3Ut��w���UU�2��Wປ���n���͘!f�8̥}(Ko��Ѵu��1����O��6l4饝�d9��ò��0y�	dp���po'�j+��Ѯ�NIy�p�"���[D�$a��5��9'/��_�X�?ѐ��y[�[���]��"^�p8~\�F��]��LQ��,���n-����ےV�<�'�������ϖ�3��Ǎ¾ǠU��`"�)J/�p�>�"��~Ŋ6�7?�A]}=������W�(�� j++1����I�d�~�y��y�%����Vᮇŵ�;O��8N����E�������gH�>��l�JZ��+�UG�W�x��:U�N�OvH����YQ!�y��fPOBȧ_|Q1^fpȄ���a9p�a�	�"��e�P�'Ie��$J��G ��?
�xY�&2t&������g�2[R�~-��|���#���P~�svI{�~	�riAYf��'�˾1:���z�YGLQ�|����2,t汣����J.Y�Q{�ˢ`R"��^x/<19ȗ�� �5C���j���%k�ToA��F�+bA��9���G��5W]���-b�+1�Õ��V*�UG+��K��#���HD�Q���&y�K�ұ���
TF%E�1�õP�h��Dj�n�ф�����Z����'�
eQ����񷛮Ց}v7��;���uI�ŤF	��;�eUuz�fRL'K�u����ҋe���t��L���55�����q�b���M�M1=kx2h���c/���/�X;�ӧ�¾U�P�9)+������E.������W�#��x���}��:U<��:B���-�ʭ��7n�ۋ>�W���`�5���k��#�R#~��4�Ս�u��XOG�:
��/�^ۻ$�e�|��i�BҔ���77a��f��������㯼��.\�Aɥ$:Ł����5�? ��>���K�B��o�>��Ͻ���_����_�в��H�E
vu^x�	y#�N�=��S�/^~�-s�ab4F���{	M�0Pf&c$��|���#At�,���-��T��r<��38���J�P({}4��g��iO�m���-�F~��ZJ�Pc+��?�yg���E�DΦ�%���g&?~������$�N�!%��%�o��a�䒛6�Cy�\�T�� F��#x����Z���;��wAst�l<���8��Y(��0 )A��Fl��ɲ֟}�v�����\�{(�Կ��'!$� Aq̏=n:cY�e/775�9X/�;j�,E���/���Ԇ/��&��Q�-߃��^M��&U�����#�
�=���Δ� �����񷫯@V�֍[u������;���ri�|�AK�� �,�S�j��'��.�[�r�o�F���a����n��/�F���"m
Vœ$�G%��wދ[�z�
}Q��)iQsK�B⩹sǝwK4\�C��Kl����_QS���{���������J�Q-�˯B����MF͐!ӕXފ�xϚ�u�V1�5Օ�'xʪT�kSS���K�j�L�m�*�;.��p�Қ	q8�,X��H���ǟ�O��O��.��k}�)+����U�F�f���N$QQ^-�<"g-��Ũ��e�$f!�Uz^J����շ�W�`���%�kQU�=r�|�Y\r�ɱCb���378�F�5���a9���H��p(�8Aari_|k�?�P$%$rI��i�~y@��l+S��y����$�@�/��O��3��kT{+���߮\�"Ov�G)�x!��Egw���~��E�g�=��q9L�J�ۦu�$�hQ�S���K�v4�vj��$�F�����9��yKI�8������k���L
۪f`��������B��^b!
���P�B�j���%�e[��l���Z)LM�`E-^~�C̗4��0iǨ8�˲-�=����=^o)��rP��%9�L�U�>���5�d�ظy������e#{6����}a�y8���� �O:Q#��ۛ1���ښ���+�ҌP��
IwyAh0����<E�7��CO?�1��Q.S�Uъ��������EwM_���1�fy������e�im9ƌ��ؐFl�]ʬ?6�*Yo~)�2� �qM�;�(K�����0A�~����*����k��D`c�ʤ�܌�ha1S0��EcC�oذ^�y�r6���͖>u��V�����S��2mu�I�H#^C�u�1�^�y�$#�����*{ʚ�=?���rȕ���7Cbl#�SS��K��y�-�T�m/������y�J?�Q
�y�����{�9T�5�e�J��H�?1,a�ʫj̈́@a7�NQ�2������{p�����UzD�d@6����Ҡ��V�l3�㥕����~mѧ�(��Q��A `�}l�CBj{��Y�S>����
��h1R9�ؕ�i;�
[9�(��'��0���}}zY�����L[��V��J�E��Ĉ*��ݨ��̌�n$U�N��s���o�'�`K�A
�r T�`���' c7NixO9/$��їCv[��G�Z7�Z8�Fc�LfT�D�b1j���iY�@�H���W�pWUЋj4�_���\�(yH��)~�D�Z�ꗦa-w!�� �h:u�˕�����|w��IpɅ����>�L�M7�_�Q��CY�X!>&>�0�8]��<'�Un����G�_�9/RA��Sy:�Ŭ��e�v�R
�$�<g�D5-�׈7���O��g��F^B�u��d����T� �:'����v�*���V:NO���$iG�pJ�u%���E@"莁�����p�s��I�M]3�[H�hX��|�������g�AG�G��i����$�����a��@N9k�e�ցgF�J�47�xMS�jf�
y3OoQ��´�	V��%)�#�mF	�LD�Cl�ʁj�ҙ~9��B��ݦ�X�MQ^��G��Z�����6^���C��e��Ć��g7c�~����b�X����"o�K��E[6d)����h�Rs�R=��TNB��pP��d��[R���u�a�(���\6�Zr�~���0f���0�R��_Ga80hLiP�b���2���$l.�6nzAM��*���jD�sT��K�f%��-i�F�]/�u7�C�xp����N��eux+M�!\�F�6FT��-���K¢�UVCX�ZuS�L�:/bS����Ou�Џ�0x��r�)�{#�m-�?ԛ!���AE�ZJ�Nco"�v�,%b'~�/zΒUѠ��%��nҤݓ�(Q�J$6��u�X~wXR���YN�r��� Ϫ�,z�ͥ�K�E���
��t��
=(X���s.�7Fg����F?�5�����4�Ԕ��6��q)�h�n�E�H�`U�eA#:��.�΢�Z��+�ն,Ŷ2�m	 �25��UeUC��E�)吶|�����w�����C~����D2�uʛp	F5i���Ezu��i/�f7R��+E�a��+�M�he�v�*���D�9ӌ_��Ō��6f��xMs ��u`ii�X%g�	�J׍�2Ki�yY(U-�8��� ̳�,�'�ǰF���D'o<,�,S���J~*�[�@����	(	��1��U�'��I��C�:��h�׈oa!�\2�h���a���Lu;l��I�Mrx@��		'Y��ER��	cN�C�f?(A�2� *GGA+ݹd\[�N	��5����})1V���/�TǄe�EP7�8ӕH��i�	qV�;��.�s�E��p�0��m�F�7�8����Q2�y�f�<��3������I*��]��`?����ҵ�?�����b���2�}H����t���Z3�U=���2�1M!{�����p�d��
�H��Y�`�[�DrD%��8ޟVd,j�lB�zP��au�&R�h�b<BQ��$�O�\�|�QD�Q�&Z���yI�������kT^4�JPd��>��G���e��r�l9lm�@eU���B�]Ke�J!�ʁ�=ln��ڌ��NP����Ơ����˯��WÞ%@��$�4{&K���H#�X�I�����:-
u0b��Y%iqh7��9�bhֻƇd�J/ ���/Hv��k?�\B�l֡��A�\�<�&5���%�H#"M�����1q9�a�XI9�,2�%w+����0h�Vɰ�^�`.��ϩ��O�ڪ
��	I��H��� �|\�p��lܨ��x�������G���эj�y��+�����}�H���v�޳A���J�	���=M�X")�d��}	�w���&Y���C�yLX[�&��p���g�d0]�����_���x�p�9���ɤ\��bFb�8�S���J�b�+���?�^��2�����9'�SCjS!dvZ�5Gv(b�>��A�l�b	|��rt���#<w�)�\<Q'n��BrQΟ?-m-�<�D�صs�Z��}��E�I%��?���&cq�n�|T����oF��R=Y����98�Mj��V�Fv5Nos��,���Cr�W����!��q���N�el�+OjI�MSv14��N�8x
�=l��nA9E�'I�H%��uW_��ĉ&-�k!˝��U�/�F]؏yg��Ά����ڂ��_z+����Y���+HN�]�yd7$6����*9�a}�������!-��_�q��'"�)�J�ҁ���z[��s� #w��u�'j�D�>� ���5��5�$�T�K�S��)N^�Ǟ|���~E:9���۳�@kL#���³�! ތ�6'�{��?$��o��!�)�֥<��D�gbpj�A�9�=�Dp�(���4��ߗ��u�CCD�CӴ�������2�>�p�{�ffE�c���H���g_yi�WјJ�V0�^,\�YZq��9�����0�$+y'��^y�C�Q���(
G�M�������"�ɳ8����hU`?��]�?���F*ѫU�Z���,*��Ƅ�8d�	
�Ƿ�qpY%D,P?� ����"�2�S�7%��}K'���c�ɳe�{P��j[9㲠Z��:,i��oV��?R�$6�Rt�ܖ-\Kb'1�\\B[����ƏAWg�N�6{}�E�*�������#{N�'��O:#*���t����bF�^.<s.~��qH:��gg�F�]���x~���-�5�_>��1g]�ً�=[�B�Ն����7�����q>�_q��(��v/S�Q��7^�G�v���W���P�=kF)�{���oOL�w����1r\#ں�T���CcY��k7i�`�V�v���w�8x���Ed�R�D"�j�����6\��[P�َbQ��H@d��h#���3��_"$���*2:�s�x�'{�PWnޮ�m�8	|X�����^��v�¤�c��5���+�(\�������B]�(=�K��,�u�7]�����Ï��:����U%�kڊ��]9��Ck
��19t	\��d<��{��W"��ᴶ�84���8c�	ڦc=�['RQ��h����p�e��o���Ʊ��VU�2��"\�,�;�9�CC��3|��
bbh���j�!{�l�, /�V��@���p��=rx�(:�Z +'�|^����
�z�)�*�U��ϠN[A.�.���9�koŸ)��%=�l"+��%��?g�D������!q5��E�o��1U!����"a�_�x�@��Qi�w�ix@�蔙Z�9�!k^U�qG�\���v�"&�[6ۯ���x�s���#Ͼ`R"�O��1ԅ{��[d����S��{�U�c���:����1�G�᧟�$(J�KC�X���)
��VV�jŜ�ͺBHm�=z.��r�k4�z�
-��{1s��8�f��C�<�P0�޸��F"�>\p�<,^�%~޾K�Y�&N�%7o��Ux�$�ءR�e�h�� ��`���g�}����AȢͯPvM��<��5᲋X}�(�F��=�=�Z�����V�v�����[�K˔��*{���>����f����&��@Ήo�n�S���^�D�S��[���˾�'U�M.U·�UFp��)J�W]=*���_,Ô����p`W�6P�ދ���rԏ�C�Q;Bb��b���%jУ��7������Fmy9N?i]���S��F��w�b�v�>���!ή���/W#!|t��޳��,]a�:�H���b;Q&��������߀hy���h0�����O�5���?�g�}MY�Ə����OƉ'%F$A�(�����I�dw�4,L��&���?��>������	*�"%���DM���Bv�'��0bD��^a�6R�ܹ��R<��kp�4��(JTQ��YG��$�B�uX�j5�	�/?w�>��u��9����S1�*�dg�"ޭ��W^z����~z�s���?^WW���=]�y�{�q�����a��c6�/a� �;�T�XO��*G��'_�иu��1s&�Ve�:l�d�~\��m�r��&ؐ�`�~{�>E|H<B8���f��]���{���M���\�����b�f"Z4����p��3�δ�~�$�X�-�C�Kj��4�<\p�|���w��t�x�Ut��?���W�E�pí�H�ӫc��-8L��!��$��s���	���r��ؙ�5Ҍœ9f�[�)���4���f�VU!1Ѝ����/�ݏ<W؅Ik��a̜~ k�t�ggK'��MR4%���1e��H��a
w����`�bTS̩) ��Cwߎ�� *��-��{�rǃH�r�]�?�㯣�D�G�8�}�#자&��t���.Ԕ�%id�;��_~�Y�#����n����e�<t?���V�A���1�5~$�>c.�{������#碬<����}�L����BTF�P1�k�:�C�]�E睍ۛ0aơXp�e�n�R�OZ��1���K%J�c��������O�
IPPֺ�n������8y���圌�֫���O�P���}'*�w��o/�B�QPŘz��q�W����.��O�$픔$ނ��y��m��7^-Y$I��c�>_��^kb۸��?���h�7ߎ�r�G�iT�6 ���oW*�������}�#9�8d#N>�0�:�X��:q֜9x��7џ�jh�����30����HZv׿��֦V$�d�����^��߭:�Ϙ�/��Y�v�@0L�?�4��X�M��쪛4��c�6m�58���b��;��x˿$\j��FJ,�_$�J'tRu�/��3�Tm��v[k��x=���"�}a�-��k��X���=6�9�@�X���P�P�/�3�����b���y��̣0u��5b�u��で%��"^�x�t6�])���k6J*�D���Htr�Q����L�iE�d�n�[q��)��E_k�N=��z^z�~�s��S>��/X�Q�x�0�w�X�y�fI�.sN<^�؃�,N��x۽�����������c���8`�TH�)�V�Q(Fs��מ�M�����^��JFt���W���/9�~D�n�Յ)�Oƺ�Z��$��s�=�'�(�g��mW���$uy���$m���n��Y�Sf�;y
�%�P'q��%,OJ�n�'_-Ǜ�-�T��0/^����r�$�9�r���� R_��EN�V��d\Źg]�p$��Ǧu+B��r˿�k��8[�Gu4}������q�E�ٺ#'��O���ѣ�9f�`oN)�W�x[�Bȶ���j���'��:�32v�8���|Ĳ6��Cڵ�����O�?�?)��r�{QW]�x v�HaP.�^Bmtv�aѲ5:%�t�B�SXy�'�	�_�I������)2�;�N5TW��n�G�~����\�D�, �p��ރ�?oĤ1�$�<,}��Ds~1I4�W���J�=�\�h�H.9�I���|N>���lډw}&j�?Z�iʢO����N��"��r9�\�)җK�5n�HW&����?Bk�0|eU�Xe��%ULKJ�lԥ�6����~#��`A�t�x�����9D$��'3�K�����5���W٩#�	v1��!�C�|��|_y}	�rC՟5�1Td�p�2�9�x�#+�D}��S�j17���_D��D�b3EF���~�{O�S���hJP*>rJS�%�p�azY��а�neG�/a��7v*�}��2U���X�8Bz_~�Y�
�$�Dcv��O�O����S�BL��L��~Xo�L1]��5��FD��Z�c�?#�L�Ҳo��A��Q�oG���+s�Ek1I�jq�巈�i�=f�N�?��z�:a[IDh�I'pYq'��ڞ�u�o������D*�--/{��:�����O�'�\=�Ԑh�av��N,U]]/��.MM�_i��Qo�֒Oq����qKHT7���bX.��t��ò��<�2��bL�(m�2oWK���8��/>WVՎ���"�Ł;���p(�Ͽ�RH#�2V��F���J����#n�b �)8�$y+n��x�ʺ1JK�#k͂2CR�<W�l�)I[j�����=ۺ,�k++��S�ï~�p�t"	��(�_�~9'_����s:=��k���(zP��Zy�hU=bb8�.
6�%ʷ�%Nh�W�c��J:���m�UI��RI��c�.�iz-F�������́O{O\����r�9�F"w8 ��D��K��'���ZҎ�^Y��J���`w��N�l���ʋ���>7�O���:��`l�e����`��9��"Q��J��j̘>Ei�?[��tn�"���6����0S�D\:�
�����]�Ćb�+/;������LI�ܡ\\yI/Gh�E�V��y�d��6G���SS��V�6r�VH�����iC����bV1,�����-�VD�G
�&����c���hN/~�Mv*��a��h3'S�nي�S�ԙ�����ȦݪU��:�Ő����rٵE��.�P�E_s���X V�]SS�hI�Ϧϯ����$�+o��%ʠB<�IX
i5عTFuWhH��˾�5��Y[�������\�2�!���,��q��K'$�[��K(�(��%�1�z+f�*����H�4��۷�l��w��P�c�" �kIm

�3�d���	I�|���� �:�W�""��Im�3b$��F��ce��V�g����j���a�*6�lEU�X�9]6C�]��c�Ic���;e�%R�S��Q�.�b#?��y�.@����(��NY_o��󞲝�$L��ml#3M"�B�DЫ"OWV�8o�zԠa'@M�7.�X��2R�3]'#�BeEX�H���$p���u���J[�.��v�t0?��\���Vp�H�V��@�d2�S�G��������h�v�â*�|@k
�ry1�K��~0�.���G���F���y;C�j�	�H��ϩF�7����]i(f�&�ۃ��>44NĶ�m��$}*(!��er������`��[.�]���*I��Q�ZY���8TF�����noR���LJ��#I�� �e���P\(�A�VO��?���+c��R0z#���AK�abk�G����B�J��h��� �vi\��Q���_�H�re��#*���Me0%�
�ya�J�R_Y��1-$;�����b�'��1���8I�#V�d�,��l�~m��8p�<G^�r��ȅ�"�����li;����Cj�6�W��k8E`�W8^��6#g&87ğ%Y����)d��mB"ɐ�dMh��t������a�V�p�*k�a�\���Ϋ����=�n��KI�#S%gu����U���D�h�"�^�DA)	8V��L˔�U�gj8�i�����|]��R6,%Qؠ�w1�J����qj�E-U<2�<� Qu׮&L?
;�Rr_�1��p�U��؄�����"0Z�fq��N�#�z�j݁C�,i�*IM�j��$��K*:I�ny���z\6ū�e���w`�ĉȧ�CQ	��F�M�T��ȡh=�	1xiy�u���5� ��<�~b�%!�AD�Y�bx�P�ﱺ܏(uB$:(���Ǯ����_.iM}�����a��֞�d#g��rxe�3r����Fkg
vθrZ$�Yr�{�F�rR5U���E!{/Z�y���X���ɡ����䗟�x��;�L�Znz`���z�˰ �&���rY�Ց��eJ�Iu���~U&g{��;�)�:(C�#S��ǂ!	A����>X�1I�l�*��
�E�wco���b��C���ɝ�j����#µ"����5�1b�4�jCeS�/ə)�(^5��G��QrҖ�8�st&V�R7�Z��Am%180ԯ�A�HrZذ*�#�9���bۄ�y�Zw�`�M)�y��
n�v|��P.�l��ѺvzHgHk$�ʭB(wO{r*:EJBy�^���A��rIK��0]�d%�PW��*�<��ɳy�R��{�ƒH��:[Z����-ۛ�{th�J�P!����Xx�uzt^5�ެij�V���t�QW��e�gd6w�!�ꠜ#!��^�:�0�J��rxOT��A �e
�^���oLvvK���$-�w��iS������p2��dr�b����&g����9�<��v sr��m��b��˞JJ�R5�ak�`�{�_[]�q�j|��cDe��)���f�qО�8��iJ�H�c�re�c��g|���p��%3؎[n����°$`�o@�g �^y�2��C����U.��b:4F}ا�J�h	��9��pY]Z�*n
��V��F�D`��p��EI��*��c�q3�~�*mQz�^��Ȓu�G>c̨z��_�"P���D.����==��N<�M�Q^S���/�+\��,O �K���*9������!���F�M��I���D"����ܬ�LM���X��8�D�$��u�QX��w���s S�]����L�ܰO[�@�zl�C��}�=r��*�>6}���d��x�.�ˆWH�0�v��xqq�_�^e@5ri���~��jg�8�_��J篒��!k�؉�3���'�|��Ͽ��R��{��7��s�ᴓ���=��
L
xhon�)'� �C.�x�X���� #C���\�X7���<���#� ��99���h�Qcᕨ!K#({�IR��
s,҉m�m���c�8{�1x�Ű�a���DVVZ>{���IZ1�`�d����1�?^�.8�,5󎙁W$UKQ?
��,ڦq�ɳT��bsc˦-��Tɿ�WfqZuR5'Oe��8^{�#Tɥa1�}�)z��b��[��_�/����69�?�\�1#OD{K�;l:B+�ổ�5�c��3�#��VT��3�g@Y$����nc�q(���p�ygc�GK�h�"�9��v⤙�`�	c� W�}����6�b����n�Պ=FU�/���^��r�W��#�p�p�� cS�u�֣����,�LR̻x���Z�q����m����*I��ʣ$�봹e��i��E^�H8Z����3~�9qTz����Sx G�9����;У|��c? /��.j*F�A,�-�p�!�$�N����<�ʪF���%��F_���0 ~��i��ǟbGo�T֠w�'u�V�{S����3��W�GY���!��c�x�*ɹ���3���O�Q�\��Z��/8m�������W
6���`��݉3O9Y�س�;�o؂u�~������*mY�,���9k�� '"' �}%㠱�dC,8{މ�^��*��P~ڴ�.�..�ƒ�^Sz>���ŋR������E�����n=m,_��==�ˁ�TU�c8Xk==޿����Q�(B�x�����O=�h���Sx�)dd}���:�x3��
`��͊��T���a���/���i�՛���+��֎+V`�x�����۷��a$��bxw�gp����� �'�>�$�[0O��	�_r^CD)ֱ���D�����-�ƭw�'�VkQE���,��{�VV�*�D�DU�,��O��mr��5��qNT��xށ���ۊ`�\E��B\><��8��3еsΚ{��}����]�T���Ӂ��=���I��W�G:���r��ȓ��%�c�ۯ�B��.�
y$B�&K�[�U5���&&�8�֮�۲c$juJd1m��8��K��yXR�8��֬�ſ�q�S,R�,����\{����jL_�yߍA1">yn���7�tc�'K���P"��]��
Ͻ�:n��:M�Cr9e=��{�B퉪uy�Z ��/e��)ғr�v�9p��ុn��og؃��~���I�~��-���g����d9�N�#*��y��⹧���P��](��Q����*}�TΆX�+.:�-�Z����j�}(v�؁�q�௷�"�C��|dp�޴x�}�/8]�G'N<�PU?':��4Q]m-:��/*ѮU��:}GO�����=u����鳏�\���K�;�lPV�>^*QB���	n!F�UDvk�Y��5�d����Af���n�Y�=}A�T��ϗ�gE��C<�ܤ�a�fxr�=f\��c,�?},z�Ȧf�V���S�?g�J��2��EkO<�
.��x���|ġ����B�x��.�����A�WS���;T߭X�}�'iZg�9^5[9��&)	�J��
,���ݴMF��^�a{�����h�5w�x�!IG�8p����S$�FR��7m��u���U(�B����'��1h�����{�|�!$dݜV��������\�\Y��Xr��NDG��h1��~��'�%�<pox~s�6"F�b)����~A(��7�E����O������S�Q�u��ݦ�$����X���rYCZ�3�jf��[7�?�n���òCή��V�}[�2�����s���e���t�l~�DHK1a�H�%iL~x}4�Cq%^"�k&?�$R$��ԤPRzסBqd#{���p�e���ݢk��H����V��.�#!���&S�tF9^o���z�	�~��K�Ė.9T:{��ؾs'��.ӽc]��e"�Y���z�t����i�]1RC�������O?�rEi�)��&�G�e݈���p�C��xCb�2����,��"��G�>�$��x�K��|n��$B�������l?qz�Fb�8�,�s�y�|�r��e�c��d���{�Ҭ����G;���:N���~��>��n9�I}��v%�oݥc*#9��9��ƨS«��xN?er���$i�X�hE6�A{�R8�a��Ճ����
:t�V��g�P� 
���S۳������FY�,e�\�+���@�xŇ�x����*���ߏ��ݛ�p�oچ��Aŋ8346C�2N�a\�a��b'﷯^R��:�$���ү�����Zmg���/���mw�4T}�'8�#���y����_��\�V�Y0Ek�;lNT���S�c�9�R~������-�v|���ʹ��8��ڮ�.y$7����?)��&����LA55�z��n���M�g�����*:l�H�'\���?�ܹs�5,)��^����K>�FNX98�GxC� y�7�<�ݏ=�æM���#��ޅ4��t�\h���	���^yӶj�����S��K��e��������-���Kf�4>o$%�H�ig9�d��?�c���a�]�c����4�h���7H���)���-rRZ�/,Q��~���Օ��v�^$�o���GK>�3�Wz^��D��`mʡ"+蕈�ko��fk���0�6�l�)ri�NiK�#�����ˮR���.�����_���>�3���|sظ|��m�%^�P�WgL-ª_V}I��5�HO��*Ǝn��"��o� ���HEY`C�_�U�� �΢B�߭܀�뷠��]�%���o�c�O<���E�ڸN�6O�=����+o#�s����1q���y"T�2�I�8UY��p��_��~�&g`�N�*���-����a9�$#|^�L� �sIYrbX��.�����:x�ux���1�n|���͜Ci�$�=ɭm��D���\��)=:�j�! D!�'��Z
�u.[~�.��y ���{��Q�$ȩ8���SS4�~:�efWr3����-Q�c/���y�I�[�}"NYy%���c��fV3��c�Vm�e�.��܂/��Q�Z<�3��8��"�-j�l0S��_�1;i��J�賯h+�ғ:E*F����ьj��b�*F�֋���dK��Y�]����a$aeA�����Fe�������h���� �?�iW����$-"<5p��;X�PB蜒:�7�/�����N�O.a�l��N#S�X�I���g�&d�����ˢ��v�f�ZK�F�ͥ��o$s�:ς`Zvw�
N�Hə������A��Qn�|�D�>R5�ľ2%J	k�^���/�D �����pF�b\3�E���pH�{�@����zz�N����Ý͕B,�q�l���
?	v(����K�m��M�Ei.�ӧ�.-���6�"�
#�h1sSj����1�CjɤLGIE�94감�ޢ[^����5(,t���\ވF.pH"%�ס������DaQ�]ւ!g���]@[�,�f��MCU��%k���(�����#��%��H�R��I��d2��l�j<��:dƎKA��f���ٕ��li�]D���S3�kG�[����ҨyI:�D[�Ã��Ӝ��:���M��Y��Xw:I�y�4="l-�kTԈj�C������ ѠO��%+�FǕ��"�["/z*_I���5�΍��d�����9x�#��++u`�h8G$�ߗ��'�C�d?(����X>;O���)/��Z���g>���9@H��[��v8~5�ʁAt2`�}t�̜�<�Y.��6{Q��x��Y|��8IH�C�C�8Z(p���6��e����B�0v�r3�	C���3$���Ѐ���X�/�^�������Ɍ��8y1�䡑ˣl�b�(ɫ�,(�	9:�:�m ~*e1�#_������PU�F��s2�Q`�0���Iu&��S,�yu *�aI�Ĳd���r��&�(t���YiC!��X���$>H�JV�v(WR���[��b���}A���d��]�jY֪���n䆍�:���XXWф�L�xxx��j�&��R��X���Yٯ�h���s���ɭ�)���LZ�I�"E���ߧ�g�Cb+*����(1ly��2��qYDָ��� ( �Zе�"��"����x�:�<N���/.�&��I,�CV0�5�y������ᾐk��_,�K��Rz��F]J&CZ��=b���kA�̌R鹑Hh�c��AC%�/O����jIO�j�
J����;�f���3�[.��J��9+�
��*�0%�,���E��g�� b<I;�����S~?+�:�����L%�F���K㖕���5�ۅ�ݤ���?�I���Q��L��m:���c�p���Fn��a���O��*���J0YZ��2���1ԓ�ls�yJ�vf*�7���ï�Lą0 ���6�ץ9�M*�F�D���]#V�΃F�nM#A
<�Ga	�x����s�6q�9� .:ܚ��J��D��ȪӿY���z:���R�Fc�(�[Qf�c
vr���Diϔ�h��PFe�E����V���!�H}Fr�|����r��>�d��OX(�W���4LP��� &5$�i!�0eĚR�Y�+�����j Onz�C�jh4R�%�"�Z9�0���f���|�<R}��w�c������krȓC�%�����LP""����$w�K��Aa�"�JqP����<���=�����Ԇ#���02r��C�J@�	޺:�$M,W���[��+��H8yȇ�d��
}
)fH�u�NE��H��Ң�^0�"2$��&88h�����'iTɿS�g�M�ȝ�ұ]�Q,�A
$�O�ġOU�k��$=�(ӏ�R�@*����I�C�0�Vm�t��8܎=&L@yy�[�4գ���da{��^�qE
D�ȬfD�^��zS����~���r��P�vdǢ��F�������3�jo|��9�>yo��>�(GnJ��U+5��X�X�V��Sy�!G��"��u���T0*ux�kW+��!�Ħ���8f�a�S��b��L�F{q�9g��<���~�Z=z��F�����$�b�<��p8��)hg�i�$H(�zq�g`̨��)�S&������?�G˾��T)�С��(�5e��e�����+Q�W֠y�1���Jj���<��㰗�3�9�8�d���E�v��˯��@��X\�	U�ƍ�KDґc��q�F *��с�0ǲ��q�|�b�����kZ(Q͙�"=�PO7����ps%���]Z?��{䉧��Tィ�ba��j�K��mߎ?��<TTV��y'F���R��K��k֮�$զ��(J��!��ebYS��'�C���xA	f���+�km���Q��(ȳ3�Ɉ��X���{��X�~²���n��f|��rm�8Eb��2��|L$�q����٫"NϚ�(�ER��֍��c��䂵P�dԓA��'9��M�Q��Z&Q�y��"��T�90K�Q4���dF�1cځ��32*`{0̔A�Q}m����pk�j�HĢծ�ApYOG�D
���5k֬A}}�z�#gL�]?��LI�T��!�����r)Z�q�Ǣ��J���Q9I�nl��@?�liò+Q�K��ؒ2�&i��R61�C8sΩU_����������<���+�E�F%��S]��I�#F�R���\�];��qd#�q$cCjtgL��?���鼮1����vm��{pǍW����u#4������(�|���O��_���~�
oeZ�Ք�n���*�P&kT��+���L�B��y�!\��K� NE��n�F΀q�۷�ƫ/SIS���(�s�Zv���;�[�\�Y14�̥��̣���?���'�+�>��DY~�S�#+�p��þ��9��߫�|Q}؍�o����#�G[��^�*& �#�p}����]�8o�g��>c�+u��� ZQ�ş}%+,��A�)�<�������-���� �ף�����b�$�E���\����j�YHdo��v�\�����,�|��V=��@$���BWOj#^����o~�(�ө闦MLi$���k�����Dw�!��$�8VG������\��q�jG)��MU�r
�qX�w(�<��XR�ӯ���
T��\-a^Dz/�X�NM�T������;>s���!H��ax��:%��V����ᾇ�E9�b��"5
נ�6�5Q�c�k}��R�b����?�$<���ڮ$l����$Yh�w��*ñG�@r`P���V	���x��^Ԗ��3N��ϼ$�k�*rD�'�qh��W�a!�D�Bȉ���~:�VH����+~�[���(�W��ųne������
8+��u�c�t1tH]T�@lŮk���ڊ���zQ�F�;1E)Ab`�a�����������w�*0�<�?�^��j�%��!^5�����:���Ė��`� &��������,` ��6��T������xmc��RhkS3�QJwJ���#܃o����K$�s^�Hr�f^r�o�
��x�lTBEKBø.y�k.�Ͻ��J&f��ޓ�&x0��ށ��!�"T1IA�9"$�R��,�=�:<�����O;��z������x[�q����!����p�Q�L�{
�^~�:!��1�N�M���%�|�V,q�b�Â4˪���D.�����-�E����ꖖ���Y����r����ZlA}����b��z^���'��[�p�⺜\�%���q�}sv�A�e1eS}�3���ŭ,I1[�K��M�WB�1Æ"�R=���1vRޑC����\w5�%~bf=(ޞ���޴h�Esc=.8�t����ȇ]jڋ�ۋ��������w��ƶ�aqj����TG�3��K����O
�`�b�Z~��G���U���I�h<ŀY�pě��}�A�|�=�{*m �+y&-8�*K��-����v��q8����Gp�1Gc��u���m��T���.\(��0é����c�J��>T�1+�����~1^�s^]��ZW'�����W�G9B��*��ֆ&��|�*�M�8�`3K�p�i'��Ͽո��\&ϙ3*/��P ���b�e���������G�E2�)݅�μ�-� .o��e�R&�6��M��K���_��
��Q�f���(��mx��;q�O�9+B"��s@�v��Ǩ·����>��v�fp��OɻI��ѣ����M0�|��H���kB)�L�t^�Iu5���۶���qƌ}p�{i�}(O=� n��~xK�t/��=�&q�M��Z��0�~�n��)�?l,f^v2�i�]����������jk&���q��w�r�;�Q:j<�y�{|p㽊��
�:���0v8�(�:qх���+�L�e-گ�a~q0���e������W�1cFc�쫑a(a���Õ��YgV�@½�x��;��y &}Y;���M�*�s����i�y�)H�zp��[q�e���(�=L��}�->b�d/[�'��}	1�(-���oc�	�I�x���%uc��/H̶UQv�������A���7]�G�=#�â�	�3%�}����!���t֊���L��NL�0��|���~鞓��x��6
��k��ˮ�y�<pT��"��5�s�\eҦ�ˈ�r\�epGj����,�q�}�=Y��|�x�i�uU��{_<��[�c�Z��v��t�4L7J�e��G����S�h=v&%S8�c����J�����d���M��ݧL��� �����K�ˢ�$L�&a�Ig� .�Xq9���8�E����g,X[߈�O>|���V�.xK㗈2�(�"������"�@�H�lw̹�vkM�2�̼H��|>@.�������:�<J�{]m�#ԍ��[n{mrP��rJ���W�c�A��:X�W/�>�`����ZF�
������g�H�S��Ja֕�K(��
��_����O�g�qÆ�F�놼�:�\��$F:�JAA�@%f��6��>��ȼ�p��W)������N�g?/W2#&�(:<��J�=�2\t孲�N����Y���GX�n-�8�x��Y�z�Q�S�٤CkY���N?�@�
��w�y�Mb�혼z�_{�K�K�}�Iǈ�@O�}�t,[�IG��Z�1���� ��b�x\|�b$��y�dk�N�<�><pϭ�gb:	z��g��ǞE�4�Y.?�,����)-|a1���Kc��A6v��ɧ_ƕ���h��ċ��<��"9�c��d)� ��-x�����+�׳������Ko���c@&aK��b@�ʌ ڐ̮ ���zBeb�����u�u�L?S'���͸B���E�%�tHHً�'M�3�-H�s}I�Gi'>1y��҉U7J�;�{�<����`r:��Wc7f^w'�~�n��}��A��+�!*F*ƌ#G"��<��-;������lX���|��/x���S��+���`|��R�)���\b#�ˮ�Pz�y�Wz5�,u?{�3�u�����¦$��o�I�ܕW�Tf�Ǐ-��P�{�θx� B�sx��%�"�s��܄q��~K�����ۥJ�p"mv�Ͼh]��YSX��C��|���4 !�Y�R����DCu�I^|ml��RZS�i�n�(1퇟|�iS�T�r���`��!8���nN�v�p�z��p=�=H�}2R��zV����-�<��Y��z�����8>��������S�z�;T�_��2�PAU��)q.	k����;�}��JYm���jˇ m�5��x�Y��5k0��L�d:f�9Fν��E���Q#q����;��Ǵl�%K}ފG�z�w��a��| �#/��Ii	��%b���߳��d�]�q��j�ŝcz���dVB����8�I�T�)Fk8��	�E!�U�Z��lT��v���\g� �5���?���>1���L�7�4�g�Yg�V��cN��≅O�;nT&7��B���Xy������b>~*~Y���]%
f�/�x��_{�|L�UD��L�k?�ը�����y��G`�02kvi��V�8~_Y���X��xq\�"C&��(2��O�CYE��uZ��r���lVTU��7a��s$�iUD��ظ�.�s�<����(2ɾm�F�Z2�bן}�9��:ֿ�z��{ű$�%E��~�|�D.�^p������bq��\n6�Ț���.�h��!���������c�ÏKy=Z�:��R�(��7?�bi8ɪdu��~G��E�\Kܖ�Cٛ�*�����*��'��@�bJ<�S;��]�:�	4�dq�1�ҫ5���.�u�5������EJ�9���9L��@$���"�t�#�k��D��2jrbs8������#ɜ��l��������X���]B	�\����3&���r�S5Ll�H��bBD<�[�9ٍ�-�;`׾ ���15���/_���M��%Y��Q�` .�"��\������Y�C`�f�);���w��?�b�Ic���`�=6�^�<+)*#H�3J���s"��B�C�nn�a��*��ks@2=((ˋ	%�z���uM�(g��AJ�׭Y�\�z�

B�:�:��K��O�M�)�/����ߐe���-;�N�\[������11b&�c^D?�a.���,��6m����(Ek#u�]*�H��cB����r�F""��Y�W���1�<{D��sT<������eO�r}8<�!��X��o��M*\�=�"C&�����z1��$��IаC�/��@Ό���@�%%0y�r7�>2�d���?#!�ˌ�pl�ʊ�$m�ë�T$Cj۱M�Qò&��
8�;�	91���$�MjK 9T�/[ntI[�l��P,'��"_�G���T��Mny^"�8{��AX�b��cI�˺-�|� w�hgg���1�`��5���׊&il�xխ�+l�8�].XR@O8�@�M͝����6���wS��������]Y��bͲb�l���$P�L��U�战�i�l�fevZ�z���&('5ڣ��7����փ��pJ�c��	fZeC�|�����a�@�x�M��8|���tl�!��Qސ���_:�Ғ�'��Cl�l8G���9J幒P��Xrc�n��ZYCw�19���F٨�� Ge��$�$�����c`�)���~1��X�d�Lf��5��h�č�&{GX���Bǧ�M����/��o�%�#�wRB2��mgP˳V����������24Mپ�T�a��ې��/^2*��\�Y��9��s^�&���7[]�Ύ&8K�:��a�B�h�*K{ť5ڰ�Կ�bȽb3$���5�ż���в�68�M%���c��=�[���)�U����,�M��]�R7ס�%�Dd��81��QK���D�|��'NP�	�Ɗ���Y��F���2?<b�9RBF��ݢ:15l�$Q4g�8�l'�����o��g��|�11�DTԑaKz�gj*J1�3�F]�P44w�{����7l�((��V�\p  ��_���,j+F)�e��VA#�}q�G�!uR8<Z]S��p,r1yϴDf��s� bS<+ٟ"f�c���\`��8k� J���w�Nm� VE� �xU
"�dCKZ������_��P_OX.�,D�][Q��X�s�ŉܤN
�I(�e+�X=	`X(�����+�8u'�� J�rZ6���J23R�usX6�R�y��(��8��D��Iȣ-۔r�w���Q(�o�L���(�$7�%�J��%�~Y����`�-̆�SR�u���4�C��׿�%d���L@9������5b@�*~�R����MI�᭒'��sI1�"6���(�d��\bH���A4�E��~��ě�%<��e�P�"(���Gj C�*�r���1����v�g��.GyS����
�cy�ƍ�Y�L����eS�)�A���w��8��ͭ����\�twr��R��2��L�����0Y{&=riǏ�æ��t@l �n���J��$1{�&���+Y2�KPΓS'�'���[�"��NZe�\H��+/�Y>��6J�:V@�W��)vȁ��O�#��.Mv����?E%4�֙�����Z�]>)�*�2[:�1���>u�U4B��b4H��GM�%*-+V$o#�1CQYK�3�q�֮6�w�IX���(�`��^i�d0��V�˩�g��gw����^���S�ɒ�P\\)wR;A�.y���&̚y��4E%�������AM��>�I�8|�~���;1����#���hŌ+�3­ҠA����raR��a�ٰ�>�(1�U�?�Ջ��Z%�2��f���ȯ�!�D�W.���l�w�4%%!��ႊ�E;��̣�U ��v��6l�x>��HL�kJ.�����ĩxD.=��������T��hcF����C�l8���������9	6���������6^6���3��Y������b���xS��Ų
M������-�Ɔf%�a���(ĒWg�Nm~?�Z��"y�kq�q�b���b��=J��ZbY��`+1`Y9���aٟ�� ��C�;���wl�G�{<�ښ�I���*R"��x����y�'��c�[��=5	����l�H9����Q,*���K��v�RA�;�_X����E�s���m�1v���15Y���"�1����j���6��#���%?K��BOLں��qə'�%�Kh`���P��;����C��)xj��RW�����w�J����v��0�=���c��CB�#�k���ى��2%��mŉGMײ7U����o����T���+���q�h؂{g]�[n�G�9��.��*�>}�=���AvaK�V��I�D�����+��Uk����p�gaxu�rv�?JB�k����n4u��M��J���r6$t�ɺ��hTm9N;�@���"�8�X[]���oP�y��(���7i��\�_V�������8�\x��d�}{3%~�s�L���i���^���ǲ�u��AVy\8�?x饅�ik�+��5Wߨy�3ʗ=������W!k����m���=���V7F�oE^P��w?��uj����g_-��'���.9l��ڋ��A��x����{�	h����a���������Ack���O;
�&67�hU�e�|*�+�s	�{{�Z���O̻?`4�Y��yl>n�e����5k7���'������>��w��Ģ>��Ԍ�)gES{� %z�q±G�Ͽt�R�Jz�sN<�;vH,�ζN���+�jVy0�x�-u�~��A�g�$�F#���[��p׬���y��h�"l�ވƦ���au�����5\z�9J��a�c��zp��0k���7]���:�Ia�7�X����0��?����3�p9������_|��ͤ�_#���i�(�Vy�p��X��g���?7j���gz ~_����Ƃ^l~����X�5�B��.����,n���K��sNGFB��t3�9�~�1|^jK������$�$��[���o�J��tJC���6���`xm{Z1��3��ۏ��;1u�%0�޶7&�*T��_xu#�h㛪������S�g�-�&p��W���;[�4�Mau01��g_R�hu\{y����wK1�J���rs̽��oB�Ν��>��с~���ᗕ��`�T8���b ��.��l4o܀W�}�k7蘿�i���T�8*A�j�|��(��g�g�&�(Ƶ7ފ7^X�XG#Ɗ�|������h���;���Tw����΃7�.n��pz�������>�OD��/.|�۷
lEO�N&;���1��7�AMD;�f]w3fϾY��<>�a��A�ь��Mr��ں��SgL�p#�e����x���>@<�ݝ�b�����G�\�,��9�$!J�@o��%N=�L?p(v4�`�ڿ��7������M���������@u�*?�"	�~VK��o9d�=p�!H�mZ[��OI���c���j����!+���o��.���\�R�W��a{�(F֕c�Ƚ������GdcX�2P�^[;Z��q��i���꒍���@U����~��ȉ]/���yt'-q0QW<�o����=ʘ0�1rH��5KQ�ˏ�:��Y����9=l�@)�}y�}����8`�IڞO���.1����
�g�t����00d�0���ǘ��T�;yz���	�C���X�PMղ�Z%�aC����Q2 ���8>���{��*y�!��S�a�l�'w��s �|�#����"��9j�b��o��Kϗ��X�N�岬�j�!��N���^���6�`�-���ï"��ah��?��xS'�7�6����|���0&�٠�J�U����cΣ��+Ѹu+J�*$$.�K�t�R�a��_|���k�\���Q��a�aP���y��K΅���
8-�{�8�1�Iȹ_��j|��2A�A�8�������ڃ�|�3	���x�� �4��T!��JV.���A��Zg^�q�M�f�%|9��+���۲��GD���8'���~����4�CeV���|��E��/֞���P��>mҼ���]����E	��`�O��vZ v]~�%�x뵰��!�ףk,�ĺ���{��۱�Q	�����55n�%��O.DK�@1�rm�R9�T$�������Ü�ga�م���]�{Gސ�'�|��o.FPb(�KR��Ox'��?��\�LMQm��c�+�!��d��Ͼ�^90�$���}V�>KWw?�,Y���8XG�����}L%���h��1#��+o�pI�)�X�l�8��Co��%�v �m݂Q#����-�L^"q%jh��SdL6R���Y��j�`��)��"2Vvl���`�+T�w^\,��R�\언\���gLV��R�������8	��p�"���~����T�v�\X8K�7f,�yB~TYl�L5X.���,(��-M�4�I���l<��7-FO<����FN[�3���(���}�p�1ε+���a��iw�ϵᛟ���Z���d2g�,J�S�&,|W��h�JZ.!��`����5�>�8<�� %��)�9�����\�)q,��[�"��ݱ�E��c1����b,r:��v�5�����.z�[�rf�pU���%���#F3��A�����^�O�yu<>�VnMY0�U��_��y����e%%�x��%���������7�@��Mٳß�x,h�����'�`pgjj��f���vò�+侼��A\)��YI�z��&�2|�=qݍ��.5��x����Jf0羇�w���7���i��Py%^~����R�$�{I��ehmk@kg6nn�e��֯\����b�:���҇K/�3��9�A	��\Hv���Q�\kI�P���Y֞6���o,�M��P�&YC����;#a�?o�?RbF�5b��ۻ0j�D,�m�}�ET,f�9+/޼�0��FZB���?�9`_��FL^��~{�K����?�)���R.�ʋ
�Oo�hR	��mm,����np��q��#Q���AP�,�ϫ��!���O�����V�W�;Z�Ջp��ێ4�����!�\k\uU��H�e�4%/�~[�}�Vlg/�Ȩ��OF��ݏT�Jp���%�2e�Z��Ŵ*bd���T.��`CG��ء	�7>�Q7��}���VOB��\���
A��er`�n���Պ`Я|4z	�J?X8l*���8�FX�+FA�ϴI��5,��9������:�=�YUy�h"�UIX$tx��/t���HBY9p:'$���_P&�?����<6�a�O���m��I;A�Dǋ�/F�D<�@Ҩ�������VGl�=&�ޜ�qqۼU��'�t/;"�(��bf��9"3����g�D��G΢����JK���[��	g.^	`����tIK�� �E@��aqtdu�"�u��B�S�� 9�L�CGoo�a���B�i���ťOFb��ܧߒp���c8���$�S�\5J��� OY�_c��-��5܋��#b�N�#�I��a���{�$*`�>$a��<�<X��O��؇�d?Nr���z��_�$)�Y`�o�خ���<�X�l?'�"rɟy�Uՙ��@e���W�m�B�1���k寷��Z�j��e���4Kj2Hd��R�pg��cMi�:xf��=������f�:����Nj�
lt����e�{��-��PLБ9�S���Bªmmb��Zf$��U�sr����bV�AƦ��nm;GC��������_2Dٍ	��àt?Q&&fY�s�R�y�����d_K��_x��2����ݵ�lt��.�Q�-�;���Ցl��!{KTHJ�������f%�VpX���#Wr����VE�<%E���`?�Sa)�yC9 '�禮�1m\�Z��]Z�B����p���u�8_�d�����<?���(�cףӤ�:R������!J:��O�i�@�c�?�2?w{,F��@	�傒$oֲz���/�G�IJ�S�ư��w���%��ܵVԠ�D���:qrV]?�Hzau�Ԭ!��08i.,�;QI�����I�?Cx>�ʔ��?��$�|.����P�K90�z���	6���R� |��L�g��|a�g��38��7gu��&��VTi�G�|^>+��U-�!����0d�_��ٜY��G,�.���Q1�&>-��L5�D�+Y4��̣�m��g54?��������M*
�-tB��P+sh����Z��ٍ6@�Y�P2#��?�L��3��h�I��V�Y��z�$�H(ِYgf����Y0�"�t���0k��i!ъ�0���x�JCV~yK�Г��C���a��*v�lޱ�tv2���S�2:1,q��1�[i
h$�8�Ұ�R��&K��`*x�,������$G�*5���6o0����EB�ԇw*�y��d^�eU��	����Ry�����:���,\J�ɮ�~���Ԑ�.�2(�Iy;(0j1��IK�95�a��Ϥ\3
	���~a�:�k�|9����w�L׃F�ݖ)�3ՔU�G��������yE|=�z:���P�6�)ѢIk��wM��0�#ǆ:�K9-�	l�-d=�
9�=�-���9C"_�r���PN�DQ*�g�:LI��\�H����ɓh)�	�X_�"E����d 夹ͥZ1V�]m�<����"��h0��u�x����f�6�X
MF�7�pC��T6�����$<��4�"6��k��v���'B%֬��ұ~ne�6Lh%��~�e� �H�n�xR7��<Ӽ4ym���c��Z�`U�-kx|��+h�BD�u��jρŰ�f��i��VPh���H���T&'����jV���8)��n���A�g�fL�[۵ׄ(*k���%�w:W�� ��\��4x5��8lF-	��G�X�l�4�<�.�G/Y$��2�����$-�+���|Nw[��F+�jhUՂB��C���ƐG��ZV�w"0y!�u�|R�_��h�f�Ԛ��]f��NX2�����p��
����j`�q���?W2���ԩ�P��:�l zG�o�56`�Q�N`>@>7BBi@�w	���ax�p
�7�Yʑ�!����y����h�!�$X�p��pƥ�ϵY����yinj�qGO�>�:(xeb�j��v�*2�p��|��9YK��ӌ����%lv�]������|���)�g^ٴx��g�z�/��f��Y[��N���U�I\~�PS7Jsiԅ!��I-�ܧ����;��sQZYslIA=����=��5l��	kk�B%���t���'�E�C��]�__��O��?�*�)��5KnB�74��*�q����x0��S��dr���8��1c���.��X{G�@�VJvK,���fdG��ŨuIE3ټL2�����*���\VV���/�@Ye�6��C� �l.��������u�,t�ZyF6�쐐c��5�I���h���w,!1�ǎ��f�3e"��AGK�\��lRD�q���GJ˴\���
G�㤼���b��d-Z5�dh�?GS{V�\��ٽ�#�lz��� |r(w�؆�o�%��|��]m�D����oCfYlk�[�ДͲ'Ņ�a�W���;w6��r��{ �w��<���dd�Y)�.eZ�\�r�`N�1zT�̘���zF���s����=�#F�Q�Ng�9�:e�#��x�I�}��w�H�\�n9��0n�5>�zQߔ<�jظ��3��C��ϡ��Q�h����S\�%+~ŗKW�ޔ� GLN3�aY?g��|����g])(6�r	�I��&D�*E.��:T����X����ɟ�&?��C�˻ĵ����,�V3t(N:�<p�t�~�!��1��d;y$�կ�.;�]��^���I�8e�d��$�p�=(��U�P�M滈m���ۚ0�����"�a#93{����.�٧�����(*�T���0�N����&<���rV�`�#�~xq l"k�3q�g�'�z���(��KZRR&Vދ�;��ׅ����r���v���|Ig;���?9`/��ø�^��9-��K��y����R�)됑�3rh-���f�� ���i�V�Ho.�[�J��݄�V#�!Cz"��\��]���X6��Ҧ'�F�ǵx��e����'�;S���;���#���E�(EI϶ܲ�2�����;��e�F�2��gί0��%|��b�ȡ
;�Z;t���
�p�Y���wއ3P*d�x>_��`�IE.?�2�ww"&����D�ihv�0]�����<��@�4l4:��xt�l��������*Ɣ�dW\|�~�������@U:��Ұ�_����b�6�T����ɶ��q̑���O�D"oHE������lV�����=�5^yR(���f�q/�1̽�6<����UR&E�dcS�1�"�SO;۶��!���D�7�Cr�~~J.�7��7��ɦP��-�\ZC��`J��jl޴Q�3�Vl� �6fY�#>DyX���vA>Tzc���h��6�<k���8�f��X�ȭ���ŧ��+�A��/I�x/��f�|IL�u�����]��p	fJ�XG3��<������CZ��v�I�bHu�Ο�}�N�(	R^.$����{��s�D1u�Lq1�8���q�g�Z��k��Ce]j4h(+��wx��Gpͬ;d�]ꂙ>�,U{S3{�A�|���+�E8�	���{�/A{[f�]����S"�jN���U�GKB�{�9x�ŗT4w���.���т�.8CJ�1���aq;z�����w��f��/�G�褟M0�&�c�D����բ?�����F��T!��3N��o}$0�L���@gKY�tng��olZ�B,k��r��i�:���a��I8~�x����h��P5�P9ttt����B��m���:Z�NK�N����.AU�e8q�,��3�R�Q�_ʋ�X����ƎX��55��aayk�C���v��gb�_����ɚ���^�LO�g�|"��$Q�6T���q[S[������#����M[ŕ(Bbʢ9��/@wg���>�_�E^?��1$1�=�;�R��Wu�?_�H���jo�i'�k���UgeGCL;���"�WQ����O��]}zؙd�0��Չ�=
�GסG>k��:�=��^����&\k� tt����������j=��֝�'���sϖ0��#G*7�k֩�_(�5���e'n��*�{�eE�lv�	g(���7\/��@������AF�4�U��6HF<�>�M@�ć�|GqH��\Ɇ���LB&qer>���w#:qD���|�@u1��=>7̾6�s���0�����Um�ΦK������cFV�أCV�D_�ه������k@�y��=8yƱ�>�V M�xl�s�߼6	u�N��.<I�q>�\s��[�N�Ilv�^v��o�$-���U�[�`KC3��=x_\{���v�I����9�]���a��;�:q�m��/�Y�o�����XG2��*��7]�ɻW" +�ʬ��H ��&#����<�~�v�Yx��Wa8#� �f�}��P�b�J��Z|��
l��O���c&�Ŵp�:v�� �V���b�)cq��dN^�(�߯��u�dS�H��/�Csg�|�t���'(�*�Ϊ��D_#���${Q�/�?����_�!�1�8�����b��9������
)�YN�d�8�$x���������g�"[�?��.9��[G$�quA�}�Qrؖ�%�+�f��������b�\hq�����>�H;�8��������pƌC��'K�z�,1>>�'v��L�x�*�M¿Ͼ{J٭	����9�5?d�X�$�X�~����C'bݸ��3���P6l�d!�nhQz:�1�_��K/��P�%���1��74>�����Y'��/6���ٌWn^��]m�J�1���d��L��q���e�r{��Q�$=x�	[Y�3%������_��4$K���F����:��P:p�����W��.�(K
ל���1r�i��懱��sV��k*���mW�Ebz��}�L�t��p�Vk<��u�3e=�T�������T����!k��=7Z��ƾr�v��X�i�B�L�w]s��\��o�o~���K��y���+9��u�b4(�x�7��G�AD��+�q�>�P�N��*�wk��������}�l%��f�=xl		�u�p�E����p�Th�����1�!F3"N%��ϻTP�S�̙k\�z;���a���S:�0iT�V/D}Iq�ќ�q]pU���']��bΌD%zZ��z,Yr	>xc!��6q�8����+a�����C��x���mx���P�|C99�x�a�{��$r�ي���ψ��hB���w�&��.h�hjǡ��o�)��X��`��`���(.��N��I�^|/�l�d��=�I��(���:�Ν/^��В�p�	ǣ�~3\�b�~��Y���i��a�Xٿp�9g�8�B�ˋ1#��%�҄(��Gq��
:�~���X��.AK�>�l�������nT�0{�g�~:^y�#8�Nm��Jz��������+�Y9a����^�0m<�>l���
	�|rY5�/��*\>����$��ށP�<���f��>��=v�؄�R�M�8�ަ%.f�GM���}Ḏ�~��(+/��de��2�9s^��^�݂}���𫠁*m�N�Ώ0��o��&(��h���!���k���k1�߃�c&h��ɨ2��a����câ��E� $$r���_�G���gϒuϣ��O9X��ui^����n�!Y!��{1��v4�>3�T\Q�F���<���Y14L"'�9�!��1l������|�5�QY>�p��GJZ�p�}�qǭ׉Gk%�m�=��g���)�$�Kj��gK�qc��w!MR��z�pߜ�x~�\�Damm���ذ���v�﫮�Wrk����(%$i	��c<��e�T��94���G�iUU��Y��@Y�{#j��+145������ࣸ��a/h(���-�;�VV���Kq�C�(�5�ȹ�)Y+��1���L�2v�A�����K�cp9��9���b��J4tMg"��6�?��Cj����,A�v9�+׮�'jPF}�UΠ_~�(�xL����tؕJ:���6����ا�@�Dg�^�u�C0wέ0�u��-� ���!־��\6�y�w?_����R�v�yh�l&�~�)<��,�,�7ճ�|�H�;���G��N	_B������3�j�a��zL7�Xc�Aw}�f�?���/�+mv	lo@��Q�S��S��j�����-ln"�.ɉ�r�)�p:�)�6_�^qy���fa�U�+Vm�1G/�ա�TD>L>iÛ��A�_��k�/FqeH͹Ll�f��_\�O��ZP�m�)d��z��p.bW�ɺ�[Q>b�A� ���.���Ðe|�sO9mr٢nR�aC,'���Kk�٪e��.J�����~q��[�Ϙ(T��Q�[ s�c�,���T�<��N�$��Ub�o+����Āˡ��F-������~���'a�+��`uA�,�:�Ki�>�r���HK�L`Sr��VJִL��ʵ c��D���z쾠�{�xo������8�j��������O���pk����>ٟ�8��b���+�߿vSfq+ݙ dW*9_��߁�>�H�Q�V�XfL��c�aGK��Sv���=Z=2g��v�fı��j�L��H�%4���'kf���3D9Sʁ�����)�e�5jdEI	�ύ��~�$��4s=���������GCt\Y���a��|�¼��K�_���;iU�yKԩ7��������'�\���S��Ĭ�F���e��T�!=��Z*qA(���1,/��!:��z���S��w>���'܁e�&�`V�}�A #G�����-�E��� �҈�X!1��o�I�`�x3^TZiN+�"�r���w��������c:s˲�
�l�ֈ��x���Lֻ���n3���ۥ�3���K<�Y�:� ��C]	Wy�!��v9 ~�Y��ȍU���)oGJG9��9r�oo�A;YVZT�ٮ,��xR�����3�'X.��,��/�ӯ������I��(��s��b,
9��f�	�a?w%��em,�!&�J�2�˪��#�w�R��/�Qѡ����*�'��R{<،SVV�ܫ��A�C��ɋ�d#	{lJlU�'��X�a��*R}�D5y�r9��|���X�3�#����e�\v�Q��1@�ONnJ��4gt�"�)��%�>6���-�\���1���`��a��¼C/J͙1��9��5f^��V1�2��%�&c���D��P��4w�K6@;J-Z��ی�zI��n	����Uv�+�IU�`�MmF���K�!A��l��ay�J�'?K�Hq���/��T"��
oTؓ������%�
�N�]:]�J�ar˟���U���\���Y��ڦ�`¤ �ᾰv�z$6u�~fRV�3������Z.��t&GE<,�x	c*��>!��odyYS�s�f,�������ȣeFV�9�CgJ�yd)3(��_��B�^��d*�HH�Ͱ+R`�\R9�l�ul��ܠ\�.a�߳&�NR%FM��ď.	p<A9D�N��T��e9�/!��uP7�"BL�r#�-=�9bq��8�l����	�6� �5�e���t�F�z�z� ���]Jn��@Q�lu��Tv:���?i�?Y\nV��Gދ�L���Jo1g�&�;F{]X�e��hn32�6����R���%�"���<Z��咞���<�?ͦB�IV��(�h%�A	�(/
�_b�[����R0��u���%e�k�1z1�U��g�ܟ�7۽���z���}r>F���Լ(���WBw�#�6�^dU�xxj�X,M���Xŉ�"}(�Я��E�k�9,��RE� Q�.p�N�|���
W�	�9��,�Ҥ_�+P�~�9y.�K��Alo��/+��"!�����Ce������2g�*PZ�nKs��I���?V�H�W��I�I��`?FV����e�y|Q.��$�r��z0b�,X�ŵ:B�pV�X}p�Pb�n���]Xn�0YĬbp�_��/~Z�}�p�g�<b(P��8x����=#�ř���*�gK���Q���O� ���up��:m�ډ�O=Yũ\N�Z��p��!�bu��5ᤓg`�c�P��5k�/!}t0����&vG�E�I@$���4��٨4vᙔ%�\��9H����cGT�*S��X�~������j8L���<�^��j$���d5���E��I�k���*T������&U�f��Q���R	l�
�Į�T���ތ�����h>k^B�Tܪb�t3�_�p���lS��?V��G��*P�t�vx�N9���2t���'���s�������żp���,� �F�8h�$�5x�����cϊ!�������i�Dل��w��dCG���<���)�q�VT�ӵ>�K�w4= F��Ue��Т���R;/Mv��b��y�ޓ��oI�G���:��	�B����NF�+��ҁ.
	���!��_t�-|E�f�!R�23�T	"#��:��0�!�+��+ψ!ij؊�O<��ހ��	A���J|E(�
��j���o@˕l�2t~���Hc�ɣ�js� 7��y��2�F۪ә��u���ݷ��DVR%�wn�Y'���xG{�r>�2�ňt�ʟ	h�rL�~0�T�ərZ��%\K(^�1C�$��c�\������S�y��7�h:�j�e������c��y���4,��[UG��O�d��^w��IXΜ8H1�&e��kJ�W��#�0!�x���`���P�{��%b9��p�3PY^�ܼ��;TNT���,�Ry햶˹-������&1
	q�daoߺI��$�溷��?V	��D��%(��ǟ��3/��ѵx聛p�-����D�s��cO#!��kk�����P���|(�K�X�����m�&�Щ*ElJ����I�s�rN����Q\�3'z?��`Noo�΢�D$%�&��ˍ#��Q���?)0���m(oT-F�J�=ꠊ��	G$����ӰSQ���Ǎ�x{�<�>�j�Z�'rP6w.�0CH�]���A�<<|VA��4���	�b�xK��t���NC�O�C��/F��,<���d?��k��$6{M����I��hx,���Ǡ��M�+a9@4t��0�Ac���7��=v���9���/�߰E.lL�k9۳Ǟ�P[�Nq��-�q�H')�ǩ�Tʴ&�F��#�_U��t��3��?���x�HKM�W���nb�+�@���L?R)�N�q���'a�>��!��3�J��t�o�A)�O0��-[�N:�P�F�DskH�S^�B{K��Rv��j0�3>��k���x@��6mބ�&�E���M*^3�_Vo4:~�P�6��M����ۻ|�re��sxL;z�x졹8����0[q�a媭���p�J���#�<�SW��z,�u���DȤUS�;��Ξ��֝��3�f�m�c3^M�'��܍�Q	;�A�y��Z�e�����`��5�kʵA�ܓ�į+V�G�N�8�����@�8����h9�d̹/6��v�}xt�� ���+/DgS3�w��΁��Z�$̈�cP�̋��.��Gښe�َp�%�b��~Ep�IǊ�b�ʵȈ�:�kѼ�A�y<����eJ¢��9�[����q�'��u���c۩����bQE��ׯ���}w�Ͽ�&qu���:d���1�ц��G���W�V2��%���],��oL40���|ƚ�����#0�
3���b����'�w>�\�[�4H��q���p��'*��:k7l@�X�Z���k*P�K���x�o��	��Y�^�j���}��S��-/B� ��;4>a��Q,b[C=��~_���X�4t�6d��3�����8`�h8=6��A�`�:�DS�
�8y���[XCU��9q1ci��-[�c��ۆ���Q�ֶf1��\�Z���,��{�~��/���9�(~GG?��g�r,zv" ���C��d//:��ڻeÜ�a��ݺS���Cp���/�s�������N�x.\s��J�F���׏���,-E{g?��q�x�PavA.��-;[���C�K=��s��sUA��0bu���ܲ.P��M�z��� ^��s�4�d{����8��:�tw���(&)�Z�ʯ�[�v���k�d�9��J<��G����ݲ�'M�a∘(T�Ge���G�8��l�3�Q�dսt�-h��~��bh(�9qo	%�m��,$%!�rAA�?�ه���K[��T���G��O<���[0����w�VSb��E=�,�B�y�xJ��X��e�X%|���U8h���l�(��o��P4e�0�=�����Ș��9�'��p!e��9O㦙�}�_�B�s����T��8/���{�l�a��d�e�v�����9x����3���<m�:�M�*m$I���!1�AP��9����%��"ω�N��nA'~�j������?���?�����N<V<M�R��۱e��5�1�?� %��[�3$�Bİe�m�9lځb(����ŋ����B�KӬ�_����͠1�1�������Eo⸣�PR� V�ݜLr���n8>��k�sz��_�0%I����7b��k�l�Pj�����ukQ!��)����K�`��~9�v�}�Y
��VnX�	vC�j�^z�a����S���rǝ(����!�l4U1���7�(RaՉ�>V�C���Z�60 ���o�v"��B�1��-���$�X����o�`�5 ��+ތIƾ� bAzk��(-)Չ[�38��#��˯��sNW���5��0��e��ra��������ߘ��\M�G��j5�r9���lk���Y��v��xB!<:�ie�%[�-yMvT��x��q�駠��Ҝ�u�`�qc��V5�ϿlHn�����	y�7)��~�]�~��شm�" �����I!J#2���%�}ʱY�7��11�-��e+p�qG���O'���A<�p�������?�g�j[:s���
�o��&�s�M���~d����̘�ufq�]sP\;\�殌�����/��òe�^)�p�	I��r�\�#�����`���J�&u��oB¡�,xw�r��E	�p�v��_6�*�5Q�3�o`L�2<d��/�9��ٸ����^S�(!#��YB�y��X�b�!ё�)�����;��K��7?�ۈf���A�$D�&Vc��_tP�J��ޮT�~BG�V噰�a|H�o�ȑ:��̰�` �ˍ��w(YJ�jZ�Ƥ:%�-��+o.�k��}���@D�yz�8{\^|�շ����t^����gjk��/��#I-�1�e��'x� ҊU�U6�*�	[j��0��'1�o��)a�O�OL�ڝ,�%�}�}�݃1�U_��C��JYQY���Mk1R&ռ�:_�&���ȪI�w��,XZ��>�G~(L�11��>Z���xK��CuX�lhw�1��|>c�z��yω���k��I�i2lG[�v�pW<�Kj��t"�.^(�}��1�0�fx)�ty�"==x��O�-*Q��):�]�Ո��	l�s�x$;j����w�$b��o��L��兴��F��lL/+
\_^��>��y$6�o�x8��E�)3�y�-�tn%���kN�L�@V��&����K���hC��O<-x;�zz�~k|�=��f"��\K:�>ge/6�h��/��c���ϣm�6�C0�e�N��B�'8UtK<5��$6f{>�
�>�8j��8���a��p��@%�FH����I;r��u:�[H�.��ذ}�B��G�)s
�qG3��`Ę����(̍� FM3萐�<,\1Ks`Ѱ�Q'6�ȡ��F�8t���&�hP��	e&��'y��Ex�g$�j6[��� drƐ$���=c
�q/y�=�bt��0�����,��C{N�|���g*ݥ��&H����ەC�H�8v���(�2�^'��X���W��Vs�/C^�O����U/@��~��{�."Γ���8�?�4lC�9I��P	��l��㑸�m���e6����{��_�\��+~/Lf�2�gt$�H��قX���8��7��i�=�I���Nmɲ������\0��[T##{4���Ҧ��*us��]T�%?�*4^%�fl�j�9�KOb��+���pc^��mr!�{�(^�U�T:��<�dۢ�gٛ��g-LCU��%wxC�h��X�����pr����|����9vMW�]ʙAvlA�Wo��A�ڂ|��閃���$��T*%�Ʌr�j�}*9񮄢���3ې�i�6�9��#$c)7���f���)1�d+����[��Ԯ�0�B�/Ɩ�qNs��U��{4��X�Ó���H.�Y66���v���M'jM:ʟQ6��=I��p�+�G�k�����u��}n+�je=hdȖ�^��8>)��:�ъRo�_.qN����Hs�^BV�l6�?hc�f���&�y���h�ѿN0�lNm�$M���N��g���ȯQ�=$�C�Cg��,pl��!�k�[,�Z���z���ȳaQ��3��������e���۩�!��Y\���x�{!_ �Q^q�U�<��]�yJ䌵�h8��yع�(��6&���{�W:�m�+z镸1!�#�W�$fz-ʹ���#�%C�J�ʎ;~��dm������o� ������#�$R�u�ZS�rC9-x���$�$C�]<0l(�p,���1DA���v��9^墀&7uwL�M�~���(��;t8�C��PG��^�ٚطQ8dZ_�$������A~��$��F47��IE�v�Kwq�����Ť�cπ�d�z��%Ƽ��a�qy�x�P�nL�>D/-��\Z ���F�utb,�]�=��/4#�	��j+f9G bׯ������+j*E!�|N�ML��g�ȕ�r�ԛZ4E�̦$�xHh��Yo�ʕ����F����19��G�~��t����D���J��\��}M� ����QA�n�MPv�g͜�?˳�`U/m��X���.`��1���w۴g��a���JU���U9휶�ty}��ֳM�0�39t,�A�����(�Y�kڐڵy��[��qSS\^�>�hXu�篪��ĳU/a�@�@ߴ፬ּ���$�dS&��Ŭ�F��s�!��Qi�])08-�]��}w�����3;��l��]����?{� �&�����%�-�7���c����  ���;�;;��wf~�9ﬂ��u��gX����~��<�|�y�����ʬεa�F����V9͡a~mR#a�ǒ�4Q�䐵V���I!PZ��T�Ԁq�e���<Y�@�b\��K����Ez�cIk����АM�8�����'c��w����_��F��%���Z�Eڞ�h���`����N���rj��/,sH4�WteҚ���-�c�!��1�D�WԨ�5�e��$��J	��ߣ�!�!�6��� �UQHiS�1�b�iP�FBC�!���7˨A
CPɫ��Q�����[����অ.2�����9� R��J��F���H�W��GA��Ԕ��J"X��
)���5C#ٱg�"*q��煲S�ȰK�u���r%]���"՘B�����hE(SN\1d���V�J�85����
1�x�!��'�|��Q^Z�H0��9��ke����ވ2J��8�ln��\���>~��Z��I���)���c�wk0��!݅��/��h�
%�����^4�3�!ˀ�4	_�a�_^��摊�$ǖJ'~ȫ�b��6,~�I�Jk�{9JK�d*e�YW1�)�&���-2�<�1�P�:-~/VIY�L����U�Q-��Rd��u:;�X�2KE�p/����b
R���	�,2�����..�-/�D��Z�e�9��"�d0V侃��Ҋmo�6YM
	-Ũ���x�d��g/!u(itt�j<h���*K�4�Z;��VU*�0*�A5�aƐ�4PH\�{�j|\Rl)hO���2%{�0r�9#�8/� ÷����:�0 c�i�To�R����4������C�9���.�������_���J-pz������.�Ȕ�3�9# fE3���ؠ3v�ePo..D:!��Ù����z��&�� dԈFL3F���b��O�}�[v���ة�g�%�����9T�������:^�$�iWk+�����k�]��Cf�dp �4C����~���j�B�S��4������IftO�i>�pJH>�]m����0����u0�)r��`����/��zX��J=���ҹ-���zѹg��ѕ����g="_0�j̞y#�%Q��`�thug�1c�4L�|R� �>��
�,f^r�}�%,��;x��9�?�w�B]䇴�������2d��1��#ڼ��ޅ��|W^v��Ŕ/��r�K�|�oѢG	�kq�8�t�N͝����_¬�.����rL�0^������9��6��۴�,�]ӄ|�H2Z�/FF�����N��<
��1G�̜����[ SX��٭�̜�82J�$Yx���pΟ~&ꪴl?��܏`8��>��[{��ߜK@*�]�:
Mq���_|>C�A�+���խ�βQq�>�|%��!IF>@`_V ��{�q��	��*ҊQ�ruPS��c�%�W�=GX�Y�B�Pq�	�.9���\x��ڀ�/)E"BII	�3��֗���K�i@����tK�٪)�ݍ+ϟ�ۡ��wsKqP0��/�O�	!����욯�XS`h���c��Q��=ϡ��ߋ'��үVj���;JӡP�I���\R���a��(�Ϗ��4�W�\^�1�t��z<��ex��,4���eh��"�됟��%睭��k�+	M*��{�1��c�|�|��&��E�٬FQxO����W\v�;�"���ڴ8��Y�G���m�܏��J��I� M�u���b��M�oW�$�����5C��=�H�Ge�_��`I�Ra��}j��">m�����!_�)�Ϳ	���Jkky�f�Va����@��z"�j�C��V}�x:�V�S����x��;���'�E��t�� M�EN.�z
?�����Oq��`H�{��'�_R���_����P��̝��㞛.G��r��hAؓn�cAԕ�;�ă���[�fD�H�%
�2���m�sO�^�̥c�#
�AXK�ŉڑ��Ɵ�|7,SϚ�8�|P˪�Z�,�B��X|^,_��^ç�u�K�E��p��t��ůn��{<@��c��=:Y^��(�M7\����=J��?��e�)�T�X�ι�@cƸZ[������v�#����k7mך ��ƨHa�J�Hī.�H��B�8�f �ݽp�h�Hǽ۷㲙3��ko��J)��2v�VQ��|�!(-)�i�YGC��5D��V�s�9\�"�����Tg1_��\ c�i�&s�%+)C�S��ĈL��<�|کx��%((�2l��C��D"Ҍ�������=5j��܎�ؠf�M>���m�<�lLj��X.���O=���f*Z��]H#Y��0��-j�.<gz�	���%ڷ!���_f��Q�Ŵs��@����AE]�Ӭ#	C��(Z�������7��|�lV�54J2�4g1c��u:��+%Ӆذej�ׁ0>��'�e����@��������.��;֡�����غk/�'Ch^�V^COh�3w��w��s|�yJ�ػw��:-:���i�R��s�:��L�߻�݈yw��^։��5I���}���S�(������7�x=�4��8v�1�Qƣ�<x׭X��#pWV��r���ݸx��p��њwȳ���?�{�����}�5W`�(�����n,�}���I�[�:�:0��+P)�|���z�z|�d)eَY�OC�^e�.(؛��_���!���Zq�ݷ��ā�͋�n��r"�Nj��s:.�l�6���z��.,X�[��|���ֺ�>�g�uE-�\p7��v�NS
��ê�̢�1��E�������ب��ɬ.����.�l�Qk���HI�c�)��x{`!fZ;[���عa���å��#�֊��/����R��A ���u7���Rt��VA�ISݽ�4\6Z;�*�$��ʰ}�V�"Ŀ
J�)D�zp��b��8��hv�Z�}�X��ࠗp9���?u2�{�5��ZiP�NG����5�U�R�\�+�Y���bL�r*,D#���ꗳ��ҥ���|��^�8���.E�����K�����_ժ��&M����ظ~5�63.��T����0]��{�}\z��ыĬ@�}����S�P]Y��x�7��!�;��_x
J��g�K$��ig)����;0n≘7�N��n/�P_W��7߀��6bDM=�����w��)9��؎c'�S��گ^�Ͽ�;H��_d��;�q2�)�����=�� �D$�"7׀��������X���x�_�V��QU���__�A�哏�5�7oS�[�Ō�}�q㕳�����������n�v�DR��xuѓX��k�]���v̙w;ʪj5� J{t᭚`�8��g�b��@ "���<�@W�3�����PV���ɦ��L:b�*���]�-(�,��E���x����=���(
�.#�Z��2W�LƎ�ĸQ�Tv��9��%����̙^���ᕋ�ڊ��^����u#PL]�T���U:��hx3fθ�����I��_?��y���/����d6?�� ���9�`%z��_+�ȟ^ցH��(O�;�|�.�s��	Dc~�

4�9�.�β-�o��>��[��ZuƬ���u���s��T�wA9�z�O����[�8�6�$��k�@���2�dD.e�����&g��w���{]��T���B�w�YQ[LC���s�╿�3Y��e�{���q!K�}w;�x|>���˼�K/�'=�$�.�}>�x��J�XW��~�����7�7��Q�Gy(�Y��-�;��&lY�5Úhm��/Wj�Jx�4PG�q"RѠN���{���ta��V|���}�T�=t$��<��Ǔ�t��^�=b��WRH�n�N<���r3�D�^|����ϚF��COg���ֶN�T���aTvSr ���E�2̸d.�>�Z6����o���.�-�7b��s0��ߣ��Fs@r��X]���'LY��UT_u�΂�dx4�{�`Ε�����JJ��赒DI���5��\����߬^{��C��������p��E��ru�q����5�f4QYUFTB�X\x�������Z�.R�8��'�����vt`,�u3�F��c:�"�n��r#���ү����Ұ
5�G���H�^y=�~�n�vt����J��%���^�N�(�?�y5�|�p�J�������5�z�n��<�oŔ3Nǲ�(�AW[;θ�BD�w�����P�X�!��f��K_,����G��t�z�1rx��)1���c��:�X	8�N�<�ȵR��$�#	K��1�B<��B��h�	H!V��0�C�:m�$��λÐ��]�"��8J�kpٕ����_F*�K,�b�ϐ#IMœ�`��l��Χp����!;����1���e��N��haW��M�,a��c���i"��Q�����zڦ�f��������7�QTc�_~��e�h&EMv3n<v��7�����i���T��hւO�\�HB��C�^[����7�B�=�C3������o~>܅eX�؃���(�w{��ϼ�*��d�Nϖx�z��ު��~:��cPZX/�?_e�N�$"�g�p����'�#����B�����8�DUV��o��7x�D rl�,�VX=��`�2�5�`��FlܶM��")��cȽTV��?ԇ������&��9�s���+�o�n��M�ZgQZR�����0�72]����,U~�X�"a��\xb�sx`�uHh+'Q�/jbIo@l����j��&Ɍ�XE�9�z?^��N>Q:���"m���ak��3g�Qza7���
����F��	9�"���Gc��3����u���v�l��2*��k4����8�lل
��d�����&�gh�|�VȜ�cS�ո}%x�W���{��M�^��^�������b))�
D�z,��/!��ϼ���j%e�H;�$�]��/p����_t����������yl�qA�e_�)|��4�o�#Lh�%r&�d�����FB���ە��NI�A)>Pn�>�5�q�����t"]J[��@�z��M��42Ke��.!Ҍ��,?�)�4�ĳ����m���MdLϥ���rh���BZ
.-�ťVĢ}���������2�����Ñ%QB������D�{�
�+�B��y�		�S�C^;zc2F���E��	���W�}�2�aɲ8d�t$��1\��$�H�.ZfiW߲v+��k�&�xGj*��G�-��<��F�$�L��)񬿬{�`<~.�~8ڣ1���m�|��v��q����fS�d�� 9�к)�IB(YL�󗤭)mAk 3�G��z��f0�$4z��En
�A[W|�rD�0fe,���JԜ���;��P���dF_�,�D���tz�FDe�5��<	ޏ���+�⨱MjH�yܔ��5&o���Z���MZ�rXt�xذX�a+jJ���5w8�z�&�RR.\�w;�����D��/0�H,:2��)3,��Xj" ���:X'N�(]�k�m@	�2�gWB���Xt̾�n�ne��I����Y�Z�����a蓹CI;n�A��o9�K{GJ�e�q�a��0�΋i����.�Z�/�g(+�!���O�~_G���ZL��ƌR9����f��:=�a<�?3i�JȜ%����R�1DJo(C�dv�Ms��}��hUg���F:�uMi���ϋ��!\�=��J��g�$]���wӓ����ý4��2��Ak
|:--�i��%Ǻ�J�;i�ǩ!��i�h,q�t�*�
qut��Ce�@�b�����Pݳ9�t։�J.����	��p��6즞�)��9��N��ʘP>�Ǚ�0�%�]�R�p	�E��X��rqa�*�A�/�C+^U_��K���ԫ �i�21JN"*�����g��Th
�����$�l�b#Q�&o�Qh��j��L8�y]�*�v�&��8����9��ɇ�fXz;��%&��$���}Kܴ��N%[�dyQ�~~tP�T�(utn9y�~�T�(�UN.!�0?ː#�Nt̩�
��\)^���KQ�a��)�
8K*��wk7��'�.^6͉�ɩ�6e~�*�0!��ϘrC��^��l�A+)�gi�̰E���8�L���6��XD��\Z
?�����{��	���WT�!2�䰙�m�"��4��n��š�sF��w��X;ﯤ��I�#�TQ���"�H�����=��m3����Bb��n�5�d����K����� =m�_K
}p��.�Q%��&:�H�G����R/!�������,	��=������tʐh:Q�+�(�p]m��ԡ��[��Pɽ���9ڗ�ݼ$N;�d=Ζ�<��.^{JɆ���{2��i=��L��%Jm�*�t�#�1J) �O9$��OA�R�1���/"��B������m����c�Z�P���aѰ=�Q&�ؾk7u%��`�H�}����u��v	�;v`D����`.,�u�:*��H��:����c�b�::_�E����;�PuR�n�:}��˄=i��dS:'��'`��/@�0��"�r~Vn,)W�I���H��x^8i�o�@Ǟx(`m}$�9n�l�a�Ç�� ��걫�G�OQ��?�{,��{	����Sk��=-FZ�lB�����c_�ι�S

�z�Dj����ݣs@�Zw!e1���V��Q��A�.�î��m14yi��(�Xa�
y��7��ʘ��V^i�T>���0c�ʒ*�Ǩ,�qH��`5����Dz~T)���&�h ��]���c����{{�0��`��f�̽3��u~��� ��%��1�)�X�M�6I�d�a>apr�P�=F�ZZ������ܨ����l"�)aWOn�qh3S ]�1�6�V�Y�-*/�#G6�����>x��*%��0Q"*�����[o��,Ё�y�|:�8�b��.Rta��b�=�Qp$!�NW駡0��ދc���-��~�"t�|;<�ǥ����K/":��c���B���c��:lf��V:A����=d4ٛ��|��� ��E�i.&4��8�:��ڎ8�?*�P��P�<В�Tr�����|�)�qa��ߏ(u�"��U��PB�"B�J`ֹS�\��� I���,Y)է�^�z3&�q<�Zp�����?U�k�UN ؉�s�E��-p�k�_�1�N�D�:x��E`�V,�n~��?��K�چ�"98����S�(:ϗ���ڔ�F¶,�Gu�m�F��r�M3p�ܵS�X2�0Snlyq�~�mJ���"|��F���X�٤�.�Ś���0"���B]��w_��Jmaxr�ԟ�	�h�|��e����Mʏ�6�J"e�`���+�����b��ס��M��V�h���"�~"�*\Z��=����&���-�6�j���_y6�8K�XW��C8(�#ޛ�p"�G������@��O�g����ϸ���Ҙ�A���W�T�V��J5]0�<Ҍ��أ�aU����0���UAD�j$Ċ9��I�U4~�]pñ/QT_�ػ�'��I��5?m%T����"�6:���_$�`�8
�ؕ�A�J"�^
j��D���q�'Ӫ�U��j�2�׹�+h�c{�D1�Qr�x|��s��M�k{�N#�>��"��Fq��OB��M<h�;�L�hL��q�-jc��N	��b_E=b6*WA���.��G��?�i\�ۑ�����e���^���t�D��9
��~V?�݋@�=����'}D�u����sеjR�-���a�i�Ɨf?b�Bl�ъP�I����S*t}�x|��ۨ){e�VE��G���E2�Fsiģ%�=}l�4�ĐE牸B��ǡ��B/
O�c%�[LȜ�����ga-��ְ1��s�V�:l����|<�����2lh��Is���|��5�BX�#�ш5v�0�!WY#�m1R\�	�jܭ�pO�2��?�1�h�!:�2i�������b���M�C�v�jN��e�4�M|N�� >�h	C�rD�&�Q��Q�N�[��g07�����K�Tq���M�:�j|�9��n{=]��S�8�V�/載W�um�|����:|K
2��Y��?+0���R&3#���y*bDVB..�o_J�ua�{Kay����S��E�~�����>���#�xsߔ��[�� ��8���K~���=��i4�������kT
"�=r?h��wo��������K.�7���M>�������8y�ׇ'��?��O���	���K_0J6�����GH�jvҙ0��������u���g��.���G6jP5��iT�p�����k_�$�<��{ܿ��/�~D�I��g��Ds_r������0��_�g?����곡k'�@i��Ce%�{�����7�l���I��o�+����SO���[���ԟl��}N �s�z��{��C�=�3����$Ŷ}��<��4$���?��~ߑ�*r'�4��{_������m�:t@ׅ<*F��3-�ǯ�܆�qK�$����}M��B��B�z0r�r�7���z��`�f�)�A� =dͥW@�JA��|j�u�5��jY����O9��5?��ϐ5�	����������pXe����!�(k.�<�v�:��jW�u9��f�)((0�����E�Ņ�6H�    IEND�B`�PK
     �8�Z��I2\k  \k  /   images/35c60fd9-1fb3-48b8-b3d7-7968b0279531.png�PNG

   IHDR   d   ^   ���   gAMA  ���a   	pHYs  �  ��o�d  j�IDATx�4�gt��q%x�!a�{ｭB(o���ڳ�dS�(q82�Jgݏ=3s��3���h�E3�'ۻ�e���{�H`nz�S,0����ｈ�F�{e��pd1��ｃ��v�y���?��L����h����@rL~��ط7��ߺ���5�..�t~&�郯0����_�#��60�k%���N9Ʀp��)�z8��}�^(�O?��%~���g����x�r�僻�\���Y�KK�'O*����yـ��~d���օ|��^?W��W�{p�)qx��9��r\>}����֍��0|��e��v9JrR0����O�!��?��������_^��z��`O�/�{�7����n�ɇ��l=�_�m�L�ceu	�K����8ğ�{&��Z:p���w��[��n������g�x��y�����5�v�y�����?�=��|���"'&f��'\�̀�vl��#���������;p��� }���	�����#3˰�wNVgxy��a������q ����
]���'g�a2���{��zW~~�8�?&�	�1a��t �ח�>�����?� X�Vi0�����?��3B�C14����0lno����l#+=k���M�ᔙ����GxX <||'�;�XZZA���H_�\\y�,�,#1!ɉ)�y9! ��]��ݱ�l�
���GG�����[�0L8q� Ss3��IGKs����l���+�04>�����s<;��uo�zU�C8��w�y^V'�� �ַ��iUF#0�����e�������W`q�`av
�c�pp�ں���k�e�þ�E�h�"�x��YL--����M���Է��3Nc�~ 7�O��`�;��%E8[����<�i��l�W����|�g���ǳ�F�Ǆ��V�++Ɖ�T9��U5p9�yΝ��޸���Fym�.ncw.��o��6fO*����@k�0�=<�o���X��6̭�������7^-�'���cs�M�Ђ���\Ԯ�4u���g<,��e�`uK�'������~��7/�$3#�#x��Fl���wo^���ct|
�N�!guqcC-�Gxʇyy��W��o�x^���(�ӄ%��ȤV�24���E~n���6��,Z��(��a�8���G����JϚ���ܜ������},3f�������ױE˲X��k[�]^	�	ۻv��}���I�y�����]�tǳ}p�;�k`�d�pRa2�ڏq�Y�8�z�!'���D�:�C.���G��/n��ʛ{G�58�#�w�� N��`D��,�6}ψ]B�!�Hc�<��9��L����V8�93����_|�ق}"��j�Ǵ�����ǜ#�]�C|����oo�Ǝ��pv2"<�_ރ�Ox�D� �-F����:�|�'�3����`M��?���^c�7z_�?������Y&�7x��a�1l��z_���A~�02fm��pD|e�!Bx�`_w,�n�b��p��� 6"3��蟜���@؊�Ch�/��7�=<�*���X����z�������(Z�j{�hX{z� ��(5^祥oӄ7>�>6��̀����u�r��n��6\;�WwZ�9�=C�\��bQ.�9C��i����iL�\+�dx|� ���� <�lT+�ɠ(3$��8d�8S��	s���N��g�U��%9�p�����"-6���D�8���� _����\��6�,�!;))��XY[GBD^zfV6Q����d���">/5m=��A:'� #�3���pZ�M�����D,��"�A����=���ق��#36���'|v$c������C`��<=���D���&tyy⍳����3��N��?��1B	���S$���{x�b)zF��g���'`|�ɹE�y�K������b��;�G���,sNzf�q�0��Ղ��[�0,����K������s�\�ￆ�`});]���p�֟}�&-��|�;��~[���o^��7(�|����|��o�qq��d0�
	����kdP��aX�R�#��5�����0+���"."�L�	Z����H�A���B��i�Qx��)Z�0�bQ^ׁ����8�u���ǐ�O���Em-
ӓ��/�YCb�<{����� ��{7�M�M�
���,����|W�ǿ�cxy���:2��������pQF�]���M2��8<4!<��a�س�ӌ����
���čƅ�`l3�?���,�Ŭ�4%ɿ��[[4z������~�,���d	;����l����ܽ�އ���3la�xm����i=&�y�+fJ��h��9�`vU�#�&�L��ǵ� ����1H��	G&�221��`dl����gW/��{j��x!c5:�0�z�B�g�3Z�h<�'7O?�|���!k����x_W��җ�p���u�B��i��H%�ŝ	O7+��\�M��M���ALR*���z�ˆv��0�ғRRӰ���H2���A�5Y�Յ�+ˋ��L�����6�L(#1c@��I���7.1(Z0��L�����&.2��e���\���Y��#lp��{�"a~�N��Z��A��7_��m +�XES���^�7.�&z�𬮁񊟏��K�8I��U��^t���֕2��"�W5��`�@=q�(�q𳹠������;�p�D>2Rb�+<Q�آ����3?;A^n���u���������/wW<�����.��q=(���U��yO���V����g�W߽E�?���5�<�4���n���xg��44Ɵ�v|��3��.Σ�c�y��˗x�|)���$,�*�9&<���s%�T�L�Y��g��nwH����I,���:uM	��dI&#�����d!BDG�--��\@j;�7�Ť�Yݠv�>�hǄPf�ܾ�z����54��Jnn&e�&��z3������E�v�h�gg&w�=����:��$�p������il��Xe v!���s���nr���.cՆz�>��ыZ�E�Āx���/^�r�<8GX�\��I����͝�8&+�3���Z����0A��aeN�#4�a��C�0E���{s��/y_Qgf>ׅ�0���_|x�������{t'��I�fHS���C�*�s��V �p���Ͳ@\��E��$xG������	k���ǚRq��p���� �F���������{��g��M�f^g������H����Kټl0l�Bc8����y��Л�`�6sA6	e|*�̓КE�E�� k�&����������0g'���fC&I�����,�j�و*��i$>F4��e}O>�\a&��<���3�kLp��?�Gc����4;:��f�Q\�6�y�b~e�k%p�����<�k�*�q6/�P�7�$�|N|�?�G)!&,�O�����G�0ۻ��d�"�q�K�8Ľ�F��id8��T�q�T5RSl#):��S�C�-���Ay�^�Ġ[���{nҢ��[�YIJz23��h�ޞ�i����"CB���'g�N�G+����p���GF9��y������N�cnv�!��f\xTߎ@/w\-����2�|�QV�O	%�V^�T�I�#3����q5E��](��۾�������,a��ST�;�'\�:_;�u����	�*�y��"ѓ��k'A)�QX(.�p�l��w?� �>�>�Q��JgW�?��
δ��S��ē������vw���W��ΡaĄ��g>��_�wn�CFt0^4��%�?}�.�÷Hs�Q��ɿc��M��	�M���rvRAMs/��\.��O&�V��a�TV"ic6Y�
�7�q�-5!��)D��4-=��ۈ����&�~��94�G�	u��ן�%����_� oW��=zFɲ>}�.���B�e�7�L/����"�������\[!�������A����hd��{B8�����.�����	���������~G]�NRrDz��&�zw77���ocg�A~�i�i�.�͕6u@(���K��q��'�a��3`��P#X1���y�Y�&�6S�7�O�X���?���
�"X�[Z��s��ye� �| �
]��-�c��}��<��P�Aؓ���D�Gs$lP�vP�X����D�$ɧ�+ܽ����� �MD�+� �Ãɦ<>�m�^ApY'�)��¶��!��9�IʜHO�0x��GG�އ���r�s�\�6�ɂ
{� �����9�:[������YD�}-�,Mx=����,k��Y0���E2&gl>fW���}�
�T�ί�[����Go�#Ut��n`0��",�l�Wϓn��͉\���k���"޹q��}	����n��"��A����Q\@��C8!;����?�Kt���4ą����L��&[;A�Gk��2�o�Pz[˿KOf#:2���L�Х���Ջ�%��H��/�����38�3���o߄߹�����dY����u.�z�F1K<���w@����>��(�%��q2��&�R�12¸ӏ��C�Ե�/�}�����<�������w��0f2xo��O��=�ƛ�^��L�Ih��++]q`hjF�(Z�qe+�����v�%�i&��@bh�ZxsG/ֶ�8�N���E��0��47��%��ه��UX��磣X"m�Tk�0����V�v�a�lǙ�qplN=��ᅚ��Iq�P狉��p�5=����f�m|a��}W:�Q�d5��ܿ|\I��ß�����]f��#�>�����D�����q��rb\�B0ɲ�%q�e|I����Y�x�仞шڹ�|}��
QĢ��@���%I���\���<�'gVu^Vy�C�2Α�9��Rz�`e��t~m]��}�l��γMW���uZ9Ap���A��'I豳u�GX���?�;�̂q_�%N���_��¤��	�mr��,��@c����B�����F���߁C3�vek� ��I-s��@���4	��k�S��>W���1J"�.C2+$�&�'�戋��cV�F�����I��E�(��W�zaA�Jww��k|?~��11�$__o���3Я��W�rzr<����G106� ~�""Bh��EtG``r�����'�#:8H�sln	/�:scÐ���yeu�鞢�S��Q@���ϸ���)������T����M]Z��
�Enz��D|�l��,TL`0N�&����/'�̯o ��%y�J]Rk8Ή�u�Zw\>��E���;h������^�X̅7b�L�cx\S*>�V�.�T5�̀�;<���~x�:��A�S��<\�J�����:ɀg��.�2c#q�#�x��I��\��kg��J�߸r������n�Çw�)���(���)�<_�G�h���+��2���9����g	�ǻ��%?��|Up@���G��V�}�1!^T��T����O�G�>�yrL��mvR,n�ע�oQi�D����%����%Fgx�ӚT���Ǆ��{/115��_9�L����4ꀗ��x�ء����$|���l-݃��I�j�S9���C^zZ&q���i�J�y��_�ٿ~zၾ��+��K���M���Z�'��E�ޓ�06���|t��u��k���p'�Z\����aˊ��*��IR�ļ����H����".2�3�L3����[�!��n!/9˫�!�����sSx��Y��gk,M�O����O06>�Yb���!6�fH�65׿F�YcpY������hafZ��ؼK�4:��2�1�'����ʁaz���&f�L֡r������m����u�������.ۑ�P�_���r��V�E�3OL�K�H��=�a ��U��R�ϯ���I�����5PD.��q�j�v�
I��ưZmʰ̪�%gg�����`?�[�L|�C���������vS]=m�����jusr~M�@rh��8�o�f��uܱ�;�u%_O/�39HLv����������E���,�X�\WR�o�c+�n.�X�!��k(�.�TF�

7;'kze��3��@R�5u��yoo^)� ��n����$����t�*����Ֆ =}	��� �����,'=��^�N�����kl�A!!1��%:��{H�3B�r";�W���::5�	Ԟ�a���F==,����a�0~t�{N��{7��I(����O��C2NW'#f��15���0?���y���DvIX���"c�!	��[e4T������q;����42Qg|p�BsEm-a�,�O%��`�p:"����&������jvb�~�}̦��u*t<��n�V�T6Q�ڍ�xɈ�et�Pc��pQ���O<v#FW7Ma|~E�H��b���6WԌ3�i���Dlq�n��k�Soq��OS�l6��u�1h�V�� ;A!��Ԅ@oo���c�
ܕ�f���IM3_�E��$.��X�a<��Ch` U=�ynUk>�v���zmj�4��D�H��c�(|aVc�~!&��}PQ�@���֗V7�yR%������3M7c��G� y�ƞa1�	�8����l%����"��;ֶ6`���;���Rd���mR��R񊸳s��F_W	��共�mHYT�<��Eb!�;j���*%� /)�K�h�]��X�#M�O/p���r�ɠB�B�@�&Y���L��vee�� ��P�����v�h�P��H���a�qd��RS�z�2R�<�-FI����J�P��V.��\�$88N�9B��������36��`s�hI�5:Q �hQ��6T�J..���T��4�j3�(����;��,����#:)��U�fǇ#5&J��C�ɒ;��I\��Q�N���&��}����!75A��'�ec�� B�=��+Z�9Y�Ă@�DU��̫h��K"�EY��u�k��4�%�.ϕv��������,��^��d�*H���=k���urD���L�w|6Z��L��>�Wa˅�y���ك���l�,��Y��yp���,�PA�'��˧r�����$�����g�Zm����+(+��������X��А,,.�LQ&�����d!+5�דe��߫��7���u2�rU���/ӝ-x��i,.�&�N����:u�w���B�=2��xR�̟'��ǅ����Ih�D#E��3��N�%����b[�(�{�'rP����9d$��K��IW�V�Zg&ģ�񡪹�s��A�45ۈܴd��%��4�0%��$	�<�EbT8I�.>�{14��/�PtN"6"����W��7���b�#12S��?|����2\%|
c���	��?�BY�7�j^O����� ��߹�82���i��E����i�{d_�!'%�um\���=�}|��(�BL�K�����!L~��30wpB����YK�r�vb�6g7at�h�������54���uZ�<=]�&��ͧV���0�E���u�Mi������q�C�3�͍��/nh:):\�Xz'!k�1KTxNZ�B���F�m0X���`��,�[���.&	Y�����T�����b���HO�3Y	�Ԇ�=��_��yx�A8��hU�Ѣ���I�d"��'�wB�7��@Qir�nAXgBOlB'x^���)5X]����m�ۡ�>d������D��OR4��\V�������F�����k�M2K/�^#Eն��p��)b�"R���{��։��(v�O�V�g�oPpI.*5&c�s�v��K�S��E#9< =C#���38A���RƑTL�I� ˺T���i�'��P�089M�LB �nrt�ΘB�0�'��Z���f��+�ı�Ee�[��"��+|�����©���J�E�0:I���*�}vz<~D�!8�k���-Mw����o^���L��a̝�r�����k�\��K��>cl� �}�{db�$�yD�oGk{;��Fv)��H{S��5�Զ�k���[��J؉V����S����D��AX�C�VmS7&8�V'Զ�"�4ؗn���G�]Tk,�%	��
b�N�q���:|������e�-���a���G]�M�9�	�܏iZ�$�%k#|J�t�ZhG���h���4Y��kml�EM���9�C3��=��%[���[4>JP�����Ć���M�9G��>�hBRT�4���)ؿ�?��E<!��"1gFY���S2���92K7�E�8�����V��i�ՒN�]^��Nh%���!���.����YYQo(~������n�z�CrvuV��&d�v��V�Oa&�`����5m����|�����J	���KJ��!����dVB� �@Ƒ�z8E\�]Z�f8)��f�B�Y�.�x�d�i0��u
YY2�Y�WH���+$ǌI,\�S(�����Pi��Ci�[���U����"ܦ�����KV�I�[$�O��^�����Ѿc�"֮�T2����2���H�u\���,$�m~��\:��RBue�Q!�ڞ)�M�=u"�h!�~��q��]�*V�BZ|�`Z���-�KF��EX���+YD�������{�"�S���G��`VM[���_*H����3����vj�]x���$;�J�J�._�5�Jޕ�����U�T#hq	�f+�e�dKlu� ��2��B(�����EJ��QWOf""П�aD[���{5R�)Hg���@�ZX^A%I��ޒ�d��s��N�إ�,'��4MY�:Y�gO��Wq&;i�I4�-eV�>�ԲD��bi�fz}�`��i��q�t68�B݊��+��ʋ^�r�T������
�,PȽ{��B8��H%�7u��}���#%U�ǩ�<Ba�C^�rJ��%�X���FB[#�YV)�c�Μ�X�t�O.�1fd���dg�X��oBV^z2�W4��Dy#���}DE�bI>>)�!EN@��EFR$���~��	1��=����I<|�΅��@������_>V8���.jEҠ:Ȍ��������5������v��?���"�cSH!3�?��r?x�
HL$ٚ����/����ӷ����B.J9�JN���%(�߹r��q�=�&�k[���.��w��'�k�a@��d��:����Ur�u��N���M���#�z��0<�@l ����I���&��"��;Q�K�ub~c��S��Z3ӵg����M�[�AB��6]�;K�aü��eqQ�
 �.o��s�֬��q�!���=��d8OB��v���Xi�u��5N�[����6TҊw	L�A��=��X��0;Q�6�(Wb��'���������C���//���M�%�ށ~��?Mz�5�fu�ʦ00sQa�><}��3>�-Xr�O�7LK�U�|H~�lV� ���R\���M�2�fĄ��o�0H�Z���Q�L��z�!n�*�JI��1"126}\��u�h�)�ON|$�Fp��]�����7��T��8�E����g&�j� 6ȏϙ��D?Wiv*��L62=��əY��G~����xjְ����Ҳy�6*�c��IZa�#�6'��݂��A�A̒�H���d�o��&��pf�dL\e<��a��[籽����PBV����y��-��߁���j�A�jj��{��0��b7����L+����%�Ȋ�6m p�B{�YӚf>�Zp2+!�h�dI��D�T������Fc�'P,�~^����(��%�M���_7���}����3Z�Ĭb�7yz3U� '؍�'��-R�P/O���NȎ8!B{ww��GG��?M6�t�)c��C�l�_�G�41��%�<�jD��7VfI��)|u� �u-�
 E�bl�����H�Z\h �v[�MO˾�����-
K�I�i��� �����qN���Jv��ϝ�����	�&�t��Ɗ��.��.�������gV�p��#�P�9W6�(���KYWJ��Y�8�g5]0҃$h[�R���C#����vp��)�Ւ�E+Y���/-Ɔ���������y)k��ࠗ�c��d?�X��/ae�\�ŕ�PaR�̎�Hu�0���9,�;	d�����dق AXJ������H��@X���V��֨%������dM6H"�F&�	�9���!����$M��*�Wa��J��	����IY���v�R���+WW�=J��Ƿ�q���H����3y�1����8��DqN*U��?�47�1�=���Fؘǋ�~�ݑ暄e�.��%Դwc�����8��jue\ZEy}'E��Ȋ���8��դ��d(n|�b|o��=NJy]'�c^����\@Y�����wɲL�I�Aq�p����.GWbyiV�M��$Ҝ�"�j��𠸔����Qe�R�-!��	!�"�6���upTc����pi���=�9���>��Sy�8`���ڗ����Tf2Rⰷ��F�9I�2�Rvb9��(d��~t���2�R�q��I��%�dBVyM�E���K\�����j����21=�P�⧘��������맑M8�c�-��eОE;�ѵ����:�q*+�o�b��].!ˊ�ӆ..j���'/P̅,H%��kD^V&:���Z{p�$�����i=r��Nv-�۹�YJɿx�HvOj���~��q�8�E���N�&,���W_�A~j8J
��aZ������K��@�r�3��^�njp���l�{�/�7�vm6O��O>������Ƴ9b�>R��_~�������h�B�����.'x���W��>�jAI~~��������Ù�||��Ε���>����!�u�4�5�8�ݦ��#�1b�I�x�x��O���h�ɰ ���l��EZw�"�]��P�:����"-)B��Y(�j�G11G��5�Ei������T�#�R��yĄ�i�A��F��k���_΢%Q�5���m���[�s���G�puG����8~�(��dU��X&Ď,l�4?����ލ3bC��Z,vmˁmȎ�=M��F#I�/�9n�`�>�Ĥ<so�d|��R��>WV�u.��Cm?0:�`������f㡶�n�]�l�� ૵!kvz87͸b��

��1`�M.�u�U��U-�+��*�Ec�+gO`�� %>�,gJ���`)��?�I)���6~�2��t�e%`�lG��v�p2A�QH�b�Ls����/��Aj�*R"�S&�����3������iEP��C�p"+�����n���&S[�.�DhH�B�0����p�A������'�롵���l�	}�x�r1<�h�dS�k�����;7N����b5b�Lp�
�J��&��������Zm�Xߦ'k�FBx >~R�y���o�>��3Ȍ��˖vlom�`߸z�(�~2��G�J����^>	�����JK�lZ>�Z��wUk7�3��C?� 8��k:��R��)Nj���E7kQ�%�Q)ϡ�wHsJ5dY�1H	�aanF�]�蒢�4�/241M+�����Q�>ّ�I/�x�F��Ӡ*��%�k7�$�{`|V�:�Âi�1PRS����D��`�����\rSۄ���vM�K��YO���c_<~�B���ݶN�R�ٹ_Y�Ҝ�長�Vc�Fh�'߫�E!ӓq��ǕJ�%�����/O��9B�.�?�l���i۪�oS�jg;Y��k6��>|�p���d'���b֣���Ik�$����T���$�6? {t��.�:��Am��ުj.�v��	�USҀ�I��b@��rvqR�#�����"���p�����0�h�0'�R�Ѥ[�9��O�;Bք�	krG'Ⱦ�ևu����
�F���u�1��\lѢ�\p�Ni�h%�����<u� Y)��%�Ml]ٔQat����tW�s�_���
y�v�4��h��q�����s�K#0�&v٤�L+ �;���!7-S� ����7��MdM.("�b��4�q1���f� Kqvr�}&M�D��3Ey�ts&+��.�]�Y��%)T��W5�R�����N�������./[�e�I��<ޫ!�(7Eu�����V��$�x� �|Y���L�>~^F���T:���W;ŨN�'!6�_�����M�i�����L������}x
�m=��eY	�(�J�r���5Z��)с�x��bsׁ;/�	q{H��3E�1O���n�vU&�[�],��$ˢ87��O�M����n��8�����{��|�1 ;���E��(�W;�����P�����$6�Ny�"m��4���9��|v�i�n(�d<�n���$�/]�(��Є⣺6��H��[(�n E���O�݊z\.�Q����WJ�E���H�l�o>-GQN<!$�?�CVR4��a���L��I���'z���D�r�bp�4��P$�0���'����S'��WT7E���������Λ��X�ܡ��ů>y���>���1hh�AfrY�=�l����<�k���"���G��	���PB�E8<w��������M.��a]?��f�3$�+�́��'-C\�%D�#�,kjr��� O�z�fF�(Mc�:�g�jtg��h��Ī�Н�7��00�3���dc�݊*���{�ѻ�t��r9ɡ��(�A���-����Ƅ��MjJe���C��ؠ@�'� TI�W��3:��`xf%�ч�q�-��Xs�1���5z7i!%#]X���Vh�vB���d�,=ka�Ax�����b�@�זNWi�.�d�4��ŜܼAܤ!o+�x�\Ê�p���w�Ɖ�L"�Ɂ$�|��dʜ��>���Bք�,<I+�^���e�B��8I+�	�\�,i�@���!V7/Zm�ޖn�[$�!1�B��ѩ��,p-�'`���8p��e��+�����:H�0�Uzjb���:kp��t�B�OmD�	�q��db�1>=�R
R?�@ąxacsKk3�E�	�~���v��˄�]Z�4W�v��ݭ��%vڑ��o�M���Ia%�����2��RE�� |��J)8� ���O��M�Ň��f�5��o�RF�����`��ek�����F1�i��0�E�#����q=�X,&�I�V�l���B������L�clFZ���f�&�r~��bّ��PQK
�09��7C<��KM�i	(N���N��8��¶�S�}�073����c�ſ���0owB�
�8��
�#���X=i���D��b�8Ş�������Q-,ɦ���.$FEb{c�Q����]�6u #)N	�}B�^0�U5�h}Cb�}2�9�讯^T�0-Q��O�0��
}PU���dx��p��CDi����s���A��*ϝ$.B��?�A��&��p�I̟?�Uvd�58;�Bv.o����%U;���DU|���t��RJ�&�e9��#�23�H�GY�������G�ʤ�Az���ĠU?�&
ŭ�rX�ɓ����\����i��;Ўt��{��+���5�?Z4��[����M-(#�����Aa9J���0��pi�3�d_���o�\�;��=Dؚ]����FM6�8H����#��YC�
W9���u�j�$�y}�e,a���w�ܗ�E�H���)/&�m�����C��&��|��S��i�CS��ks�e��j�10:���	��V
򒵃P����0��5߂��R�_!�ֵ��
�w�d|=\�9���DZ=�%Nd����ʲ�wG�P�wg�&<��&i��R�ϥr(��kIֶ�:�'Sb�	T�|�ʶA��$�BS���g3^���֮�&Γ���rom�
=i�(��J��U:.{Ȳ�v�C��I�������2?R锘P�2�nZ���.m8��Ǖ�\����q���#}+����Wo�'��Ƙ�@�+����2|��a���9�xAn��Gy�2����F��������8}�������B�XFt�&ℭ��_t�+�J�%�Fq^�Z�4�%�E);zTۆ)Ѵ2W3'"�dE���Iy3Hsq�y�s�P����/�u1�l���"�"�(-w�[��	O/��A�	��
���<�,�jq���$�Ĺ�T���K�� ��ǵ���s�>{ZoOW�D��_=������e _�!cBNJ~��.�>���U�r<ȩ�<���l����W�����SI8���Z&���_Ge�M�q�~��}�����%d�E���s������D/�ˍ3�0߯h�v+#�(�������y�#��CP�?����7��V��;�'��`2����}�dF6�aл�|lx���X0�V���pZΡ����ft�M�c��!��愇5�&+s�������v�Ѣ�w�y-〄#=)��L���16�m��)��,����x5��M�5���$28+�Ȧz��C��-'zi
<9_O�h�ó�p1;�p�(�Rf�1��P�ޢ`�����n��S=�R(��^s�glp������S�3�G�E���t�vh鰗2�Tݽ��[�͉�	�XCTto0��%�S��J�0!)
c���$��@�n�BVf<6�� �-�˜"K��'뉠u�($H�A���`EVl�n!������$�橋���#�U��ߟ;�/$G�Fz�7�D]�@yhrBZ���u��,�v��I�>��E�/���]�FJ�=�4�-P�,*�"��e�k��9����(ܢ�f��g�P����ǉ��컻���fr�f���.�������h"[+d��7y���&�c��Y��X[Z��7��52Wo�H -s��x�R�W,��`�T�ȕ�`��s�/\X�O\�e�a�1�kt��iE�XJ�9���+4q�+�{Gix�\i�,U��fhӋRp�d��MJ����J'���^͍��4���;1���.��ό�
��p�NK���EnbJ��6	�/����H?����eD�@��ԭ�:|��� ������Q݀�z&�m�m(L���o'�ە�V6�����[��GO(F�� cA�'�i����>�!<���fCek/�G'4���S��}\\u��&���<ù٪������_k�^����|�}�	�OT��ʠ�g|qc�+�gg�d��R�%�s�/�ۈ5���Ǻ��ae+�@�}��V����5%�NNF�$s�0�%)�4u��_��|,�*Z���'�M��Dd�r�����s�Ɨ��!UwS�(��B���	��-<D#?���l �(�2�nN�G赦�-
Ւ�'\I3ơV�yI����&�t��@N2G���:n?���C��j��h�A
m���*�v��N�Ɨ��u��	��4|����=xi<�Q��) eF�Vj�R�J��"���E�H�L>��l3�3�F��Ƹ &�qNF��n�����8��&����'��P�>�]�r�s��{�n^�9$]�\��0��>����A�N���,+���ty�\N���9G��磵��]���8����"54��m����M��
S�� I�I�����^BD0����%�-������	�n�8��>�!(�L����b.ѐ�d)�c.�Ȃ+��<E��F�3�y{�MB����P���)�ɾ�9�[z�t�Y����Hg��i�ޕ�\mz�%��O�b�3��u�8K;+��2N�ee2.4�/�������W��R"PC�*̊!4���/���DZ�I}�?�k�<k [KG	?�K�<Ku-���*�Dz�,�vU;�KKv���<'��<�|��ѡ82Y��ϐ���|���D2��_��@��eR�����ClT8>�ϱ���v�ei��dYܭB ��+g��Z[�L��s�X@#޼rZ��J1a���*<���K�[���jY!�_�gR���o���&G�ܸR���!�u�B��\?[�O��ҙS�'��l���'a��y69Ɂ�6��+K�l���G�IѦ�m4��IL���;����T�T	E�Tʟ�7��t~i�_>��4�2�K��kTvM�ֹ|ZW/<\]����227zϫ�"a'�n���&W�l�FRB�n��%;z\׍�a*sR�o^.�%{���sj	{G�ZB�S�̛h���U�W�B2�~�Җ�)}�4iz:)����	� 0�yΉvJR-&:a���?�g�>![
v�һ�����Umk�Z�Fi/�OL鑇s+��xbfV�iܭΨ�$�l��{�T��+�_��>@gw/�	q�_;z �,1W��d����#+����lEq)I�e2�Y���w4vH�zi�Lb@�߰#?9Tk��v�]V���/r�#���v�ߝx*�TF�R�Y��L~!���P�X\mȋ����'��� 3����	���+{ɦ��-Ɣ����;L�4AZ���'RC�&��%풙��҂�z����Mz�BY|�RC����~��mZ���.�΅���`ʂ��1��.�{����3d�kH�\�fr�&�������@v|��,��j�k
�;4�˄���qƏ]=���k����&J�����v�sK�.�tBuK��NJ����dER��c��F��eNn���տW�B(��7.�hZ���G��+:�9���^��IZ�� aS�A����I�;�Z��\�����h\�O ��&.�jN��w ���x�,[�z\��H$'�zP3�ϊ�i��Cȃ����t>#V3��� �k��\n���j��=��Gh�"��R����')Ix>���Q�j��I]��=�l��e=ΐ5y�y����#cz�ԗO�p�8�����n�uj����S.x6N�%`���E}ٗ3�<��؜�H����_<����,N��G�V�ԫ4�$/h�$ʶ腍]|�F�@B��`d'�7��g(�����ܔ�vv��`Ma'�����:R={�ء�R�rr���d�����1z|�-_z�t�
.��!91��c2Y�]�:�Q�9���Μd� ,$��֊���Po��12���9�x�Jg.����3$03�O�!�y�љu�3FIN�N/�J�(�0ˀ���Z�c2D�Yx�9�o��8Xz�I��=��>�<>�s$�[��_�F���0M��g��(Զ�
V�9��à���]0J�����ךM��Λ���j�4�q�ĲmdM��s�6�rd%��^rĆ�q��'`j�7c�@FɃ$�䨍B�@?��u��+��ּ�ąa�X�ő3����P�Ec��OZ��3D��3b���V3`� ;<$k
	@bl�nmn�F�J��Y����eh`��[��s:~9H�X������32�	� /�<_�Z��s@�n���p��	�/��:��|�=�֍��p�c�g����I?ƪ�^� ݭf��RE)_+��}�J�;_�//o���X�х�i�!�Z�F;��Bq�6�u���Y��4>S+�H*9u]�0Fq��K�H1YH�Y�ԋ��d=丱�%��%	x�kryMd` *�����dS�ds�zv�V3@��Ba&�z�D��4N���NDy�:���"���$,r��5�Ə6w7�!_4��x��l=�T���{=��&+����c�J[a�J��Nl0��q��q�]��+EK��.�ʥ��3.���B
�^�����\E1��������<(L��p��v����r�� �z������e9o����eđ�om�"2"?��Z:z���R�(�,�in>��~�v-��"��?6���@���K�qA�����}h��I�xI�$��~�z�֔�3���w�H�'n�%�B/��7�I�J����L��������}蜜��w6����IO��h���A�����nh>I�W���{�D�e�G�P����������ψY�>�z��yJW"�HM��ҒE�n�+�W���O��/Gz�WzBPd.���06�"��o[$:��H�	���I���<n���%Eyz2����VGgW����A	���l�Y�R;ř40��#f�~����N�@�	��� ��j�e���1���}#�j$���;��V��E�^ݣ%�讣C����IIZ��N�У�$�*�&��4�A6�'$�V�E�])a�D5�᧹$iё�[
��&\�y;��r���ZD��+�.z���3��DG!��4��E�S���!���<q��J����_��?�
�~�1V�=����4�˿�0�����Mִ����o\-���8�1��y���]ݓx�lm`؛,/Mw�JsanW)���P�����,-�H����NΈj��+�)أp�%�S���O.}Y�dk��6ٮ�`��p#�gϷ�^�E%��[K��\��b�zl�$�u�Q����4��^�2]��QC(,�|�t�6j������q��u�+�IZb�l�S=@��!�^/L�����'����y�B%�&<o��:'wc~��:���5�R�:�yj0!
��8+	O������#��ӜX�Yv��T9���*\.)�kZ4��uO���>n���eȏ	D��8��:(^M��,���gQ{B�ZEc���>�WN�yY�N����\�Х��d��D4h'����"�i��M�PB�k��R&]r>K|�O9@9BB��L_��.'B|I�6}�E$�Dٷ(�R����RaX&�x?ă�V�=���Y�X%�I��^e�@ /-�2IgK���}P7��Y��29cˌ�\�*�Ci���4]/��j-ٲ&���1=ܙ7�'+ծtix���D
M������pPqN.=�fra?��?�;h�^�#�R��~���&i����� �I����4!�%=�����P�:k���GL��c|�T��C����LK�X����TMG���x�W�D5/E���px���A���F�}GdA)�!��mp]��Z�K�����O'و4��o�ƞ� o�Q!w�Li~��.�� b�?��:ƨ+���ǅ�#��K�C;Y��H'���� �Ek�}xRi����	�Ҽ�98��PL���:9f]2ٓd���A��Y��������Q6�x��(+�q�L�"N��D�	PZpB��R�hwì�q�$|��G�-d����[���q�ݽ�0Gz���8ww(vV�vp�*7<0�X@V|���TC���zɉhS�	_K�90>�S�qRWϡ"�Q�4�O�(5Q$
��S��0=���} Y���������i]G��a���I�GSW?b(>�?n��b")&
5-}��$3�ã�D����Š�����+'2���&{7R�Lԓ�Fy�eeQ'5�:p���;*�рKder���N��wNcc��?/]�7ˉ��N��o���|���0��{�L1��$&�����rn�/F��*j���w�*�$���EL2�>�W�7����̸��o�zO��1@&+���������{W��I��@zR��ww��3����P)�mr��o��Ek�։S�+e��2��]��bgRT�ʾ���{M�h�Q�}��ˉA.&<O���pʂ��~�����׶�au �����)�}x�${������ԏ�� j�mW�]��9�����S{��1 a����;�U#	��\��o�zNo6�o��:|S���p�ӿxѤ�@?O=�_ח�彊v~����D��$��P^ۡ��M&uW�><)=�V�E���NB�ĘP44w���_~�f&'�l5���k�V1Y]	��X��7��
W�m��-��U�
���BhX0l>����9�C��`coaa���	��{���V�d󽜏��IB���]�G�4��5��� ���"",�/{�i
�qJ
���p]t�'�VI	S��3K��?=�G��d'RfjH0R���ɿ"[��£���`o�$�;ȡ��	qHKI�3�%��/�ןT��zj�ߍ��4һd��l�(;%)�uz��D�F�GMW\�y]����$=�+ZІhA�]�E,�`�0�Nb'�����N�ig�i3m�N�&]2I�8^H��lf�		�о�B����s�#0�C����}߽��{�A.����k�TS_���V����&n�T��~k����������c��pl�^�T����_]�M��a-t��˛M|���#����K��p��#B�MRJ��0ӄ)�^�gGO�?�ק�C�r�ڐ�4K��b��P�P�3 W��b�<k!%����\�t�.���\�v�-�2�O^/+�|�V�eS�E�N>R��R07�����	�xk�\$���rVC�Shni���b+���t2:�ߔP�LC\��61H��<�\�Y����'@�M{�f��@��䩉�����C�/�c�fxi���]�cL����������i��`Vk�ى34a�P���R7�[�D�QL;^���Uh#�s�x�2�z��k=�+����ԛ��Z����s��EM�!*��ǧ�@#Ģ�ĥ��|��f)X�4����i1/�ghTŬOT�R�C�d�����3���V>�ʥgF
~�/S]���Qqc?g�|��&tRn?j��o�j�xV�*�꧸��1��`�v�&�����i��ʴ��I���Jp��55�t�#��`�B��&�e���/���aZ�`�|q�����c'�b�0�?7k�0!�?�qhI��R��8�à�������v�d(�)P �;(ЊY��#�P� :?.��v�~�K�i7��I�DrP�DA	��I��NѨ"�Ni��\+Tj\��<S�~��R�)����dKs<$��S�/):��!�$1OL� [}��O�1]dp����Kr�d���T�W��m��)�hO� }T�Nl�k	���5Kh,!��#�����?�FPI�����~=�KBY��h���!44��CJW�3�S�;��6<�k\̢�+���]�XE'�$;�R'���&?�H�S�M����Ӎ��tܡ#�a��3?�v4�ݝV�S��Nm+2�������gل��A�y*3��QR����N����9ˠn��({�Nu�=�5KBq����{�V�����EE��1O����|��>���z!�^����W�		u9�����u��Y��"�6td޽~�տ{�c׶D������bl�n^���175ӗ�_��o�K��v��������N��J/����߅���x���!5Ճ���?�m���_-#�:y�0��ػk��Kk���?~sDJG�n��(	�/�Y������ؼ|1V.ˡ��1���'/���z���F��m�E}��k��aQR��W����ĕ��8s�r��q��hJ��-�u�\\�,|�2\}Ѐ��t�",���-,H�Ʒn� v~b"QV=N^�I?���I4�y|��#�Vt;�7�܇>���p�0�=�W(Q��f� 6�m�)����as0�ND�V�ɫw���u� ��g`��||�,<<�����lhWgWN_� �����J<�Q]��.ܩ���3�}���mbiR:�}���4�RpD����~FL��	a���EoBGWRM�����q�	�d ^�~��D��#%Ճu23�~��3�IMCRJ��a�`I�5H�,*6ʗ!`�+�#ȅ��DDФ)q�ԉ�=%p��/H���#�9N���H�g�a	?�)'6�~~jj
��n?#�J�HÒ�L�&/�K�L�W��njrq11��m�6gM�Y]��	��Ą��.��(��rI.F�{��GMm�eV��}C!��Z�q�qS�-��v�+D�^a�"�fm������Eh��DI�"8��.��TBt�^� ���1m���֬h<%)��{܈�ŋ���hl?UЦ� /1�XO4U� �4̯��W�N�Sʵ�;_S�q�('��;/,�Ar|$��zy�#�w��)Y�8�	�|#��D�x�*�e�R��u��)�}�T��J�r���`����I#�%�D��-KL��A}�ɻ��3/�����ƘEQ�L��4�I=�nYm	¦�~<��q����[��
Q�[�xO��mt�{��!A�h��滄�߸������l�)]���m�(_�����c��T-��O*T����ؿc#�W/5d�lj�1&���U�N�!��C���q߀��'-� �r:��0j��Tqk�� MZQ�w�dƕ&�#�;�rsQ��;13g����i��*�[��#��
#�{�߭&7��9?J9����9D1�Q��wf�i�`7��i>(��u���.߭E(���eg�����[z�J�H�@2��]N�*�H�c�\On7�5�j$�G�q���#;x�ݖSQ�!�M�qs�y�8�4и
�x�45����oO�h�@��]*gK"���;�}y	F�J(�% ����6�O6v��V�e���!�O������$�ꬍI���p"��a�͜��W��t��+(�6�/W�NպbK'%�v�d���Nɛ'ӌM�8Kw^I@�܁H��7�@�uص�9�EٍKe��c8E�"��CA٣�v{��찌� �ڵ�Y�n1<�����f|�54j�V�K��_h��1����aC�a��Y��E��+�������s�:Q�-� bg�zk��iT�����=�wrM����Y���v�j�'/߱&̕�&�*>nj�`�υ��LBQnFi��u����?������J�ݮy�:uE�+%����m�5Mt�1X����z��"�4cH��[M����ˎ���e��<���k�M�'$ԁ^�蛡<���.� Oba��X��r��`��p�M�ߵ��\�m���%�a�Z�)�`=��VZ^��]�o�|��5#��޺�4Mz������RG��� ���ʋ�0s���)���N�ӇG�]8�c��i��}h�K�vw�b�ܨ��ΑWw�Au+���˛����'����#e�!�w[T��_~|���_?��"�$e���cV�'2Z��NG��Jk)8q����DXk��r�H$���M��Մ�DMt���נ�AzL��~]���ڞ�E�/J�ї�Yǭ��l|��%�;.|����MI�'4���|t�>ʅ�݉�P7c�����h�g�÷ Cjq��Ó����-�4/�S⬙S���M��2�ˏ&9��y"��x�?8�9���$y�1>6CS��N���@dAz��@44�������И!/�@���!42����;@ ����.B�Vw0:��Ϗ��s�"�������>JO����6�o^l�E���^ڽ�M�z}s?T}R�PdB��!H��+�E:N/�[LR��6���>������g��%\U�BQ�>���LMKGb\�	�I�Z�F���N�&a���%�,:�e�Sb@�f����j-��Z2W���#��]�A��5a6�'��5�3�|�U�DE2F0�di��G��H����C#�P!�0/�?H��^�O{(�塷�3RMIH�e�ɯY���z���O�~�Nauq�:��
r�<\���2�'�_3���n�߼]}}XLHy����1u�<�K�?2n���h6�S��8#y��H"r�xPg��l��	�J�5ַ�K���A�[V	16p�VM���i,���HM,2���*�G�-�+{}�2�pћ:�@�V��x����Nс&�~ƨ}i��n)6����oy(e"�b�q�t���*祩S��;�{����h�5�U~Gu�^*�fG����6����m����ً�{��t��f��b�^Hs>�s7�Z���/Λ�t����?}��|����62vX�k ʲNZn�Oա�A�.�VUr3F�Xn���i��<�ͪ��A�j��ft����d-��F\��Y�c.	T��7�)K�^hG��!�X����Kq4/�7ˁ
Xh
υ��
����0�:�f���y�mT���nMΑ;w�>�3Ȫ���ƟR��k4O�N�����l`���O��Z,�����]���K�J�$��h�ʽGF�Q�8�|��Ճ:��X�k����`����PW�d����Q��@��Ԋw~�17���#�&�ͭ=����G��s��y���J�zZR7�7��'����`Ф���r��#����О����(X��?�2�_�N<;=b,v�\ u� ޔZ���,����������c%����O�#c029fܬ9�Y1p
x>�O#�{�>���,�ʦ����E��������9AQ�g��-"��(pU�Vm�w�s"�'_����18fp8�k�~e��UO����6�hi˚%��=T�6�O��}8�}��߻t�**���O�������^�S��}��-�G�nT?uQ�<��K'K�V�Kғ��2'˺NCi��^�D/<5.V䡟'#��^c���p+]� ���j�C�nK�k�ZGW���I-������/a�'@����}�'KY޲�+���B�-A��W���i��]��r%�*��%���s0&�'�=���VBRAgF4($�����ly�t����$����/�Xgؾ�k1Σ�y6���-��'.2�Þ� xx�ނw?��L��vmEτ��{�JF����kG�'���C��$��Y<"�}��>�2�����-p���&���M���]����8v�:j(�Q��K۴2t<��m�чx��kI�"��J,/X�/.W2�{����XS�c��Y錾��jPR��eO�ܲ�Sp�������!�ç��|�qh&����UӘ����D==HK����{��CR\���N�y�J 
��a��WˌO%��Å����0����o��w���o?G�s
��>,�C����:?��G&*���ްZM}s�B���w>�wz?��Dav&f����7�����k��Z�B#�������A^k�UM�x�1F4%q�ŋ����A��3go�;ޏ��Ip�����{��jA�� �]AƖH���H���a�	��.���ܹi�.7"�%��`��s�����NLA Q��s���U�22��S�<P:�Vb�<k&uH����������Hz>{�ߚ�������&ЂC��;�)Q��on��j.s������J�մ�:Ӯ��0� &@�:i%&0I��v��EɘG4Os��ӄQ|���a:c���M?:&�q��z[:;�(U�L�wI�C�^ݝn>��D��wӿ�����@7����\W�	�g�&2�|hzCk;^\�O�<�%�zU-��@�qm_����y6ҧ�ӫ���) �p7�te����&cq&�x�<���#^__���i��Ѭb�k�A�$�/]j�:��e5u��H�o_cC\ԫ2J���vo��V��osg7�G�,5?��.7g����!��C��zY�AgUD�ۻ��f��҈o�-��W��)�ӏU=�Û�׃ቱ:��Va�3�������6�VBdWnU�<��+�8�m-}�j��.�a,��ş.�،9ާ��߱9��~|�wn6���R>����ś�hF�KR�X��Q��T��5e>n�Є��]�Q�c
n�>f�+��2���	�6��[�]d6��Q��b���oW[J�3�J�*1�`B�	|Ej��jז�����W2����Ҭ���8��s�ם�o7-:h����bϠ/( ���������[k��ڧ��"E
��k����|6`�S���7�Q��T�T<#�JMq3#v���ߨu�z�N��J�ω�χ/��i��\�	@������_�knx�q�5�oU4cGUhJ���	���ֈ!_�T����ӎ���Ú-�F�K�^�ii�E�>*g����&�'E�oc�%���E��wX�Ȍ58|�.y�I�;�\�k5y�"��S��L��v�(����7xg�>�h.\����+�H���B]7b���n0���D3���^t=��p;��O�,s��v�����)@H���j��tZ�5.*�_�f!���&>�u�`��������DrXe���؄ɬN����J��{�V\eui�i��,�����+�u�>%�6E�� ��{�GXd�O� w� ����ʢhg��xJn��5v�����x3h���TM��	���#?/.�l�~��Zb��j~IM�Ŋ*�[W��Ѓ��k��*[Uh�5�Hǝ���]�{۳e�@0��4V�\����K���������S��O^@7O��ݛ��xJ�Z��l���ϣ�&W�����=�x��n��/��҆���@EuF\�qh�ua=ih�+�������N����p~x��iWl[���t\�����E�Pq߄�voX��K0���6�����Q�2���:Q��LF�u(g����`�*礧��'���X�d!vnZ���N��t3��ßnX��^F�}�m<���{���X�[�POs8�J�<N{��_م�H�a�9��o�}n��￹iI	�������ǭ���sq1���E��q�"�����/��8�;���0H��?�՛(�Y���m�����}H�>���íg�����ѯNV{L�w�2�4�!Q���y��#Le���X��}u��CXC?���h��	o�z��8JW/�s�I{ʈqx�;ڍi� �O}S��	OB�M�ۋ)�@���x OX<:��y�1��υ1g8������7��&n�y=JL�3Gc�~����L�ET6N$7��L;����M�����1:cҭ#����@D�Ϥi�b��~����tc��LI穘� ��D�%��aL��'��ٌC.S��1����K�j��w�/��A��ϙ#*��ώ�:0�?S��,�����e����;y�A������	��%�mC'c��i�e/��`o'�C�v��\Z��a��ġ�Q'�g�"B]�� ��Ց)�p��'��M��X@�����_>�D��a����~�\��N�R�&����ET����S����}I��Q�hb&�I#{'_/���Kfpj�9a���n��fRG�A����1�����Φ��[͙�wL������Q5�hl��V˹C�0�:l�1�Y��
�vʈ�����\x�(�����ǌ(w��9"q���]�{�1�����y?Zf��r��{� &�q2:�ol��f�bL4�"�����K���7v"pr�"����t�,N�����+�s������x��3�,(���/}�M���n����U    IEND�B`�PK 
     �8�ZuaKbH bH                  cirkitFile.jsonPK 
     �8�Z                        �H jsons/PK 
     �8�Z�֎�?  �?               �H jsons/user_defined.jsonPK 
     �8�Z                        ߈ images/PK 
     �8�Z	��} } /             � images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     �8�Zd��   �   /             c images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
     �8�Z�Xw�s� s� /             ;' images/49baae61-cb81-429b-96a1-6cfb8f124b59.pngPK 
     �8�Z��X��&  �&  /             �� images/9c69fbd4-c376-47ca-8b4c-793dd402431a.pngPK 
     �8�Z���*6 *6 /             #� images/a1588c66-a70c-44df-b30c-55fdbd854069.pngPK 
     �8�ZIRP4#  4#  /             � images/2dd92824-eee5-446a-82e5-cb3be823b6e8.pngPK 
     �8�Z�&�y`  y`  /             < images/8c2f1315-cf23-4ba8-a920-becb97f13280.pngPK 
     �8�Z�����  �  /             � images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.pngPK 
     �8�Z�Lz��L �L /             � images/256658b1-ffe9-46c3-9f0b-70052a8fe00d.pngPK 
     �8�Z9?B��  �  /             � images/d18021d8-4522-4af4-a3c6-358ee97fa8ad.pngPK 
     �8�Z�IQ�H� H� /             F	 images/a05d3615-68b8-4f26-98d6-1aedf7f6d878.pngPK 
     �8�Z��[?:  ?:  /             �� images/b75f5fea-d559-4623-b1ce-f8cd504066c2.pngPK 
     �8�Z��z� z� /             g7 images/00f35920-432a-4227-a0de-f9ff33566dcd.pngPK 
     �8�Z���1�_ �_ /             . images/fce5a045-7211-4fa3-86b3-f57a3d8041ae.pngPK 
     �8�Z�J��T  �T  /             tn images/91777b75-38f2-4118-94bc-a70a6868aa47.jpgPK 
     �8�Z"9��T  �T  /             �� images/0b0a0ee7-c404-40e4-9217-cd21fece1ba1.jpgPK 
     �8�Z�|��b� b� /             � images/ed998360-ed4f-472d-a3e6-52adfa722a6d.pngPK 
     �8�Z�GR�8  �8  /             b�" images/08988072-c7a8-475c-9331-8aa77c72a02a.pngPK 
     �8�Zj���� �� /             W�" images/3281a32a-bb08-42cb-a591-9481e2c9eb0d.pngPK 
     �8�Z��I2\k  \k  /             G�% images/35c60fd9-1fb3-48b8-b3d7-7968b0279531.pngPK      /  �:&   