PK
     eO�ZYQ���  ��     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9"],"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0"],"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6"],"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7"],"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8"],"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0":["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5":["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6":["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7":["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8":["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9":["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0"],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14":[],"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15":[],"pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"],"pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"],"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13"],"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1"],"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"],"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12"],"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2"],"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7"],"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11"],"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8"],"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3"],"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"],"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6"],"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2":["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10"]},"pin_to_color":{"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2":"#0a0a0a","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1":"#f70202","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3":"#0300b3","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4":"#0cdf2f","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5":"#b6c11a","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6":"#5df4e2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0":"#f70202","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1":"#f70202","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2":"#f70202","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3":"#f70202","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4":"#f70202","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5":"#5df4e2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6":"#0300b3","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7":"#0cdf2f","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8":"#b6c11a","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9":"#0a0a0a","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10":"#0a0a0a","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11":"#0a0a0a","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12":"#0a0a0a","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13":"#0a0a0a","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14":"#000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15":"#000000","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0":"#5df4e2","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1":"#f70202","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0":"#0a0a0a","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1":"#f70202","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2":"#5df4e2","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0":"#0a0a0a","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1":"#f70202","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2":"#0cdf2f","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0":"#0a0a0a","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1":"#b6c11a","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2":"#f70202","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0":"#f70202","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1":"#0300b3","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2":"#0a0a0a"},"pin_to_state":{"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2":"neutral","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1":"neutral","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3":"neutral","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4":"neutral","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5":"neutral","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14":"neutral","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15":"neutral","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0":"neutral","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1":"neutral","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0":"neutral","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1":"neutral","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2":"neutral","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0":"neutral","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1":"neutral","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2":"neutral","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0":"neutral","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1":"neutral","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2":"neutral","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0":"neutral","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1":"neutral","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2":"neutral"},"next_color_idx":13,"wires_placed_in_order":[["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_23","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_22"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_35"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21"],["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"],["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6"],["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_bd8b6d2d-60e6-4b66-abf0-62afb810491d_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1"],["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_23","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_22"]]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_35"]]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21"]]],[[],[["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20"]]],[[["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21"]],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_21"]],[]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_20"]],[]],[[["pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_22","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_23"]],[]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_2e0aaba8-f3e9-4089-92f9-fdf2a0b41a97_35"]],[]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"]]],[[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"]],[]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4"]]],[[],[["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6"]]],[[],[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_bd8b6d2d-60e6-4b66-abf0-62afb810491d_0"]]],[[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_bd8b6d2d-60e6-4b66-abf0-62afb810491d_0"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2"]]],[[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]],[]],[[["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]]],[[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]],[]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1"]]],[[],[["pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2":"0000000000000001","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1":"0000000000000000","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3":"0000000000000004","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4":"0000000000000003","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5":"0000000000000002","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6":"0000000000000005","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0":"0000000000000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1":"0000000000000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2":"0000000000000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3":"0000000000000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4":"0000000000000000","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5":"0000000000000005","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6":"0000000000000004","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7":"0000000000000003","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8":"0000000000000002","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9":"0000000000000001","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10":"0000000000000001","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11":"0000000000000001","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12":"0000000000000001","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13":"0000000000000001","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_14":"_","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_15":"_","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0":"0000000000000005","pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1":"0000000000000000","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0":"0000000000000001","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1":"0000000000000000","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2":"0000000000000005","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0":"0000000000000001","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1":"0000000000000000","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2":"0000000000000003","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0":"0000000000000001","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1":"0000000000000002","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2":"0000000000000000","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0":"0000000000000000","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1":"0000000000000004","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2":"0000000000000001"},"component_id_to_pins":{"2382caf0-f704-45b0-afc9-19555c232ea2":["2","1","3","4","5","6"],"413adb9e-60b4-4310-bd72-e4e11d56ccb2":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"],"1cb3a49d-dc66-4fa6-8d47-aea3068df0b4":["0","1"],"7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c":["0","1","2"],"6709695f-c694-4d3b-8888-654e702eb44c":["0","1","2"],"ff0891dd-490d-4f7f-b028-abe315436194":["0","1","2"],"9160c2c5-ef89-4fab-911c-be70a3060d8a":["0","1","2"],"686232c8-bdc9-4b03-9791-f090cd6c7e85":[],"470753c0-2a44-41d6-b577-b515fa83a749":[],"17669cf5-00f7-487e-af61-6dc7cec32cac":[],"78042b3a-f2f8-4275-8b35-53f2a17714ef":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0"],"0000000000000001":["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2"],"0000000000000002":["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8","pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1"],"0000000000000003":["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7","pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2"],"0000000000000004":["pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6","pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1"],"0000000000000005":["pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0","pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6","pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5","pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[1110.2200060000005,175.944395],"typeId":"22281399-816a-4a45-b5b7-1546df80d2bb","componentVersion":1,"instanceId":"2382caf0-f704-45b0-afc9-19555c232ea2","orientation":"right","circleData":[[977.5,185],[977.7218695000001,155.00578700000005],[977.3354725000002,229.19248100000004],[977.3354725000002,243.10244150000005],[977.7218695000001,258.1716545],[991.2454915000001,287.53722500000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[511.8908200000001,204.4938005],"typeId":"a634ff83-abbb-414f-80bc-066b6f1a8bb9","componentVersion":1,"instanceId":"413adb9e-60b4-4310-bd72-e4e11d56ccb2","orientation":"up","circleData":[[602.5,215.00000000000003],[602.3500000000001,236.0000000000001],[601.9000000000001,259.33399999999995],[600.25,282.66650000000004],[603.6670000000001,306.0005],[532.1335000000001,306.0005],[509.16700000000014,306.0005],[487.0000000000001,306.0005],[464.83450000000005,307.1675],[602.5,143.834],[603.6670000000001,119.33449999999999],[602.5,98.33449999999999],[602.5,77.33449999999999],[601.3345000000002,52.833500000000015],[533.6671585000001,283.83383000000003],[580.3338265000001,304.83383000000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"version":2,"id":"Resistance","label":"Resistance","description":"","units":"Ω","type":"decimal","value":"4.7","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Resistance","unit":"Ω","required":true,"validRange":[0,70000]},"Tolerance":{"version":2,"id":"Tolerance","label":"Tolerance","description":"","units":"","type":"string","value":"5%","displayFormat":"dropdown","options":[{"label":"0.25%","value":"0.25%"},{"label":"0.1%","value":"0.1%"},{"label":"0.5%","value":"0.5%"},{"label":"1%","value":"1%"},{"label":"2%","value":"2%"},{"label":"5%","value":"5%"},{"label":"10%","value":"10%"}],"showOnComp":false,"isVisibleToUser":true,"name":"Tolerance","required":true},"Number Of Bands":{"version":2,"id":"Number Of Bands","label":"Number Of Bands","description":"","units":"","type":"string","value":"5","displayFormat":"dropdown","options":[{"label":"4","value":"4"},{"label":"5","value":"5"},{"label":"6","value":"6"}],"showOnComp":false,"isVisibleToUser":true,"name":"Number Of Bands","required":true}},"position":[528.299914926406,239.30827804023798],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"1cb3a49d-dc66-4fa6-8d47-aea3068df0b4","orientation":"up","circleData":[[512.5,260.00000000000006],[542.5,290.00000000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[318.2035,528.6544999999999],"typeId":"6500d8ea-11fe-42e2-8a9f-99be354012a7","componentVersion":1,"instanceId":"7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c","orientation":"up","circleData":[[212.5,560],[222.44650000000001,567.7579999999998],[240.05050000000006,567.1609999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[570.165334,616.4889995],"typeId":"8e0ee0b2-778d-4065-bf79-38edea29856f","componentVersion":1,"instanceId":"6709695f-c694-4d3b-8888-654e702eb44c","orientation":"up","circleData":[[497.5,665],[507.055,672.077],[517.3165,677.7395]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[43.31500000000004,434.6300000000002],"typeId":"6d0c07c0-db0e-4413-b9a4-ee378c2ed587","componentVersion":1,"instanceId":"ff0891dd-490d-4f7f-b028-abe315436194","orientation":"up","circleData":[[-87.50000000000001,485],[-81.25249999999996,496.5335000000001],[-73.08349999999997,506.8655000000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[801.3969999999999,646.5035],"typeId":"1cec4e8a-72c2-4b6a-9a5c-b6be0dc427d1","componentVersion":1,"instanceId":"9160c2c5-ef89-4fab-911c-be70a3060d8a","orientation":"up","circleData":[[812.5,695],[820.9989999999998,687.0725],[829.7424999999998,679.31]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Turbidity sensor","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[57.96696427243663,531.1244549982175],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"686232c8-bdc9-4b03-9791-f090cd6c7e85","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Temperature Sensor","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[292.2231314606828,614.5459012322258],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"470753c0-2a44-41d6-b577-b515fa83a749","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"PH SENSOR","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[550.8560026663338,727.7651803249732],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"17669cf5-00f7-487e-af61-6dc7cec32cac","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"TDS SENSOR","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[772.1681606443491,794.1359304792926],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"78042b3a-f2f8-4275-8b35-53f2a17714ef","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-99.61020","left":"-101.68500","width":"1487.45961","height":"922.24614","x":"-101.68500","y":"-99.61020"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#f70202\",\"startPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0\",\"rawStartPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_1\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"977.7218695000_155.0057870000\\\",\\\"977.7218695000_215.0000000000\\\",\\\"602.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#f70202\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_0\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_215.0000000000\\\",\\\"602.5000000000_236.0000000000\\\",\\\"602.3500000000_236.0000000000\\\"]}\"}","{\"color\":\"#f70202\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.3500000000_236.0000000000\\\",\\\"602.5000000000_236.0000000000\\\",\\\"602.5000000000_259.3340000000\\\",\\\"601.9000000000_259.3340000000\\\"]}\"}","{\"color\":\"#f70202\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"601.9000000000_259.3340000000\\\",\\\"602.5000000000_259.3340000000\\\",\\\"602.5000000000_282.5000000000\\\",\\\"600.2500000000_282.5000000000\\\",\\\"600.2500000000_282.6665000000\\\"]}\"}","{\"color\":\"#f70202\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"600.2500000000_282.6665000000\\\",\\\"602.5000000000_282.6665000000\\\",\\\"602.5000000000_305.0000000000\\\",\\\"603.6670000000_305.0000000000\\\",\\\"603.6670000000_306.0005000000\\\"]}\"}","{\"color\":\"#f70202\",\"startPinId\":\"pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"rawStartPinId\":\"pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_1\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"542.5000000000_290.0000000000\\\",\\\"542.5000000000_305.0000000000\\\",\\\"603.6670000000_305.0000000000\\\",\\\"603.6670000000_306.0005000000\\\"]}\"}","{\"color\":\"#f70202\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"endPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_1\",\"rawEndPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.3500000000_236.0000000000\\\",\\\"580.0000000000_236.0000000000\\\",\\\"580.0000000000_170.0000000000\\\",\\\"227.5000000000_170.0000000000\\\",\\\"227.5000000000_567.7580000000\\\",\\\"222.4465000000_567.7580000000\\\"]}\"}","{\"color\":\"#f70202\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"endPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_2\",\"rawEndPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"601.9000000000_259.3340000000\\\",\\\"572.5000000000_259.3340000000\\\",\\\"572.5000000000_177.5000000000\\\",\\\"445.0000000000_177.5000000000\\\",\\\"445.0000000000_680.0000000000\\\",\\\"507.0550000000_680.0000000000\\\",\\\"507.0550000000_672.0770000000\\\"]}\"}","{\"color\":\"#f70202\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"endPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_3\",\"rawEndPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"600.2500000000_282.6665000000\\\",\\\"625.0000000000_282.6665000000\\\",\\\"625.0000000000_155.0000000000\\\",\\\"-117.5000000000_155.0000000000\\\",\\\"-117.5000000000_506.8655000000\\\",\\\"-73.0835000000_506.8655000000\\\"]}\"}","{\"color\":\"#f70202\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"endPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_4\",\"rawEndPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"603.6670000000_306.0005000000\\\",\\\"655.0000000000_306.0005000000\\\",\\\"655.0000000000_755.0000000000\\\",\\\"812.5000000000_755.0000000000\\\",\\\"812.5000000000_695.0000000000\\\"]}\"}","{\"color\":\"#0a0a0a\",\"startPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9\",\"rawStartPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_2\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"977.5000000000_185.0000000000\\\",\\\"767.5000000000_185.0000000000\\\",\\\"767.5000000000_143.8340000000\\\",\\\"602.5000000000_143.8340000000\\\"]}\"}","{\"color\":\"#0a0a0a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"603.6670000000_119.3345000000\\\",\\\"603.6670000000_117.5000000000\\\",\\\"602.5000000000_117.5000000000\\\",\\\"602.5000000000_143.8340000000\\\"]}\"}","{\"color\":\"#0a0a0a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"603.6670000000_119.3345000000\\\",\\\"602.5000000000_119.3345000000\\\",\\\"602.5000000000_98.3345000000\\\"]}\"}","{\"color\":\"#0a0a0a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_98.3345000000\\\",\\\"602.5000000000_77.3345000000\\\"]}\"}","{\"color\":\"#0a0a0a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_77.3345000000\\\",\\\"602.5000000000_52.8335000000\\\",\\\"601.3345000000_52.8335000000\\\"]}\"}","{\"color\":\"#0a0a0a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13\",\"endPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_13\",\"rawEndPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"601.3345000000_52.8335000000\\\",\\\"601.3345000000_5.0000000000\\\",\\\"182.5000000000_5.0000000000\\\",\\\"182.5000000000_560.0000000000\\\",\\\"212.5000000000_560.0000000000\\\"]}\"}","{\"color\":\"#0a0a0a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"endPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_12\",\"rawEndPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_77.3345000000\\\",\\\"602.5000000000_80.0000000000\\\",\\\"302.5000000000_80.0000000000\\\",\\\"302.5000000000_447.5000000000\\\",\\\"430.0000000000_447.5000000000\\\",\\\"430.0000000000_665.0000000000\\\",\\\"497.5000000000_665.0000000000\\\"]}\"}","{\"color\":\"#0a0a0a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"endPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_11\",\"rawEndPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_98.3345000000\\\",\\\"602.5000000000_95.0000000000\\\",\\\"-102.5000000000_95.0000000000\\\",\\\"-102.5000000000_485.0000000000\\\",\\\"-87.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#0a0a0a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"endPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_10\",\"rawEndPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"603.6670000000_119.3345000000\\\",\\\"603.6670000000_125.0000000000\\\",\\\"677.5000000000_125.0000000000\\\",\\\"677.5000000000_740.0000000000\\\",\\\"829.7425000000_740.0000000000\\\",\\\"829.7425000000_679.3100000000\\\"]}\"}","{\"color\":\"#b6c11a\",\"startPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8\",\"rawStartPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_5\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"977.7218695000_258.1716545000\\\",\\\"910.0000000000_258.1716545000\\\",\\\"910.0000000000_432.5000000000\\\",\\\"464.8345000000_432.5000000000\\\",\\\"464.8345000000_307.1675000000\\\"]}\"}","{\"color\":\"#b6c11a\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8\",\"endPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_8\",\"rawEndPinId\":\"pin-type-component_ff0891dd-490d-4f7f-b028-abe315436194_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"464.8345000000_307.1675000000\\\",\\\"464.8345000000_267.5000000000\\\",\\\"-80.0000000000_267.5000000000\\\",\\\"-80.0000000000_496.5335000000\\\",\\\"-81.2525000000_496.5335000000\\\"]}\"}","{\"color\":\"#0cdf2f\",\"startPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7\",\"rawStartPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_4\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"977.3354725000_243.1024415000\\\",\\\"895.0000000000_243.1024415000\\\",\\\"895.0000000000_417.5000000000\\\",\\\"487.0000000000_417.5000000000\\\",\\\"487.0000000000_306.0005000000\\\"]}\"}","{\"color\":\"#0cdf2f\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7\",\"endPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_7\",\"rawEndPinId\":\"pin-type-component_6709695f-c694-4d3b-8888-654e702eb44c_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"487.0000000000_306.0005000000\\\",\\\"487.0000000000_290.0000000000\\\",\\\"452.5000000000_290.0000000000\\\",\\\"452.5000000000_695.0000000000\\\",\\\"517.3165000000_695.0000000000\\\",\\\"517.3165000000_677.7395000000\\\"]}\"}","{\"color\":\"#0300b3\",\"startPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6\",\"rawStartPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_3\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"977.3354725000_229.1924810000\\\",\\\"880.0000000000_229.1924810000\\\",\\\"880.0000000000_402.5000000000\\\",\\\"509.1670000000_402.5000000000\\\",\\\"509.1670000000_306.0005000000\\\"]}\"}","{\"color\":\"#0300b3\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6\",\"endPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_6\",\"rawEndPinId\":\"pin-type-component_9160c2c5-ef89-4fab-911c-be70a3060d8a_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"509.1670000000_306.0005000000\\\",\\\"509.1670000000_410.0000000000\\\",\\\"632.5000000000_410.0000000000\\\",\\\"632.5000000000_770.0000000000\\\",\\\"820.9990000000_770.0000000000\\\",\\\"820.9990000000_687.0725000000\\\"]}\"}","{\"color\":\"#5df4e2\",\"startPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"rawStartPinId\":\"pin-type-component_2382caf0-f704-45b0-afc9-19555c232ea2_6\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"991.2454915000_287.5372250000\\\",\\\"940.0000000000_287.5372250000\\\",\\\"940.0000000000_507.5000000000\\\",\\\"532.1335000000_507.5000000000\\\",\\\"532.1335000000_306.0005000000\\\"]}\"}","{\"color\":\"#5df4e2\",\"startPinId\":\"pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0\",\"endPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"rawStartPinId\":\"pin-type-component_1cb3a49d-dc66-4fa6-8d47-aea3068df0b4_0\",\"rawEndPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"512.5000000000_260.0000000000\\\",\\\"535.0000000000_260.0000000000\\\",\\\"535.0000000000_282.5000000000\\\",\\\"532.1335000000_282.5000000000\\\",\\\"532.1335000000_306.0005000000\\\"]}\"}","{\"color\":\"#5df4e2\",\"startPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"endPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2\",\"rawStartPinId\":\"pin-type-component_413adb9e-60b4-4310-bd72-e4e11d56ccb2_5\",\"rawEndPinId\":\"pin-type-component_7ebe35a4-ffcc-4ac1-9f1d-a3604f68747c_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"532.1335000000_306.0005000000\\\",\\\"532.1335000000_282.5000000000\\\",\\\"242.5000000000_282.5000000000\\\",\\\"242.5000000000_567.1610000000\\\",\\\"240.0505000000_567.1610000000\\\"]}\"}"],"projectDescription":""}PK
     eO�Z               jsons/PK
     eO�Z�o�r*  *     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"vega iot","category":["User Defined"],"id":"22281399-816a-4a45-b5b7-1546df80d2bb","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"5de4bec6-ccea-4571-acb8-2cf876e4e4fc.png","iconPic":"f4826ebb-d8ab-4c3e-8d6e-ffd2265d28af.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"35.40728","numDisplayRows":"35.40728","pins":[{"uniquePinIdString":"2","positionMil":"1830.73470,885.56396","isAnchorPin":true,"label":"gnd"},{"uniquePinIdString":"1","positionMil":"1630.77328,887.04309","isAnchorPin":false,"label":"5v"},{"uniquePinIdString":"3","positionMil":"2125.35124,884.46711","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"4","positionMil":"2218.08431,884.46711","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"5","positionMil":"2318.54573,887.04309","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"6","positionMil":"2514.31620,977.20057","isAnchorPin":false,"label":"GPI/O 25"}],"pinType":"wired"},"properties":[]},{"subtypeName":"PCB","category":["User Defined"],"id":"a634ff83-abbb-414f-80bc-066b6f1a8bb9","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"3281a32a-bb08-42cb-a591-9481e2c9eb0d.png","iconPic":"35c60fd9-1fb3-48b8-b3d7-7968b0279531.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"25.12926","numDisplayRows":"23.63459","pins":[{"uniquePinIdString":"0","positionMil":"1860.52420,1111.68817","isAnchorPin":true,"label":"5V"},{"uniquePinIdString":"1","positionMil":"1859.52420,971.68817","isAnchorPin":false,"label":"5V(PH)"},{"uniquePinIdString":"2","positionMil":"1856.52420,816.12817","isAnchorPin":false,"label":"5V TDS"},{"uniquePinIdString":"3","positionMil":"1845.52420,660.57817","isAnchorPin":false,"label":" 5V TURBI"},{"uniquePinIdString":"4","positionMil":"1868.30420,505.01817","isAnchorPin":false,"label":"5V TEMP"},{"uniquePinIdString":"5","positionMil":"1391.41420,505.01817","isAnchorPin":false,"label":"GPIO25  TEMP"},{"uniquePinIdString":"6","positionMil":"1238.30420,505.01817","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"7","positionMil":"1090.52420,505.01817","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"8","positionMil":"942.75420,497.23817","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"9","positionMil":"1860.52420,1586.12817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"10","positionMil":"1868.30420,1749.45817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"11","positionMil":"1860.52420,1889.45817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"12","positionMil":"1860.52420,2029.45817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"13","positionMil":"1852.75420,2192.79817","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"14","positionMil":"1401.63859,652.79597","isAnchorPin":false,"label":""},{"uniquePinIdString":"15","positionMil":"1712.74971,512.79597","isAnchorPin":false,"label":""}],"pinType":"wired"},"properties":[]},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"TEMP","category":["User Defined"],"id":"6500d8ea-11fe-42e2-8a9f-99be354012a7","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"49baae61-cb81-429b-96a1-6cfb8f124b59.png","iconPic":"9c69fbd4-c376-47ca-8b4c-793dd402431a.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"15.00000","numDisplayRows":"15.00000","pins":[{"uniquePinIdString":"0","positionMil":"45.31000,541.03000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"111.62000,489.31000","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"228.98000,493.29000","isAnchorPin":false,"label":"A0"}],"pinType":"wired"},"properties":[]},{"subtypeName":"PH","category":["User Defined"],"id":"8e0ee0b2-778d-4065-bf79-38edea29856f","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"256658b1-ffe9-46c3-9f0b-70052a8fe00d.png","iconPic":"d18021d8-4522-4af4-a3c6-358ee97fa8ad.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"18.00000","numDisplayRows":"15.00000","pins":[{"uniquePinIdString":"0","positionMil":"415.56444,426.59333","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"479.26444,379.41333","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"547.67444,341.66333","isAnchorPin":false,"label":"A1"}],"pinType":"wired"},"properties":[]},{"subtypeName":"TURBI","category":["User Defined"],"id":"6d0c07c0-db0e-4413-b9a4-ee378c2ed587","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"a1588c66-a70c-44df-b30c-55fdbd854069.png","iconPic":"2dd92824-eee5-446a-82e5-cb3be823b6e8.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"18.00000","numDisplayRows":"15.00000","pins":[{"uniquePinIdString":"0","positionMil":"27.90000,414.20000","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"69.55000,337.31000","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"2","positionMil":"124.01000,268.43000","isAnchorPin":false,"label":"VCC"}],"pinType":"wired"},"properties":[]},{"subtypeName":"TDS","category":["User Defined"],"id":"1cec4e8a-72c2-4b6a-9a5c-b6be0dc427d1","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"a05d3615-68b8-4f26-98d6-1aedf7f6d878.png","iconPic":"b75f5fea-d559-4623-b1ce-f8cd504066c2.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"18.00000","numDisplayRows":"15.00000","pins":[{"uniquePinIdString":"0","positionMil":"974.02000,426.69000","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"1030.68000,479.54000","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"2","positionMil":"1088.97000,531.29000","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"}]}PK
     eO�Z               images/PK
     eO�Z~`�	� � /   images/5de4bec6-ccea-4571-acb8-2cf876e4e4fc.png�PNG

   IHDR  �  �   ��ߊ   	pHYs  �  ��+  ��IDATx��Y�eYv��t�cF�YY�U�n6�f7��d�(�Oz4��`��C�l�aЄ'X���X ͦD�챆�#c���p&߷��Uݴ!����Ug߈g���ک|�=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC���=     `z@@@@@� 0􀀀���-@`�[���� ��lC����`z]ב�O2��V�������}��=�m��+��~���˝���������o���G��m#�v#k�n�]��3�ɿ�5���mھ���=3+����)������,��<������gV����]S�9�v�_��Hr�7�/�/�sM��{x���t�������*J&�8n/�(��Լ7I6���޲�ˁ���}dwO�(��q2�߆�m�|�ź��:N�i\w*=�;7[�qd=ߗh����2^G]|�g��j�E�U���<�w�[���8�몮ʤ��Y�����*�,N,��$F����NZQYV%�L��Q\�j@��4K��*�R,�o����o�%��|meY�E�{s�s\Vi������f�ygY���hf\��c��ŵݤhg�"�c��(��t��)����5v	7
�U�βƣ��B�J��%~Ϫ:^��2-E�i��N��u�MV�1�hK�W�y���E��m(�*�{���2����V�΋2��u���E�<Zs�W+K��2�J���*3tQ�7����=?�s�k�Sbɵ��~����n]���\�����놛q�,�r5�6k
C�����:<ďE��hT�d������gs��9�t0����������_���������7iY���_��l�P[b$C���d����\��� ]VVQ�o�H�-���_��S�	fZcg�ׄ
�/����ci`��� =�Q�����{˲\�O�u�&�nU����^%`�����|w��n���}pD��oq�4�����6����UT��q������uVTU����9��B�pmU��gQ�GQ�GỈ.�(p<�UE��q�wF`e��+�	����V�5�eDRakp*�(ɋl\��}5YF���U�%g�������%�wɑ�p�W��H��~�bs��Gk|�c�Б2"���ȑ"7��ID��G�U��Yml�e��:�)�EF	N��c��w^��dIxR���Q^CD �A�1�8�2(f���pk�$45㌢Oe�1l�e)����X+�]��rt9���z���Ǌs��	W�f1�G%f ��*��qZF�~a�Sދ�p4�Z�	�0#���D$D|�F�DGyG�I���a�Bf~Q�!��h�qH88�1�o��G�ɖ��un.��$Kke��Qsh"K��1������2�؆���*����&����/w�`���[y}nX��o�H�@���p-�\�X2	��M�?��� �@�NkQ�Z-¡mZeY�/!�dI�m�^�9"u�4V%�8��/1>	��l�l!b@6�(�q�T��os�{�d�J��V,�(�$h����_� ,u��Ȯ�?x]�$V�i	)��k�����C��(s����>J�,[Y��J�z�%�RL�c�����5�L�T
Q��[����Z� )0m�r���U�S�՝��T�
k~n{:d	H�&��yL��V��fw�����c�� J5mh빼���<�f���mh�ժh��>�x�X���`����o���g����'�6=;�
4ͻt��J���E�j�"l>#��%��.��j�E���U���`�_'")��/J~���։����h���&�;�fj��27lt�WR4("d$��`�Ge��ව������\��U���\G�	6K�����N�;ꮿP���I��u�HP�Yfd�/�3�
��#�.�}�����h)	sB�G��>j�o>#Ǌk�݆�T�-�n������X��)�ѕ�=��1r�e]@�ʩ��l�����Bm��m�z�vI����k���t� ����b�Y/%��ث��X��+�W9R���IڐBJK�R8���<ܤGe����5�gkI�{��t�W$��k�p￳>��'syp&�������"'h����_zN�݀~�����OR��7�b_��Dw���s�;�tƈ�:�H�N
J}[�7v�i_R�����7�;�+��o�^c�Sʃ�׷���|�l~���ڃg��{�;ƃ���\�l���r��4�>��e=�+��������N��]^z���o�痃QiG�x�/�{�B	J�ݠ����׆>�f_����
7��c.Y:5��c�t�(����tgh�����	l��"�ȭj�qB�E�4�6��|�ȋ�T�☺�WJ��uDa��k�~����Zu|�&~S3�5����F��"M��r�0�����4��oή�4�/��� z1��[^�?����޿�l=O[�S94c�R��:�16�AA&��s1�;Ē����ye�5���$R<�!l�"�?��em��W�n��cq�����qK�<��/���+�.3ob��]bz�h�F粯��,s��;��:����^��>�R��{^W�Ҋ5�vx.{��9]*2h�-ʻ���͜l$����d�:rJڦ�%���+݉]w#��s��V�z��u�C�P ������tC�Վ�'"�k�vp�gi��yf_gӑMFSa�eh��!�	�̉��}��1��-�S�C+r0�B�BG��u,�2��͜��M���Zkȭ�Z*{� P�ǤYwD7�b�_
0�n�w��խ��5GG��K��+cm^��������	���_�sQ�a�4��Z�K�&2��������JSP�����������b[`N�|jղ��|�y^Y��	R��#�4Ͻ^O�k��-�oW����!���Jj��o��!ښ��/��l�y�-\ӌ#����ꯍKu��7��<rU�Xe�j�ى����|�5��9�B�����h-�ѝ��̜ �A�II�gMÇ��m����ӛ������ғ�I)�LO�z�}��=	n~��ߣ����KM�=׉�n����4�����G������<����?���ֹm1>�CDoUyթ8E�|���AThO+����%������~�j����H�
��i�hȔ�f���R��vv-����늁C6���.��j��%�I���Y�89�nN>�D�\���j�Zyӎ�l�]��|��>5���Z�K�ی��P��{���ց��4���ﶯ����j����Z������j���7�B�f#�|���$
|��=k��Xww��4r0�
D����n,ü�������M�`��Y����8�ˑ�����i��Q�Y�J���p��gG�AFX�%�uqve�re��J9��QL��Rg����'�4'�&��E��Yf���Bw:Ƃ��gK[�s�4��A�_[+��0��}�1��;_"�������"�(��j��J}�%}����'�����w�n��oa�sk؁�[{5��df���3C_��9�{&�>���t�?��@�9��]�h4q^��>iJ�1hC ������]	��nF6�ϱ�\��}I��_�x�Z��GYØ���Uk�.6�k�Ŀ���)�u�a�w�T#L����|���+m�{0��.���)����e��wZw��%������w�oZ_#0t�e�.�@t��[�jE��}��߻<y�_�G����G?��~�wF��� zR��1�%�$i81vM�Zښ�g��L��*��3q�:	;��U�Y�_��I�U��6�cxe!�3�M|�#Ɲ�=��7�(�������*����ܖk�|�0�
Ĵ�Y��a^�ZDRҼ�Lv�ʤ)&�M�l0�@���)zF�u���x/��2c��ج��|wg�Vb�^�z{|��P+1�R׃c"_<��:Fr����!m������C̷#1�uHc��uFL3���E
_�e��-'aF�`��,�5eZ�m��y�cshy�#�
�[�b��(ֺ���ز=��7T[g鍍��-�%�dFO�h�P�a;u�/-"�c�/�o�`�͙���2'j�,7��|����<9�l^lƾv�b��%�+���0���g�٢[G���s���,�Ӵ���h|fk��F�󄼄��n�%�蹒<w�
��PUN��d1pAII37רcJZ�_���ո&u���j������`��L{ K�6hu!��`�,�m�>�|MmM��W�����f�G��Z������1@B��f�S��~oS#Wcb�#̜u!|u���]�N�Bb3k٤H��*׉���ҹH����g�\��k�s3u�2i�9���etv���o� W�
�|��w�PY���_mݫ$dі�@�n$e��|�{�����CۅS�[ׄgش<U�he_��5�@�;��j�Ʒ.5�NXĺ���ʖ�0�s1�Ͽ���-�����ɛ�/��g��{W��� :�j�|Y��%9�K-�������\�+h]��+]��*����F"�qu�a\�w%XǬhr���O�������9��2f��0�X��l�:/ܵq�o�tj�#�ə~�:���Em�ӃƷ��9������Ƨ�O��.o��6ح�1vfZiU�4���7��9�̡��1++.P^���ȃ�J��w��CF�J�%C&���ID	m1����̶��ܢ�}N��ms\O풌����I��jL�NZq�r�s	��̊����V_4`΅�~V���k2�ؙ���bd�lK�b�L�4�`��h'Y3��&s&1���6���` k0�*i{���t��2i�
}���,��.���۬嗍�����}�d�c�Y�!�x6��`g�ڝ���{Ώ�J�pn$�\p�ƪ��g]h�\��,M�cY�bZ��7�*������e4�dp�5�sz�R����1
�l�z>�b�5�j�|^MS;>�̭!iNnq-�Z՝�s]�4�R��>����h|Wh����V�9X��Lp��%��6�O+�e[��bO�
ӊ����[��y��p�
���PW`ӂ¹��B�ᨼ�G�<0�\�=_��KF��YKF��c�NP���`��SYB<���5��;}�Υ��m3Z�n�'^�0�i�/t��h�Xru�ԝ��	R_q�m,c�\�Υ�9�^m])��6ŷ��ҋ�YW����+�(x�_��ƨ�Цڻ�.����\O���)����sv�Fx��/����ڵ���c�/��s<k�G��yE�aVۏ_����|����2|��WQ�m1�p�M�����Ą�ׅ-�ŗ$��{�p�n�E�g]���&J~��J���(��ݿ�n���6��HĀ� !�#I���Y͗k�5(��Ys�f�Tm���"�Y�]g�����l����������8������Eq��GTyo\;���C��-���NFv�A����d$�3�iKUN+���GD��b��F����G�#���H�	�����g��!�:��9 �ZLR�1ww�O��p b������W�J�U�KY8�%�����,�6��1�ěy�G�@�V��Z���_�~�8�z�����*�7�\-ў�_`}��&0�P�p�Ӣ�E.�$K]x����	5�N�ָFA�Q������֕c��n 1]A��f���O-�^�?1��#'Rfq��.\@�,�r�"\�,��}N�ؖ�A��g�����M˺}�����ʋk�1�mZ
��|�zM�`l��<}f��=;~s�wb��q�j;D�3�Q�ҨI So���e�¾��^�G{�v���\$��tf�/^��f��3H�r���-�(�@SB;�`��c5�6:>�+��@2�cn�v+� �d;{�k�Z���=6���t��h��ݧ�a�B!��
RC[�dT0�  ;�ش:m�G(��bB�L֋�ތz;��d�(0.u1Xc�g��{�>�`�k��k��hkY>�g�r��X�y�:�)��8rq`#M� �F�r<w����
�\��)`�����te���e&:Ba��`]���^>��}��s5���b�xg�}"�8�ݣ{��V���L ���E��K	�-�m�7�I�,����;�s9�r��Z��ӖF��%����0��,�>�t�&j����q"�ʻq�;����}hCo��"�}�Z�(_~��j��ո��O��>�����m>��Z�7��'�S)rlV�n�5M�0���9�\6&'�l�*��HR2�:��+�Q�d�q��1o;	���~egŎ���,���h5�^i��Xc���,��)U��ֹw(�/`���X2�FN��%Aȫ�G�9SS�M�f�2���zM������4'�D��8F��m�1��"L���0�F5C����� �4�rV�WV�H.���6�0в��ڬ��Z�`��;Cmz�c�{��H��v�M�d�`�=#�c�k�I��G&�.��T�hc*��k�,�e�%�ȥ�f{Z��c1J9s�9�a��1��.W�-N)C�32��Ddr�X;�-Bx	!��(����
�:�q¸\-)�:a,v�щN�Ka���3I������h4%G$����\���+��rB>�=�5��e�6��Iǹ"<3�``�Qoh�z<�Zyu�y��IF-m�pr�EG�{-#����|B�>Z�fj�)���lrqcק�x�<#�ю}���ka��}���ͮ�-�S����#\ _�{�������)�z��ZY�X������B�v�i�a��\n�L��ܝH@��3&#���
�{����8Z��z�0ދH���t-�F<�	܅�ɂŶ,�N��Ǡ�t޹�Mfpq�E� �٥�AXD(���ņ�n,�4�]0^�h<I��� Je��w��:`�٠�qe,B뫗%69��m��غ��]��h�`hu�֏������f㉻kdN����*q	�6�EO����C�k�;�;����eb���c\"��V�%�%~�`ҝ�PBa��˵��H���>)%(R[/b��:Z�c��?��l��?����V�%� :����J"@�h.�9'��K���H_��&-po��4,�7ї�Ҋ̜V������}���5LZ���̦4���'��gS��W�r.��K�Yב
D�+E�q/7O%	4q���7f��w���1��d�8���K{-�k�L^�7E½��	�{��#5
0t�����dl3h�9��@��H�����CC)֥��������lM��1�pL��1�D%7�"�i��6ΰ�͛�_��C�:$�ܜԐ�[�o��W	-�63�f��%�&!��K<+�`��]��s �$hg�;�|�1� �q$���26��iE!s����Z/l2Z�N`3�l��9Ybި�E ��cS[�[s�z�,���g#�R�iivoy�f�~�î������L�-#�.
��X����^�om�/����Khk��{�8��2�}�E������&�#��1䒉Mg�+�Z̅c\�Nۡ�#-.r1$+�&���Jn=33`�ZY�-U�g��ι���C�Kia���5��te��h!�v��4G�iϭC%q�7�L���.5�vO�7C��C&^�Y%���9k�2��Q���>�U�k�*d��oG�e��������¥��q߂�8��8���>�SZhW���4�C����^3E:m�*�SbϤHgR'��1�
Z�ڕ8S7:@&�x��g�u� �w
X�c���[3�۩^p��ՌqTl\,y���2��&%��ޥ�5��݁�uφ�l>�6ƹ���vyz��G��?8ܷ��l1�N��6OnF
8�;<�A�o��6]��{�$�6*E�p-�U6j�X�A��F6���ȜY�.�\����~������`�s�ɣ��;{f��	�L
�
pq�?v"���WW�X���r��'�����~�/����m�a0��HY����"v�	���2=�4w�
H�O������J����o���z)O<u~b�sԵg��wT�K^,E��GL}�8}�W7�X�"��m&.W3eP\[Z���롩�Q���h��F	"��.�Sԕ�p�ZЋ���HQ_�����t&��G.jj,G�@!b��.��)��L�iq,�ڬ8"�e��E��{]l��%��Y��7F�V`����(��M�� ���� ve�k+h��bj+��}I@����1��S!q#�aD�+�[3Y��&�4���!�X������B�ŒL�L���k;�h�V˥���I B����eC�rG;'T�3g�c.sh�m:0�L)q��5Q)gN�K./�;���g4cb�~2�EI?~�����fq}�Yx~[
��R�	���/��z��t-W��2Z0~�,�K��9����<>�mR4j�U�̐B���:��kGV]n;	�s�H��'�o��n\�=ص��+;� w:����ۤ|�H�Npka=�h�����=<��S����C��Ө�V�����,�`�� �
 d1+ZhG�[\�*($em��`cM��)����+𹖹�t)QJ(��L���^XA���"�Z��-�Œ!���%��̊@ۖ�J�"�˯v3�-Ҁ�p����s>���&Sg��j��. �ׁ�LWS��q���̰�ia��,*\��Kוe�p)��P.��c.#�6���7)1�S S��%�-�w�x=�8A���<�3��^G,"(K�b1��ݲ�#�w�����Wk�@V0���S6i�>H�v�կ>�r&�,�J�lu�a��'���v��g<�//�w	btY�!X�ҏJ=`N3/*Ч^L������_���i��������*�&I{�H��w���Q�B@>���%���󩐐���<L�
6'x,�YfS����U$��mV��ܼ&�EDA���A;
�i����ܦ��^�qڌ#��h�B�O�,��᪘93!�
<2���a���0��4K�ў	�_<���v��͕e�V�i5�y>�UfCINڕ�jb�oV�#FsǷ�X|"�>A���ۂ<VИF�Ii
_�m��\�`�?zhG���b#-�/�b������ڢPұaGq+H�g�)$�����l�6GKF���ް��NE(z ,d���M'�f+@�Ɖ�^ѴW�J#˺mi�ǘ)��1�?��u�;ҘV�����=5Q�:�F_MF6��,�v���q�0��c�o�F��mQ���A�GBz��5F(���n��ks|?�0���&�3_3 ?��.  Dp������fٶ�B�ɊAei��)^C��¸q=P����N\ ���z>���m-hN@��v$h�CC��!<1���*`�z
��L�s�|0~�t`%����]~5ޝq���J>T���J)�AF,���XL ���|:��7�]^\���)�na%Qp���!�UJb$:�Ay������.خ�}�АS�����%0�l�������ʎ���X�s��,��o�%�LW�{�|)_�4ȳ�[�=��P��z!����&��"� �$�_co�Ʃ��ދd�ZS�ZǶ[��`L֎`�@�f=[���Xy�&+MS�b�l�@L��i�1X\���fAg.!���&z
"��1��ᮬBtw�X����\:뜹��Z����m��}�]xMJXe�@Q��}: �F�˦`��I�}A���?�+s���%�C7WZ�$���8��C���|�_
O2��^V��',*�)�e���R��y�����+{	Ӓc�� �5���,a	�Z����끆@�:�
I�]�A���]ͧ������`�����E���Q����;�Ï����9�ӓ��?|���y���� :E�څ�_\$�_cs �]l�4�`��d�f�}�m�M����W�-���@1oF�BM���H����#A���o�1�٥]D9C�%$ �u��u
�U����c<2�M�#O�?������}�;Ǧ$��д_���1��m6�K��7��֔o�*�Lw��[��E"g^�d=����l��-�c;�Ь�`���}��?�vN5���xl#0$
&O!3����=��TE�'������7��)�X��#64��n���F� ���C������^���z{����1� ��O{�����vE�7���}��_�%4�Z>rl`�1'~������X�1 ��>}f�'`B�ҳ4���Z�;h�l3��`�q�W���x�b4��̑D"n��B�~K>ƾ�ܻ�O
n��Ɨ��ُ�Os��Ԟg���\9�; �����M�av5�����K���-�E-k���m�!��@����*-�͔/\Ϲ"�c-���=�g����N$4�v}|&!�]�2#��JC��+�qi6�<x��v>�9���_�0Y
G��3��{ᆦxܻ�Z��noGA���/��ލ ^]�)VJٜC�� �A��B�	]j��?��o_��ɉ�� sXb>*|']1��>���0����v�yss%����������:���\w! t <�D�	o<���P�3��Z���5��V���	�ﯯ�jt��}�F4T��YU� m^aO�clt�6�F�}����^�����T�L>�7������zb��,�v�k)�r�^+Q�/��4z�	j���9�t]$�*�`^�ij���(�x9�xB��t�g����V�?!�Qȹ��������K3ƴ�95�k����y�	�#5"vY:�ײȿ�g���w�J��}��W@4�'Or�X*�x�	�J������>}H�p���jd�켤Ń4{��J�X%�����ӧ�ǧ�hK�3��qa�?�����$�'x��>|���Y���Mzs1S��0��Bf�h)�AZ�Y�ڤ�Hc!m�z�1[�oY*��n��ȧ�H#f�j�ģ�BX���:�yc� z�� >#h�K.h| Fq��-@�� H��P��]�����=1�
��em����V��a>o�g��8L�xcR����2�]�k�G��Uw�O|��w{�Y'��/���i��	��T~��xjo޼Q45	��ё�Q�Jh����{�yx��}�߰��3�@�y�I0�jggφ;=���A�J採=�'O�ѣGV̠񽿶h$���%�Nh+�>��M@ti��E&ō�����ޜ�i1��\�c������́�j¼��=��#' b\޼zk�"�~w�������	���}����o۫/��W�x���������>�����Ey����1����`0�ch����'��p�0���L�G�G�?�4�>�/l>���͵(-0䝽!��T��\#}V���=Ě��?�׶�A۬r	.S�h�v�-�kG���|b{ �G�l}�v��O~����i�*΂�Zu�eu�B
���GŔ��Ԛ��v�gE�Ȝ��H��c������f����Z3��~��|�S���m�=8T����!��&c1N�ݧ�mP�0��gpyx�BVng�+�0���vro��d`E��Nfx�,�<�Z�Ogv3���D��CZ�Z��|����iu��J!�?ܓ0~>��	4��B]m #b��c�t+��h_�i$פ��{"A�p�L����E!ve��.6���~�������N��-���|�>-rg-�kyکc%���7a?�&�9�:��ŉ|�,��l���KX]�s�> p=�%v����&��rf,�y��!��]'���3U�Iq����$5u(��h���+֮<rS)����)��.�C!�,"�ݼ�!���������л�|����J�ӂ����(��s�xV�\c�!���/K�I4����|��Z/o���W��,Tp�ш}tw��;�k�և��*��|?^9���A��T�]��+�ʒ*�p��C��WN�/�{�Lj�\��\�~J����];x�Ć���A���������]C�L��B�2��H����� l�sŋ�L���U2}�jo�r��ҙ��>����M�UT�:�{�����F��ݣ�H�(�����㏞�?���o�����gOۣǏ�}d�˹L�W�i�� R���Si��剽��j�82_�hpO��&v���&ѫ+��G�|�?j��a���˄��mB�>ƓAt��`~W"П>}b{����tm�\�U���wBx*À�񜝾�������M1t����5�����N�V
h�CjKs���u,m��C���O�����N�xX�>�������t���ؘ����3;�}�)����W �;Sڅ�Ϡ$�r�����.0���?���/�E���b���������jn�8A����O>�o������,#|F�*���Ď�W׸g1����{2z{���|�J�r�b,(�0�re�&������؎gϞ�0f6v�%ȴ�;��|i˛�������y��	�h
���G�����~ޛ�k���H�s[^�@��h-��Gm f��J0��/���]���Zb	�̜�k��>���8����E�o�K �����zj3_9p@�`_���n��s:99���+0��=z�h�{�����������G��v�<�\�Bƺ4�Ҧ����{�{���zLnƶ��`��}Ŵ�u��h�V�I
��eG���k(�d�&��MW��m���D�:u��_0�p��0igr��؏�܌!�dfLs9�θ���`8��e�\f� ��5�{�c�t7Ơ�}���mRB�"�`�i�*����%|i����M&�����M��7�{��bRYhKsJ�BV��!�|j��;ߑ���ٙ�
�_��1s�����cF>���Xs�.������Ǥ�V���Й=�S���jd��Wb�������4�mL0}�y�f�F�&���op5�]^:)�c�����yf�:[9��mnQ�g��+�s���wJ�rF_;}p+0��v�L�:}Y�/�>4i<���韚Bs��O|Н|{J�s����{_ܝ9��O����S$�J�*�����.�7��6����٩]^�������;�{�;��)��#0(������R��ͮ/m~�Rя�g���=�s|�>_+O���>ܫ�w���� x���}yv��L�UL�CsQ�gY]�)�ܝ�����&�w`⌮o�R�ܱ�_��g'!��h�����]Ca RM���-�=��m<�I��a����xG�=�A(FV�}�����~��wEK���@h��..����]����ۗ_��o�> ���u���~�y��g9}�7[�q-����v�q�{��޼?��mX7s��!4�1O���͵�����p��~����`,�����u��8���S[CȰ�_v:�����6h�y��1���]�g}0tI�+�;���Ax"H�}j��4Cf�𹭴g�~���;o~�+���y
-{ъTk���S��L
O�=����짟Y�0�s�CN+DL�n�Ƭ���0w�gǵB!��r�*ɬ������H��K�����!�W���/_J!xwz"M��\{G�fB]OD}=�m��ٓ������_ڋ/�c�Aȥɺ&�Aww���	�}��{@�BpyF���3����bd3��>�XwU��f$|�j���?�m���9�����3�B;��)D� tн��?�ߧ�=ܵ���VB@]͗
2�[�Ѧ؄cH�-'<�"�:���v�g�]�כ,��b�R��R�Ě��6`X.JwHL���mwvD����%)0���Щ�+��-������w�H��K�r�RP�`��+s�H8z��HbÃ�<�pr��c��e���6=��К6h��b:�5(0ELwNU���Y���f�-����[��C�DMnF��tƜO�Y$I��$H_�!���w�������*j*.��j�M)T�����I1�΅"�N�� "0����h�gәM1���+�����'!��]��s�h��4�Tʐ�c��[�զ��G��jT�R�\:��OhE��ðK�_K���_��2 �b�2�ܨ=j#�����K�2�N�3�+�p�]�~yi#���"��B����<�@C~i� �dlLšF1������2�����vD-��Z�v��17]����=��蚵w/_K���Wf@
'R�V0�g����Z.���1~1�.���LD�s�d�3M�������5�uac���$g��l|}#��6��e���777v	�9v��;'����?�&��;��(�� ��)�����X�����χV�v%<DJ˔Z����1�||y1Q[uXl�"�ch�\3<\F�`�Q�׋���f��7�jO�n���O�����`���\m<��Q}��xbK�S��v�u��|�Mkl�G���}��=��'��\�[����.���G��l�5s������=~h�����!��;�����Ԯ7-���j^�O�e��y����ѡ��翰���_�Y�������z��\#��W/^�!�������m���wo$@?�0t�dZ�)���T�j��?�����i���3���x[0�Ku��9���=��oߞ�݀��O��&})����Gr�M.��a?P���o��~��ڿ�˟������a��B@9�ٳ9���w������o���׿mX�o~���}�Z@i�J�(8v?��:��dX�?��>�Ȟ<{��߅�4��_�s)C�3��ڔuS6u��I\Le�.и�ժ��u�`�p��q���E��b9��U�,��Cd�*�q�}�$]��:�Y.�:c�"�s]fJ����LI&a��L��;�-���;L�d:&�����e�se:M�&�����!aF4���Ꝫi�/J�*e������K�*��X��+CO��G���D����&�����sI�~a�M���1��B=�(�w�(K<{��5��`
��F���n��xЄ�Q�d&ֺN�U*z�)�Ԙ�ն���6M�$�L}+]������3��P�RK]����H�f��M��v�Z3�n�W4��ѯt�rK��'�qS�o�
R)S�������y�4�b��I��q�r#�'7�������k0�9����Y�Q����T2D�Q�c5J��
5M`#5'1��Zؼtg�nh�/�Yˢ� ��oT��"���'�^��+���^B0�U$�:L�b����i��|քKg�e���M�+�F]̽��+�Ly��9r(�k�u�2�F�[s*���`����+�<��j��.�E�N!󳗹�(U	�X��a@�[��\�7���8�2����}�?ܷ��iٕ6�k�������h����R��ЙLB����-0�}����%���zn��.����Q���޾�1�q�����hߧ��BS|�u��<����=��)N�����?S��d�gϟ?����e�BؚڟN�Fe�L��g��L�Gvvrlo������������%��˛k	r<A� }_@�>��xʀ?.6����l�aߎ��)����Ah;�X���K;}�Z���|����e�n_Lx�uryy���*Vfk�ݛ�b�o��
���ۿa�������i�<,������L�
���'ϞZ�;}���	��s��0�/��!Ed��b}J���a���,L	�:
��:�g��Uǋӎ�MU�&�=�7�0v���Ӆ#�tT�HnNӋ]>����Է[:�h$�Gs�T��z�;h	��y�R����۠.�t��L�kC��v8��.?_��Aw� �3fs����F���$�1UUQ.oշC�T}�q׍��,���1S4䓩��=�|D���J�E.5Fğ�g�r�E%�6�� f��.�b�VW��n���b+�/._=�Y��0�VcƗ�K$����.��"CU�J�I>���_/@��Q����j�?+W�d�$2� 3(]�J�\��M�LOa�;{yy��`V�5�h���Y�|���#㩫����=G����G�p���Z�@�}"���[h�NW��N//E��=~�ח��Æ��d��~s�N����"���-tAp�̓�}���L��>zb������q0���qq%�lw8�O��6Nmo�@�eT��ō�����q��݀@R�><z�qcճ�{���v|rf''������<��U�:9� �~������2��(�?����5y���s0�1��^7�� Lf�Pa�!�����x��4�c���-S� s�Kg��0�����w�ЧV߾�ʶ̘��ʉ�ㅈc 胞�d��1=�g��x�J}oG��|�dW�ҵ<�d�����&
(�㻿|�Z��1K�Q����sV*G�r��x�J���.�z�-/
뵰߽��=��a0l��z�+K���s����ͅ�?5,A��+����q��̶-F�f1��)i=���ZF7�b�d��]b/^X+�A)�=qic�L�Z`<���9���v6�5��+����B�ꃃ��@+��S)LI[*�uj�X���W�;�-SNy&�I%���0r�zT0�ÆX/��ǟA�-��gV����zq=�������V�.�>
�ҙ�e a]�V�P�"VQ$](=�%M�?�`,B$zĽ$7 ����#�n���z~Dsy��������t�PF�-T���.MXTݞ�ќd���(}~�X�t�B�{������Ԣ�y���dY���k���.���.*X6xA��w�X�q���f) ��_��w�
*UuQ�����M#��q­�yS��|��W������D�ƹ��u�/p@FW����:5n>@�b�Ǒ���h�/�)_�j5�R7a�ƞ����c�|�B�=l��[X�"3W�$�Ff8	˰�ͥ��,���׬��v0�iI4���p?5]2
*��$]S[����QZ����K[����}�]�I��Ϡ��L���
?�%����ƛp/�|��>P��Rh����?sL�p�5p<����և:��GP.�3�ay�)���T�㹘>��l�,���Q�����F���|���n&��L�^�^��9�<x�L��8x��Ώ���\�ߖx���ȸF�r��GѤ{y#a�Tu97S+Z�|��}�[ߑ@���2*���矿Ҙ�mv���xA����AS�淿+�A�L�@�Ͽ��gb�����z W�������?�J]�F���c{	዁]\�,�I�}������u�
W��4!_���7oe=�d�����R����٣?Q��h�ʘ�K��g����xd貲Y���l.��P�Dn
W��}r��,���9f \�댳�5q/����jvLc��|�uvuu#����;Ͼ��x�;���;Ը��Ѥ?�.�>t	��7�G8>��H�
=��k����W׮�+�3�-!D���}g��篷@C��!� �WGz�
c��|]K aU�����̰��W/T$e�X��M-r��b�%���D� G�q��Xx��x$�[�18:Mљ��$����)m�����qԢ�[.����g�@p�b]v:�O�9��tb�4�����.X��iӾB���p���-����X�g�� ���+���v�-��N�0��P{+���Y^��:�B4��1���I�R�h�b����������נt.�y�;<�T<խg�C���iW�V�۵�X�]�JTH�����*)0,r%�����ޓJR|T��S�%CgZ�"*���eK�l�:�ԟ>ŨZ���h��K���bQ���ƺC,j��\���@p�f��N��������<���fӸ���JeN���c0���T��kX��07ͬ�̓�hC�N"1c��DL����M-�0#!r�+�NP03ރi��A'S49w��ň)@���	ejXtoЪ@�������Ѝǌ.dF�����Rn��YN��1�V�!�y�;�Q��Q�"�ASd����(x�
�"��O�#3����̓NV9���a��t��� �������ҹ0�yb���/^�X��w6w"�}	����7���h�P���ˑ�	�������[�W�`ǂ)&t�&����<=?���s�_���DK0��̤�i� 2�VV+��K�^�t.5zVSc�?�d1����&����ť�?;����}�<��t,fɲ�=�OR�=�1N1�J�j�Zv��ӧ�Ʊv0o=j�,����9ƍ�ɘ�^8������'�:t�#�|��,���9%2o�7׶���������G�ʇ�����'V@����g��k���X��Ќ��_����3�y����������Z�|*a�Š�!��0ۏ�l�`�Lc��p�_@h`:'&Z�Y㾫셷��moБ5��'��`���{
bN���{��X1�Z!���N���g�B��GO�e����^�~�y��a>h�6���w���o�*�˜}fR,1/ǧ'X;gb���V�5����a��ҝH�9%�,�g�Y�������hy��
��s��¶1O����r�L��}�R`K����:�-r��gF���:w�U]��/���v}�P]�G�HU�e$:�$�}�MX�k�\��3��ED!�n�.��"cA�Ц,y�f��sѥ)ݶ��:���/� �A0����
�¥5l�Ģ�#�
E������;���S��N2$s��K��:1�3�F�t'��������J]&rr*�S�̟������cW��a��?�n8I�0J_�V�`��@G�*N��f���@Zg.3���`��rly�Y��w�RXw|M��l*sh�C���1�ɵ4%�zh�؁T����OIf�Q�+0�+��rg?�	�
B3['�:S������*�<�� ��9�4?Z�N��{Sj٬g�vG*��͡(o@�I?}������IxqK��i�q����z2�A7C�����4%���`�JL�Z	5����u��S�����UJzW��1��6����Sj�蜲�	ƎD��ĴC�wR{�/�1G={;ǐ�]W)+v�~�#p��"0��l�
X:Xd��X�▴'�:LU
u
�~��g �S�*W8������y�xƘ&eh���E��5Chf�0܀�P#�&�Z�}�qF��;%���`B� ���wМ'':CW�h2��eG���gN���	� 5e�-`�zy��Flt��;`Ƒ����)�?���v |�}�wbgt�7f+��g���0�O�}�r�9~�a_U��'7����I��])�Јk-�Th��<}����i&��]�;�w`�
�<q�qa&�|���;�-�C�X��'��i�m�#t�0^�l��.\���+_;5v�����|��.oF*��������sl-�	
8?Q�Yw��X'b����Q�,	�.d^wu��y칯9��-�Ղ�
YJ�,q��O���E˫�d�Φ�@���dt��9r
G��E��Q�t#N�d�Y-E����/3V����}Ё��J��C�_�]T��i��ڌ���Es�ß�S� ��zz#e������C��S��ueM��e�Zh�ry隔��Q��t�P��O��T��VO���M54@���������}.-����u���-b�D_���Xb��/7�Ӹ��9� ��Pj�4k�6�\JZhv��zOy�c�xrV���5�^��w�|v�DK37S�Hp'�N����@g�*�J��·O�SĜ]Vy���
�|��s���%��h:�v��h�Nu:�3�s�]�ەEsw�9k�����*g��S����g]:+
KT�����=YOfR��|W4�Ai�5��g��ĞX3W��țice�W��X�����V|������w���F�v���srpp�P Qcѡ��`�@;S��F�i�� *�%2u2wV�KEr
�f�A�Oe*d�Q��ie�D��b1�8u���ҤKr=9��b�C�K�f~MR��o���Z�b�N�����3[����<�D&�D�aa�U�`���e�b�8ا����.�6�@hC�;_��ԥGR�� �S+� xq~%���n_#��5��/�F�����MW�d��u9���(�*�C���D���o�!�������oU��>9������	��Ϯ'69�����:��r�Q;���5�t@H����d�r��d>[��'���ѻ���chλ�E���3{����
�=�e��ٳ��-0��Á��6;��Ѹ�y{��bx@w�|�h�h4�������?�=� P`�OW�c1c�V�cJ+-qM��֥�p8ZV(ն������\k�͚�d�
�0��:-�k�����J���i��~4���W���+��w1͔k�.�66�R�����b0��ťhS[��no��	y��(��T�@�i?���%b6m���7�1���b��@��nɥ�bd���gy�<y���Щ�sh��i]ywT܎l�c壓���S�o55�Y�]9`���ʗK��c�/�~2�E�t�<
���� 	�e�NprEe���!��ߎ�F�>�̝�_�#���E�� �'�@d.����t6�RAH�er�:�;�ɼ�G�7k�VbI�<ɉc3����;5��Jér�Ѡ-��2Ϣ��Ny{KGjZ��Ln��ѩ�r������l)�<qG_��6�@kZ�6���h��@�1O}���^E�H��|k����H���1�>�����*��T>V�B���,J'd�<�ѡ.
[J�c|D,�����.�B��i���$�-/�iYq0M�yH��w���@�����Χ汕�#�K��H`h�e:��I#i�7h	b��jYǲ����l�� s��Us4n�-M|�[�v�� ����.oA�wQ�r�B�������A���\��ȑ�3��d�/��45�1�Y}}cS������Ӭ��7���J��ܟ,��Ot�Z�^l+��\`�x�jfԸ�9�4�W4}O�Z{��Z��b?�"�>��2,���Ź�W��ZieV����y"(뵻P�Yڱ�1�k��[�t�0�
	OG���G�b�n��H�����F�|�|��U
u.��,tq�-51��DEe.���닚��QKϡkM��r���[���b��UU#ܷ���@���Ǩ��Xd2�W3	|��3���,�[�Sg��ks.+
w5Q������O���W�k��=�G?�[�y���/,E���'c&V�޼zc�{��!��|�u�:������}�V��:���3۩���]L����M((Ѕҳ��cO�>QFM�ە���tf�r�J,A�(�V���}���m�^QyQI^��g��cLrUmy����j��ZX����k��A0t0.(�L]+�����^�v��[׮T M�$α?��E��Δ��q�4���R�e�����Z�DX�U�l��\4[�Zɏ���Z���t���D*��V�7���YljW�gW��X&�اsЄ�v�T0jb�D�7�����ә��s�#f����6N62���|:�����VZ^&�K!�.e6 q�ݓv2[��:�L֐��N���T6l�$h�Q�il<Oy2Q���x��W�(�Z�ӷX��;�im
d�����J����L���2�w�;P��p�!S���1��Z�x`C�L�-U�*ݝ��$x�X�W�4,��x�d����͍{���
��i�����v�JS*΀z�㈜���v��e��g*1j?,*��?l�x��A�8+��Ч�FF�Fd%R�E�I��<��:��/�On,�I�D�&mi��X��T<(��+�<���b�f�2`)�+���z`�$y<���Bk��
ik&a�?��R��ci���gP����/WbJ�+Ю��_B�|\�)�ę(]:#�Gm� ��>�p���[W�C�:�;�{�5�Rp�#w���mn)��o��0}p���\!.�Z�in3_�(*w~;c<V�)�ϥ�(0M4-Ҝ��i뢍dc:�:8Jk��tboͩ�۩�,\>���<x�fr�F%�K`�c�o�eV�t>jg.'=�5�5���J7��m��1'<�p��JCwk�TԢv�a�A+�Fűa�����p��X��%���'�u��;���'�u=�c6��_G>XN��ڧ$W�
�re�b�؟��{���'c�M��C�c2�X����7�E��i��w��:_b�ʥ���<�A��X{�'�-�u��Z@��n|��R梋�F�ag^uy�.��-� !�ћ�ٲ>y�*��m��F�����m^�6�K&�8	V¥�'� �`"��Y�hX���;;Ҩ]!��@�dz�ѳ�δ�*ejb���3�k�f���H�����A�h>��?~���������1x��WJ�:���5�H�ͱ�rP�00B�:�e��f���1.;���N�������_��.��C�_J+M�56���XO�+6��:�n�?��pBM��S<C�;�+��������
�%�;���Xy���S�b������$k��!�3(�Qѯޟ٫�Ǌ������IUb��N����8V�c�y�w�]�z����nRZ��Ijh�}'��aR�g�*����||�΋w�~C���?@�2i�B���L�!�����.�tm"�A���v�ij$~��&!�a����	�S���Ȝ��~c�>eսD��ƶ���s�_�|,ۦb�k>ma�C_�v�v�`W5Z>Ȓ�i�'�W������p��1�X�f��C���4j����P2j_6Y̾vǮRp��:�5q'q��4�[��9�������g��]0d���B�����+���Kk+��h�v�a�QҜ��TEg�T,���:z75Yx�_W#��>�5�5��fI'd���)XB��#Ћeu���M�O�:�1�dt�䉊:.�9��B�V�.`��Y�n��6�ios�r�}t���ڕ&.n&�e��ٷ���_��:XH`�p�Ⱥd��W'���)x��}���X�U�v��k`1_).�4�"��u��b��W.a�s���0�82s���^sg����Lf4�֌�t�&I)���\�����o���'X�{j�������z[��ʜ����_9k"@f�t6eBP�e�z*�M��F���^��>���h,i�a���AF�}\��ʔ����e掅Tj�mIT�}ޥ�-W
|���iڕ1�{cg�Zc�7Z~əJpZv�B-,�O�͂��=|`��<Q+B�.�d�#h�g%�~�uEf���زj�jܩc�dO߮t��Cdފa�f#��,t2�KR����V>�>i*�Y�11����$٬�S� ��}��s���� �R��vr6��V�ztt(_(���CI���ɷ�mA�ae�Wo߉���3��4�։Ƹ/f "�1�ڳG�O��zu�#w�
K�bNX�����{�H�eW���\���RTU�IvO�\rg�v��f�X`r��.��22t�&���}��]=��a(/2+Õ={��s�1g�gN9��қ��O?�5�����@Nz�ucrh��`�TO�l%� 0��Ax�����;݃��?:&CN�-m��4-���Od��0|����Z�>P��Z�޷�㡽o��|��=z`�c!�qP�ߞ��;SO�����}��Ce��`@)��~���o��?����F��b��x��:��|/L��|jΖ�㉭�����pq~�3�	੶���������xy�;�<i����?}��;@/� ��7��y8�5�Vv���F�Z�w�
W���	Z��\sZ�s�3[a�hQ@�b�}�7��jk�N����9�YvW�1cO\P�%��a�
$8[J�<��SA��p�3}��Q��12~6��G�v��F�N�|�bM�NF�F�	�zI�m�к��q�Y�R%��aD����p����`���s��\X�RՓL���,-��s�{˞�;�< @�i�5�*痾y��������p|hӋ���2�:��V-q]��N+�54�~�M�"��P �����[U[�C�j�.>�>�7�5¡�^�{E4��v S�4p�5��I��['��O4SWB�ӣ!�W��ʂ��{��q8z�I&�*)���G���Dl-Az�1sy�p�@�@먔Y����g�aVǝ9=�R��8�,"�]<�I�eQ��H͉�<��U�Bd4�cI��e0QH ��ԣF��M��Teٺ1�LL��R�e�C����"�=�XYT k׳��Im3hPaf}��$��zd�qv*$|�k;��O�������MnY��\Q4R�+�ܜ	Z����|�R��ȀJ9�v��ڂ�m���.ͩ�zU������'�W�F��C�y�rF����o.��]�?�Zz����_���g�+[���	I]fNⰘ]���P��"���o�C붽L��uk�|?��zD�̲���m�\�[�9�A{��DY���Bλ��cԼ̠S� �����p�β��,<�D��Z���tc K�x�E�33:�����g�� ��S0b��@�12��oX�1�7WR�# 8<��~�������2.���������&9z��ʉ�h8�����ޞ��gW2� ��#G��S��8^:v����o�?�����?|����m��O+;�3Ǿ^܆˳�Z[�'K�Q}���U�-#=2�(��"�T�����+\�^˂�=U?�����Z |;�����lf��lD��A%U��]�����m��f�J�o�_�3Υ�U�)6z>���HٯW��~�Md<����L4�م�`<�Zs�
��XU�U���Ѿy�ޮ1���0BJ�g$-r��F���H]ڽ�u�����w`�����'{�+2ۅe��G�A�j
0۰�4E-X�J�M���V������\{D��<��NEk�O�ڎ�-�D�@_�����״��KC(M-�;!~�a��'�\ L���r��2�l�g�i���*��V������2qY�̼���|�^�D���K��^��gG��vO~�i�N��]��hD���CG������l	/�l51Sz��Ԡ>�1�N��d�z|�BmM�Z��Z�̙�Nw�E��pJ����e�X.�=�6F�IhӋlx�,ő�ψ�Ae;'D�l��#�5�A�Y���vQʕv t��'_~^�y�yO猘�?�9({o4%*����c��P.�����0Z`p|,R�M��!b��\=���NQHr�H��*gã�XS.:T���_��{ �� S޺�����2�<z��ˋIxg�֞�,("o_^��0�U��� ��^�����=D���v�ޟ��ù��*�bY*S��AU4�lza��k��!ω�#�����aw���Z�햜y)�����Jg�9�������#�Z��,\���i ���o��D���S��~��_�Sً��d1����������go���s�+2�����%%ˬ��i��Q��g-X��放��ѸR�����{9�i]�+֡���������]Y ���$n����A<��7Y�.J^��]��߽�(Jw�����?��C)ђ-�����2���D�|�:x����?>Y�E�4��|�� a��B�O?�5��m,d�G���>8!�z�N[����㾇R�9��E����R:nYF{l��㱪?�JR�n��D��uX��8��_�;v,����ɣ{�X��+˰#������]em��`�3o+
t��Z5�Ǥe�YV�+���M�o����=X������=>	{�0��µ�^Y�j.���_|)�E����0@��޳������_4vȴDo(�xtt^�y��
���k�o�-�~f6cd� ���sQE��@Ϗ�co�vCL�(�I�{?}s y�4�B��c�jA��}�;ۻ�\����ו�sA�����RVg��=TM����Z\	��g�����Խ��3��G����.<��T�И�{Yޝw=�\u0�)�]���f{eA�J��	��Yl�&՝C���&�����0�^S	�+�#���Gy���!��,W�R�ٜ�A�Xil ��8�gʢx��Ӌe\*�;75�G?"�,�SOT�N�<g)�E��Pl�*c*Xs�7�e���X�t�
R���˹1��Č����G��0g����eƭ���
c0���d��u#�[e�"�l�8���%��CN�?Ec	����et���F4�q����v���d��j9���*�t�g~
w�f-^qJ�u��������9/{i��+sL{�Ϫ|���dԗ�"�@CDm�ʾw�,���u8~ZXFԓ��#K3��}��Em>c�ݾ�9P�9�O4Ԉ�m��m�pzɋˉ����:\_\���Y32������Y�ka��I��s�oϿ{�)�A�Ү�z �T��gqM���F����g��0�!/��G��b�n����f7��X'��W^Χ����[8n���B��kt,k�b���� ����XS�x���4�hgaN�}j+%�*]�G���|OZ ��R�� )j^{#�$_�
g�nT�t�0><�g��`�Plw�zĉJ��u�4e�����ji�od�(��կ�m9t�Q�%>�0�!�1�}z���[I�6�������l���Z�,(�J,�<{�V2���3��/<	��T�6T��
�{e�A;�,=��|~a���*����Z���Օ��tz��i������ae��>��SU����o~��?����{&W��ؓ�#�3�7�x�8�{cݿ����I]�6� ���6�)�1���W�~P+�&3�$�B@��%���,�����G�$��܌���G9JΘdk����y���c��v�I�{������@���`�ˆ�~��u�t���XI�>���v�F�=PhU�nM�Bhʥ����1��������<�8u���SeL	ȩnA�5��D"�2�6�n 6�{96� ^�<3���RV��X�A��:v`���!Z�Q8�D�����of����F��m:��Q���2�� ก5,x����2���@�oK�H˶F�93�f
B��֢�,�5'l�wE�����n�!�5+�� a| �(���=�t�7�̜����Z=�"��e�G�펀e��V��Y����&A���t�ꑂi���
i^�^�8�/��+����l7j�ly��b��'�i��j��)�W�����8�O�lhü�J���'%*��s�Nu�l��� ��5c�X�R��1Ȝ�O(���g mQ6�-�g+,��ʉW~l�L�,�ێ�E�L��pu�čX�+�z��8��h�p�%s��� �;n1[��I4�K�����eG"J���Gc�ck��&:�T%��>;{��_�s{����Z��Ͼ�=z^�X uj�ñe���0?|�mx�Å@�������p����<����ヽph? ���}��v�I7���a��7�����{ԗ}`���*��������E�?��h�ʗadA��ے5e¤C�}_U����]P@�(�ٓ�_�-��"<�잌���z�8dZ����"|������F�������P�G.�Co�e� �K��|��{��͖����y�Z���Fs�{������/uq~~|��E;�gr|T�����s��n �"4��%�c.�p�WJxh�ĥcD�^g�j�%��뤄~�~�l`�4޼y�L� ���c�DS��šS~��:t�Aޯv�u�Ƀ״�=�.� �>-�O���Nju��v!���������z`[�HH�k���;��f����C/����=��P1�)�0�v�9G���Cj�8_�&-��,�i��`d�g�y�o�z�D>�R�e��ֽ|�	T���S!e$�;"Ay��e��0:��l�6�#Jq��7�����ɑ�Z���^�l�A�'3�����u���Q"��0#�ۧD�U�	��Ҕf�`' ��r�]�F3�X	dӈzM�y|9���F����;�#�ԏĹ<|��2�9sH?�Io�Co���_\��eI�M���N�Ȟ�C�N��ϙ_^����'�Sʰ=|�Ts�d���8<�կĜ�1Z�%��E'd �i~p=y.cF����疝����WjM�;�{�  �������u ��޹��»�+}7J��) B�Gǖ�Ϣ(�|��W���[ ��dD���r����m�����~W�TU�/��+�Y^�,&.i��=."y�s0�|�fʶ��t��EF�̲@D������1�g�=�<~(.��|n�[�k3P=�o�����ZDǀ���k����g���9Y�栛1�yD�S	�W�N_���Z��0�-#��<U����F\�X����b��(K��������ek���1�v��W��>x�4��*�/V�*hȦva�[τ�c؞��:\]]���4� �"*C6���ࣃ^l�j/ 0�����g?��gy;��$��d��V�Ŋ=,���k֫�.3���^����ZNu�oo7?v�&1�f[��l�J�J�IT?���:��F/�y���z���7P��ę[<�v>(�c��p���R0�˝Jdi[!�R��0�-�f��;�sjg�*e�Ce�:��3lڏ8o��v�3�a���kB[��/���(`��NA���w�}>^)�
�D ;�o+Bq=�w����r�a��3�r����X�e�����߷m���睙��چm�7�V����C��Tsڥ�n∑<��ttt~�������m�,	����FsW2�T����2���H9��Dz�W��L,{��ќ2�amۜ���Ti���,gX	�Fo\t��Q��4{{re,y=xt������ϟ�GO���ކ�/�$�j,nW�f�ʭe:�d��e�g1KS��V@J�h%NS�c��uC�رs� \�l�L�L`�hw��X��:�����0�
�m������nn��]���j���8��؜��J�8㫷�r���
ǃ!t�䧨c=��Y8|����U�|�V�_(�����c��$�-��Q�����ԟ�������?|^�y'�ǆ(C+e��Xx`N��wQ�1/l�	Pޘ#{gk��
�=(_|�N��{�G�`|d�y�z�}��w�egӉ����,��wo��ŗ���;�С������*�6�~cF��D7��اEd��w� ��7߾/^҃~!��Ms��v/���Ԓylk��'F��jc�����g��7ߛS�i��,G�ֲ�a�cY�q��h_��q�vw`�څ^S�0S^`�F>�1�$�X�3�{ױ�rx����噗˸�j�̑-a�+K폛ɍ�.��0)��ثm��
<q��͹�k�x�e��ϴ �}�}�A#Ud�^q�0��0Έ�{�����e�݆�Ёt����~9?��3�~oՔr$��R"��'ՙ}~.G�c���������D}��aoolA;�����CI�R]�8ub�Ϭ��'C���������s�����&���ֆpff���� ��3Nm-7[d�2�����,&	L�H;A��E�gf�c�l#�g��9?��B����҂	�6Xר�F'Ju�=��c�ߏ��{ٞ�i+PIS�<&d�W�A���cK����:l����:��n��pU�J��=���ֲ�O��V~>2>>�/KlYzOãi3cs�e&U����*�-;���*�h���>n=�
����,�����H]��?�7�x�\^�+x�m�X ��|�]�3,�5����	Ѝ)֭��R0Б���A�{x,>q>c�v-�9��eڙe�?�}f�#����s^��e(�07�BO��a\9-l�t$٨<�n�[}��|��4$�H,�L|6��ԝ����{�
T2n�{oX�|iȞ�w�kN��ٻ�p;Y(�ҳh7D�L���JV�� �B�B�Dꔙ�m��_ˊsczr=r?BM������l+'Y!pǶf��q�ᴧ�pa�Ƶ�N�0ht�@%�2*+�]q�^��支of� ��K(��\e�8��������}	r�s{o(�~z�7�e��P_NV4Z74̭��k"0"����/�Nv��45@t��@���?}'v-x�7�� �?x��홄cw��S9V��.n����ٍ=�f�mk���GG2��<D���ӳSs7��b9��$�J�Qd���F5@�w˝::�GG'a>�=��LVd<��s@��W��@|~H��.��(�X �=N���5�]��ҦM�=��9>sbǏ£��5"�a8<:��>�`	��sG�j�lM;���g�`��Ǿ탢j�����(�Ik��nI`���pі���w��UW8ʴ�y����u���g�}��3����^軼� �EC��@�ԇ���2n���X��/~x-A�\% ���[MctP˳�R� � H�x������� �ҵ�Y{{H��r���i�b\��ӵ�����|�O�R���'4{_}g�;�������&�l��p�<��	��q�bϻ�Օ�:����P� x��H�\&��q�`�ւ�����+�}zp��C�K��<+��P���mF��Eq�<O���T�kZ�66�8���4����K�J���@MRFn�>y��3O+$<
Z�5]݄�1�́S�GZ�^*���z2�m� �RￃA�s)�MÐLe��`�*h$7͐O͠�m0[�V�T۸k�A,��N-*MފU��������d�8�l!�T�J͞�?�V_7Q���Β$*��g�����$N�����*��h�t��[���3�メփR���0[I����k 
�(Y�Jg�Ό���*4&��H����-�Z�7:�� v�!.��.�9cz���{,#����'F����F�4�j>l�_b��(	K\y��٭�]�A��@�h`F�0���C��l%��f�Ͳ�l�8�,˘��]�Z���g|�n�h-DF�3�+9)�g�=%�d�݂�` ���3�y��ʪ3�?��T|�N��*"�\���ڕ1w#;h�G�I?�7���g�`�88y(r��lw������ջpfA�f��*kT�׿y{��}��y�* |��f�_��;��.�qb����>WP1���/~��U�Z��k�=��8v�ݯ��ԂdM@�2�Ͼ�{��-p���?�oN}�GE� ��>�Cu�`�̾9K����.-�~�Y{���y��bCF{gme�T����;��]�N\�7�������TE����A_T�����kUO��k�i�^{mA�5,P=��w��Ge������+6�!a�Rh��zܶ~�eޅk��e���E�ӕ����A;]��fʻrԴ]؇_>�\g;@�q\��Tnx�K]Bx֔j�S̲���BYu��&��@�+d����������۳�ǑD����Jl�y$f�8;wi��'��$:E)���l�!�SSN�=��,X ����ǯ��H�U���ڢ�K�V���A�{<���_����	��'*��'���E���V���imTf'0F�R7eo�D�� ��~�浽�Z�Uƙ���۰W�ޫ5P��$f�AX/��2��}��6|n�pa��C�,�r�͐ލl���O���Z�\�ln��< .� ��HC^Fq	��]�\M%	��i��倒<$���a+���-�h�Aܨ|��Nؐ��S=��z)�	8�d8Y�3��v��n=���d�x	�l��_G�j�❔! �@�P�p8?DP��j�ψ��|��')�s�gpwC�\��J��:�]o]��C��i¼ǜr�F)�d��Ỉ`HV��W�k�3��ͨ�j��LK ����˕�}4o�F��$�:k�h�R�d\�AK�o�8w9�����N�RT*�l��y�0%�Q� ��|ˊTp6y�p�	��,)��ID�H��Z�O�3 ���KMA�áe�j��Z��d��Wޯ$���*a���e��+1��=/�C�|}sޚc|��*��4�{-;���yUȎ�Ó'��"j�@�����Xi4���^�Da{}s�{�'�D�s~q.`�vv <b������\�3��~�:�YVO剽SKs���ٵ��0��S�Y�K�A��?���s�
^_XPA�����̉h���g����Z�B�	�����T�OUa�k���"�I�q�|�F�up�u��:E�w>p��6�йW�ot'�H��]�C���yo���U�CU���??���ֱ=��*R<�?��g�0�oY����tv(�zR��|\B�)��I�����Wr�"��{���k��}ma���s?��*�aVB!�)Z�,r�t��qx¨�vS0*��_���o�Z�~��˸�oQm��2�K��Q�"k����_~��dx����v�*��Nɕ��Z$u���(Q��7;����Y�����饲�|��3��2���f}�~,��f��M��߶�@����"Ey�����b�5!�X�t�������y���r:��t�w���C���"�@�C�4�2���\�l!ʠ��N��bs�B����,�p�P�]�߷Ciy�}������PH�N�@/55 g�v�{��pG�~j�܌��\sڈx�W(s?���P���,��^3���|����6�f��s���t�2.*9����@�����x�Ke�)��M�(�a��G�+��ĈB�̠�H��u�t:_����#���7ֺ�5 ���,]��Tb���+R�Y�k���y��'��@�[����%�]�R<��!8xy�L�닑����Z>)`& @*V��t�R�0cM��҃����PL
!�oh�e�8�{G��.]]�^BI���begֲ�Ks�7Ӎ���b�6�C4R��-�e�:�|oŲ7�O�x6m�O��4���T�l0���gj}� Ddm���1�f�U�Qh�cݚ���Q�$��S��)��*�;U��y[3�ө�p~�����3�����w?�P���3�>p�RX�̆���)��Hޗ:ke�=D����Rg6>��&~�K���:Sw���p)*"LU�Ukvv8�_vlm���{�y�Z�#���o�/�}��ת���3�:
��{Y�SͣD�@�B!���X�ckG]�1k�L�?�У�u��q׫�0���^V�B,��?,�,�����2\��p�a�Xtl�zzuFG�;���»�o����fL��,Sl���f�5㲘^K7����֧�Zd���1pY2X-ETB�	v0�c��(�-�F�����u�#�Hámb�ʍ�~�$qf�9ol�ns/�3�s�g�5�1�8��}/�}��y�?��'��7�MD�ǲ�hj����R��eq+��Ū�ő�JO	�"Q&N�^lS9^f8A*O&-Mp���u��Uk�ޢ������R0��>G����|2i S���-�&��;�0��Re�y���Z�`���r�Iʺ��F.�cK� К�
����Q�7H FT���F)��QĽ�ZQ�J�U-�(��@�ZN���������ߺ(G��H�.�1��>���������@�������T�E���DV��nl����U� `�����h]�ڦ�#�#J,��_��&%U�A�	�����bs���i3�_>�8�ӌ��u�&]��S�I����f�s���q>7��r�m��#��
g��+)�it*ft�G�z����ZI�<�"���չ�ƪ;�@�,Wr�d�{@5�C1pjז����'X�������n��ׁ� �C{��j.R>[��4��jB'Q/�(�e� �\���[�S^����W�胦j2��{J�3٢�b*��Р��B7�,I�f�L!��+�*b�e�T��oť�vr>��,i�@��~��8���"���]\9c���>�/Ǿơ���Za���p���!����H|�{�~5�ϯ3����/�W�������o�%�~n�=,��7�1 0V���'��$:�[���D�ƌx�>���Bg��ѧ���z��Ӆq�i\2^�rš
�1�~�Q��W_j��#��"�ɏ�4"�s*�f�T����c�Z���3��9M����ckc��4��$v {a�/-׈K�6_�N\����k�0ǓE�E��oI�w�a+��1Kp��,�0��j*[���И.~|N/Υ�M�zZ�㎏�=�3�n�e�s�eC�t��:ίRj��ӫ��?�G����Yã�9(t�I�C�d+/?�9�҉#t��Z�>�P������?"���V;F|�(ue-M*q��iw��,c�;�g��U�*v�"u�aU������A��&�$�y.]�4�e��`Ek���
�ǞH��e�R
T6��f�N m�X�f�2�����n%�d����cO��Ъav��JSW�J��i�����>-b/>_;��z�*n��$JKPd�Q��i�Sߋ�Mb&�$>Mq;D������:��o\���+d�z?�Zb�c� 0,���:׌lJZ���R-��k5�T
��M��K9�j��It���*�E�%3�ԃ��-kU6�� Q��H�V��+	�,��R��@b��6���f������/טH1�[%�S9���E�ݺ���F��c"���k�����	")�8�ឰ�'x�BҊ#^�Oi���Ѽް=y,���MhPI��稌B-u�����i� �Ԙa3�T�=�\���1�Q9���M���U�C���Swܜ���E�+��f�������M@h[�ɒQ�����qh��3�sK�� 8��!<A`-�u�"ʭ��*O��W+����[X `N�"K&���%#�U���g�E���_D2�ѳ�1u�1,�ӿ�*|����s@ls��)ur�Z�.ÍA���G��fr�\�'���Ԣriպ&���.����#���3���x�xq����б�������K��{���v3��M����j���C;H�mG:�dkJڀ�l����\{�m��}qc �.�:�[�4�+�� Rv NL%�1T�t�9[�� �-|���PV�4cN��њ�$*vs�8��оl;o��R�Y4���RW7�h�_��IYsc�݌D�����|/�])��Wn��8l`�U��*D�� ��&篠�)��=ow��P5�+eu(�ɈњH�39��L�1�O��p%�.�[�bv�Jo� VqR�*3�`:��>��T��l�}��:ѐ�9�����̺r2����@�c��G1�y��]8qN�����>5�Jǻp��<��s��}�ۺZ��G��Ͷe�#�7C�䪠�O0��z\��*�_�
	���N1'AB�U�JI����l��Ñt�}>-"�i��%���6�EY��j�-<i`M��9�ī �!2�+��mw�R�ñ&8l��|�)���^!QA��
^��)m����g��;o������ң08z;Ӊ��lR��ۋ�`>]կ /8���^�xy������*@�AJ+�.��8�Q@FTu�IH�JR&6=���l7���k{�c���&	,5S�:`�X����A�����eB�g�����!�Oq%�>�^^����m�#C�`���s?��C�������G���=�2���0?{�$,&3/��62\�n�C)~��N�:������mJ���9)#��ץN�R�,s�����U(͘`���ka+��]�dc�ԫ*nIR2R�&.$�Ԡ�{��É��(���8{U��/4'Z�]����?@�&^��l������N4��$��A�}���c-��pb����"y�cy��.�D(\��$����}���-�Ʈ,X��vd�p�k88KZ�e�5'�9���,�VU��KD�$yt�	U���ƞ���Տ� h��e,���|� ��Ϊ�Xq�˵�?�5dx"���[��Q�59�=��s8�/S��R���!{��IK���*�!���$�	i]��;0�¹Q�:�@�]dI�	�k)J�޹(Fs㨧+ԣM�sQVl�Wx�Pžq�
�2S1:_:i8������J{���äKóٖX!����T[Rg��M��6��zf�ѕ�TWEx�Z%��'�8x	����q�R7t'�)smJG��ʿ��z��<6S)���-9���� a��3�6�S�i������S�������B8U4r�P'���bë�ZA�|93�K)�|�����)�ɤ&s�ӸC�#��=��n��:6u����Wȡ�M-g��.k�m]{�s���"Rnץp�J��\8�[�nC�I|O��x}��ؽfcW�Oj�{�l�����m����8��~�š��3R��g6�m�E�5$yF_~��>��̷a�C�����߅��a�'P�|���lae:b��>{~<yjYwO�d-�V3J\w�dA%��"�n�%Ź]�dpP2B��*$qҿ�w*1�^�3��q�D��J�m��q_P���~�������{��'!Ck���Z!������Ȃ�W�U��6��ũ���:��4% �����3�$d:�|嶵��h6o[r|=����FÊ�7KbmN�HUj�c0%�Z�k'�R�_���F�))rBZ;S�[nc�t=^�0#��웈_�^��A��2lT7J�����F��	[Vz��|ٿ�0����;B����"�es����ⲷ����3VC��n E���~��jb����6�dj����e��1��
��nk\Xvz�j[)+T���e��PVy�����S�|E�Xɻ%�9h9�x�Z���,�ר�K�~8T���ъ�J�eL�źT1x���	θ�S��>��SD�)_#Mc��G#�b	����>��G�+/�xKc��0�:�� &�K��<�~�|���QX{�y��޼�H#0�˦X�;6�D0,��"HN��Fᦴ����;m�ꎗ�T	���mV�8�q�F� 2��f�[YG	JZ��Q�i�۪l��&9Sˉߗiܛ�8��&�O��B��SPV܊R;���9�8 �Ҏ��#5��~�Qe��Zּ�VO�h�n&=����#�gjg�����Q�W��F��Gv �������������Dr�]s�(P�d����}sٹ�b�`湏����ax��A!K	h��|�(?e�(mү�Ĭ��?3�W,�|^xjA�f���h`��({�Bqu�]?<#�Wf�7�S����C�R;��1vO�j��sLR�@�?|�P:YxN�A\ւ{�Qt��i[ljr^�g8�-��\���֬�v��Ժ��r^y��mE�ĺ&d��z֘5��}r��$�'�]�P�+rg�#JG�!�+R������U��:�)�[�.���� Y8�ւo��k� )��sbw�e�s�g���t�%�9��E�3Q��$U� e���y��n��2Ϊ�D"�L��J�*�HZ����_��1���Ae�)��Ī��G�G"G��ܚ��L�|hx ��]F�h��L	l��Ң�bf_��/��B�t&(�tۮ]�8��[F�d���PV�*� z���՞*�P�AJ<)u�|�=�-�'!оmy� ��ҫ
J�ԧ�)���;+U���c����v���6���/�wT�5+��9�8��Չ��mWU���Ȯ9W��m� \Q�C9S%5;ؖ�L"��g�0N*ݴ�Jay6B��{pc{x��ⷈ`��GD��p)�3e�J(֞�Cm\ȑۧ�*U3 �J(K��82�G9����o�*���dߜ���޽U���8	��xGM{?����G=�F��Ы���>Q���Y��Vj{���s?���5�3� ��~"SڲH?���Yd��g�F����������>&�`��Ku�&uU�T.z��T�!d�ݶ�p&(�����8
�e��b�����S��m��5�.D���ʑ�8�6�����p���{$q��.0ؕ��B?��W�Ϣ�^�� �p�P���k���ʿ�n�2a0�3,����3\͢TO�$���'�}���g��f+���T�YE�@���/Ʈ�!�R��	D'(�M�xN6B�tP,{)c1 ��*	B�Ǿ"F�)��I�|�w���T�����z���l�̇�Uq�W%��pT�a��� ƍQ0�x���y=�&
D�S��	�d���=�:혩�a(c�;"D�� 4|�A�'2��Alj��AQzW�Ի�á�+��3��<�	�V��!3���BH�4[��Q5��9�*�&A�*PAQ��G�/	�,�D�1�T�~��V� �~o�u����� W�_Xē�eMe���#�<l�27sH��
A)%ۖ�.�`��Ȯ��T[Z͖���;�4��N�g���.@���Z��θ��.?	���U�� �Z�n|�0�z[�
K�w{� �v�Ί�i"w���H���J��F�i�G[T�b���Tڔ+���m?�����6��&D��nD�����8�"�$P%��*��*���O<�Ji�46OJU�ѭ��4�?ͯ�f�>$���I�fh{�(:�$N��%(5	T-�RF�oJ^��N�<�:M^����ejj�B��������I8t���䙐f��2ٰ��j9W�[m,Jk��)
胃г�Z3���R���E�V(6���wa���Pv���Ҋ���m�={��eW�e%M�-LI��`�;9<e�g����~x�4:���o�T%�dW����S�?/��3�aǠt���C�zv�'�>D�Ϟ=����n���!�{�Α���J�@i=����4\�|*42�c��tCs�FC}���M0x���?�r<�)��\�l3�q����Ϋ����v G�������PW ��� �XWT:tu�Ym �;%'���]�b���Ѽ ��c�x�w�^zD&�o�<���:���]i0�F��ey�����l<h��5\�F�=fk���G�"�V�d�Ӗ�t����v��M%�{0�{��,������7�&��I8���1�-:*Wu5ɮTv;�X/��(�g�N�;�,�r��<�|&�b4V(�ʀI�I�|���߯���������q����	�1��H�𑞡�~d{�w�ٵ�=q���W�ɬ�h���C��aA�0E�kOA���|<����� sfM�bes���b3�ϧ��ED���Jv�����g��Z⌃j_�gQRC�����e_���^^����LQ귙��3����}畦y�� �d?��9k�������䃷�Ļ�9���Ipt�|���D���'�y5�̎��'�X]��*�F�6�"�^��s�Q�^mH�{���D�[L�D��	=>	�nv�~���M�o�-rC����ڢ̎efi�YNÄY��b������X�Iƕf�I����� ����fl;p���<,�'�@�r����?]��3�mc���B
Kq�t�^�>��Az�yU�vǓj�S"���F���G%����"�i݁�w�������񧼇��K�����������%$<���D+�΋�*�/������;A�3$@43�{�m]F{#�oJ/�b ]��uM��s~��k �����˻	���ހ�z�lM\��r<�@k��?m� �<���{{�ܷ%e�֝jS��Xsdm+�}���HX˝`ľU��Q#��
�,4r��?�4��>("xr�ߵb2��H��&��>�f��ƓTa�̛8�ScM̧WN���/Jߴo�&�ܜ	�y��=q������}��Q�z��x]�L�#�Ύ>4� �)O�����E#g���z�P���IT~�b�:��M�a��ػ$���]��D�U+}��8
U-boVh�a��+��f�s��i���ĪOm�Y���nEj�B����W�]��KP�Wߣ�P��>�Y�
������:��~C`]�~~��{<�M'�aV� �jj�D1����5 ��l���t�r�y*@!���01���T��	�H�z�0����s]�;��YXO.�q�,��j�����'��`o��+���
V8#|>���N���%�/���=�g׿��+�<Ѩ��r�}�[��	�%;Z��w���KNj|lC�;n���i���s�l��'�#�ǧ�e�3�U'<���r]�������Ó06#�)�r��xM� M//����(A��yQ�gqd���5s���>����n��O�KBU�ȧ�04�Z��AOQ��z��!��B�R��JInl�ѳ��\���e��L�~y���G��������w@ ��ɐ����>��,W�N�%�R�}"��d�E�f�:�~+��Sc*�7;�жlg<�ml�����D��p��W��"w9]X e��ʧ5>��3������h1��kDD-}�R���d�~_�b��-`�ӷ���Y]��@0�`�F���N0��r�T�STY��)kL��A4�W���9F��\ϝX��@�[J>5�QiUs���9�%���>�pc��x	,h1�Ʌ�]e��N�=�r�9�Js�?��OG������f@���^��3�^�a�nZ��w�����WC�ڛ:m�;����}��&:f��UҰo�g]�{��|.�������4Oθ�	JĴ���� 5��-�(6�G��8?T ������	l���J4��ŀ-�_�i�1Q[�ۚ�R�[�>˚}Μ�T�U���ru8)I8{�֖o!&H�qΙ�$��m�'|��1�kf�kv}�3�z#���C���s��=11V�9��U��6'ξ�q�������F��J���G����pO�e�8d��y�h�cWJ���>d�A�k��U��B���E8��%�/_��z�K;����vj����g�����6t�U�����=���(ڹ��Z�+�$��}hzu��1��	I�:��Q�����v*�8�k�渜���l�����P'ܪ�uTO�v�������GQTdD�۵E�+3�v��U���������yT��1��8��9��e�H�px�%�V�CLbt{m��P7�̴\`��ц��Գ�6Dv��e�C�9e�2u4�c�����_�H�2F���ß��������:��KR����o�O]!��W�(��6��߱5s�����O�Q:�.����}��*�/3�h���5�WW�Ci�\]�=ʚ�֌���~vy�ځp�A7R���<�����Fvvi�yqs6��2u�s&;�2'�p��qD��>3���kUuq��-F	={"p�2Y�9����p(�eIݛ.��ɡ������^܄ՠ�Z��(��Ep2��2�{0��\��|&�7am�-�2 X3[��Ϟ[���'��K{�ջS���w>԰��2��7A4�	����Υe��<�@WxE�=k�������e��ᘑ,V�%��K��lKZ,�_v'�OP�wt��}���G���o���̲L S-��8
,#�l䖭!�E�3k'����0{��uG#-�>�KI'�,}�-oo�ϵ~����$D6c��D��#�n��Rm�˷oT���U���z���k�<�}4 �A����Y�� R�&���	�F�c�
��~����Y85�u{v���q�#-D��}�>m�rc�ڹR@���g�.�)!��$F⣀���	 �<>�S��u"x U����MZW�����ZZ ��s�F�3L�1�ؙ:�
��cؿ]�=�}�g��;��fv]ţG!?�7f;�ښ?�\��/-a]X���2�r�7Sęl���A�d��i�2ɵ�Zm�jF��b�xw%��Ά���5�(NS�qrG&��v:���~�Ԗ��4|d||_6�t�(E��A)㓔:��w�,�7n��p�+jW�ڵћ��)E)�^ZI3G�v"W��G��[Ep��4 ���4���ƤrDk�T�]��f�u��F�ߍ���}��}g^o�?���kG^?�R���q6/c�����J�{�B�.�i��j����lk&�N���g���R0��F��������7h�r=w���D0-(���ׯ�AG'A�N��^�9��p��k�xf �pL��2��Y�_�~w�T�kw4�Ӱ}BF�ѥ�\}Q�G�i,�/#���&����[�2e�ڜ�ʾ������á�[sr�d����q���y����#�nG����d�'����3�W��� 0������-�����Aٵ_��T~.؏ӳk��f=��n�]�R�:G�Ů�E��̷
*s���͑g��x]���Tƌ3G�c] o���΍ߤ̷���]b"Ǉ�<�v�W��
�J<���z��Q�N?
�Ok��W����g���+u�̙����=� +�.[vo���7���q��CU���0<:>
�`��}�eK��!�B��<2�u3K�*��<ОXK���� 	�3"�dd߱Wǖ��- �r�+�R�Dw��t�sٺ�@0&�> ����z��Lm��$
��zpHTBF�g��C�����2�d� G��K�Tnjt}�P�3'��ֹI�	a��iH.o��i�ut~��}���p���}_�^W��jn��]'�Y�Ԓ$m�Γ߰�D��Ｆ������Q��9j<N~߲~�t�5��(�?kK����U;�!Tc��E<�)~��F�m�;X�x|]@шά�zF���-��	����>;�?8G�Zt�fe�"ء� �&ˆ���@i�Gl��Q����̢t8��6m8�J�_��d��
~�(cٰ�XU����;3�qWɮ��c1�z�K>����u���6q�|?,�כ8���^ Q�e��{�)�2y����Q�w���H:4;���@��5q�9� V���e�f$<ŨD����jkٜx:���)ܚs0�}Ƈ�>�9}E�]�.o0���?��$��'��Y�x2�}3�+(AQ�
A�L��4��?A*�A^j�7�}��}�vÑ�*�c��O2���i��ۈ��.�.�7���v87����p ZS`�*J�V�c��h�j �T�T_{@�����i�UbO�47wd:��kXC�n-�ztH�bt�r�/֯�,�@8��R�Ir(ueC� ��[��2�FP��*�ٴ�,wg"���6T��Hcj(y5�*�- 8:9��`��{JҴ��r7����̍��>���ص�nsqm8�������<�����F&Mt���ͼʥ��`�75x������I:��bR�S����y��Zc���l���A2Q9�?�`���ٳ��j
�ߎhrx��nof���8���P��
d����D*�8��Ye�\�\��y��L�R���Ѿq%�\�a\�Ϧ*���H�� �'���QUɅ�5q�*,� ���p�QH��C�?
{��Ȳ�r�,�|��4��V�(A�mY�j_�!l2
x�����?���g���C/�K}���ҳk����
5����}p��F��϶�BS���+y����؁��hm�B�B,�s?r��s����W������H����8����|��hK�I�>=��
�ۣ�c�x��y�X����"�}3:O<�(�fp�/��Ҽr��"n>Q��֛��{�f����*w�c2�z�"|�i�#�F
����]�0[�5������?�H�������g�w�@�3�^���[3 �Ⱦq�_�Tv�?�x��G��*!Bȓ������{��$4�f8���3f,f��t�/�NJ�df<V��I�b)�6զ�C�qߍ*��˱3����H��5wn{$����T�?8��|���!�ӬRYP$$���Ȃ�SƬ�*�����~ڔs��*Hx��7�u������F�S3l����ǫ���t�X�zkA�e�dU���á0|$#CRg��
ſ�4�5�#��=A�v���z�@�"s�v�{�,lB�c�A�#EK?T�e� �83R�2'�����J
�����n//ԃ^[��?#Q�����?�Q�R~!P�r��QW������-(A��z�`�;l��R-��p��BLg!�U
z�!*��+�GeOkܫB�)u�T�o���C'Q����ߊ�}��r����f�J�d����T�����x�!\�_��}Ɓ���g*��-�Դ��[�����~���c��8���i��+9���m��$j�؞���H ~�C ̎�uf�H� :sT{���C}��%�*���1�2��B����������gv|@�p��nh��D�K+-	jW ��l�ڇhQ�Ԫ0�]��Z��x0�Fl4��|��I��O����*	�x���f�2���=������rH�>����|7��I~������s?���N�9P����T�g\�*����N�}���Y�ч�D):�}�({ ^,��&ւD��9�}�H�wd�������Ł�z��-B�u$U��2��ɴ�
�?�B=C�D��H��#�s�Z�ө���vG��ay�v�u�Z~ q1��i�v�����$Q�b- Y��۷�MD`LG����T%���-���*KRƜ\\��rP�m3&˛�J� ������Ɯ{\4��.F��%�U��N`[['!���:�D�	�E�D��<��wQ���w�9��ߔ��K�&������A�2�\ng0�Qg�O�(q�'��}fî�lO�o�� I�/��*X|�LP�T���ϗҏ/�P
�����?q�G�q-Im��.W3���V����m���P���3�܊sߚ��� �[�+kIG껞vL��6�C��9kʈK-�%A�Ro���.5����㉩����Z�[_D�ޕ�S�]��!��Xa�jWIáK疯���"rB��&�)�s�[G�K؃{W�Yk���Q�T0z��5��<�)2V(6�b��Q�O�s�z���5��V�>�hk�	����ռ2ߏp �j��@�#�E���(���}�o#*U���d�0/�J���Z�����/��Ɯ)����;���T�Ƈj��Y2�wu��vWmM�(�sƀ5���&��h8Aj���}�:�5�J�<j���x����:Ӯ��hﯛ�e���>��F�j�^�MnLQ������ė8!�u��	�h���hJ$q�ӫY/M5�nW��`Y�Є���Y�ƈ �0[n�b^D���v1��ܪK�Ut���R�>���{����8�Vg�I��x����1̽?��}�4w�������\#���B�������eb8 �&0�B����p��V���Q�����S/�azvnm�)�0��m;8�}��,�������x)ݫϪ�rl�;��-���i	�vb�8�;J1���9`�8q�7.�e��A�/�Ͻ�q�;<�X�ȸ[������K4hߩ�7G��a��P$-׈{ �c4��^R�M����%��?V&BԽh�*GL�t2#ѽ�9 ���е���TfP����Ke$KjHr�Y�0Q3���H׸�/w����q�E����t$/J�-]k�E�_�i�����hO�G��{�o���)�/P3���!�r��e����a�Η
 �q�]8��x/�ep>��j|vV�n�8���{�|$��l[��P����kֹp����f$ui�ۀ�fG�,�&X���*��PUiׁQ�P�+(b�á'�S^��,5"M.>A�������V͔��K~�����j�s��I�7߉?�2C�_��6�D�p�Jx�Tb�e�\ |�.Β�Bf�m��`3i���k4z���~V�'vo6��^;�������񃐷�����j�������K������Gf[u>~��U<�r��Q�;B�s�>���:g��DB���es8#5@���8�\UU�:s迌���x��#�gTK��C�p>h��*�&mrnW�e�W!O}Κ�ֵ<b|�R� X�@Hg-��8j;8�+���߂�ԥ3��"]�c)��HL&�+��S�gn��3$�@ƍH��޽9�:3�>�����;�*�����߽&
�w��}����� �����u��$q dt0���l�洋��VO9��'�g <��7d9(pE��Ep��Q�Ξ�*5[>[*��r@�6�BR_��ۂ�5�a,�.G
5��\��N��n�"�i]y$�����vC_Y:�6�Q߶�6�0@6���l7��Y��z�e�vtp(}��|�q�"�~3,�	?ęW��R3���Ʈ�.ΝK[�`&���5O��釡 m��W
sdJА�@�[���"[��%��,��8%�G0Fz�
��O������T�iٍ3�>��3C���{��9#�U��v~J3⅊R������
��H'���7�l�aG|�6uUI�E��vW��10�h�)I�}䴾r`������@��wf�n�yw~kA�T%���e|}V�G�UG�m?��ki\1� �m���y��e�,8��J����[U��G�B6�LTԬ�ֿC�xM	����^0.�t@#�e�G0ސ�I(�`�R��ۛR�=��t�����?Q߿;4'iA���:dG{!x�ð����sp� ���jg5!��c�7K4�33
@�GD:wI5�����j���jS���Uź�~��^;��.u;�[�=M�Ρ�O)~hA��������]]���9@� ���EE*�AZ*��n&aa�rr%� M��h_�O�)�޾n,�";���f���4\L���$H�<�܄M��zU������)ÚacL+�x�*׀vf2�7G3[}s��e̠/9ֆ�fE��2{	b����w`����lq��?w�b��c�a�$�1�
WJ[�\Nnl�ɿhn���ٜ����=�'S� �+ƪ,FÁj�<���8 (ʈ�F�`&Cs|�r����1����_��P�T9�%b!���lL�"�J�.U�P�d�n�=��D�,f�������]3�*Ɋ�p���t2'�bи#��=[�=~3�d�U��$���@U:�i�^5}c27{���U�6�z�>j+pQ"�b���-[��Rՠ�!j�B�b�����yb+��IY{�����-�h㦫||PJ^�,ǽM#=k̐ �L�\4���r��Y�=�� ��	�@�t{�ke&�*������	��#q�H^�cc^RہR�����8���2fj�M����J�8��IM4�'�ڭ>�[~��k�
_"���͝��ք�<,��t�W5����}��=)P5���4�@C�3��֔�9ai�K����w�;Mv�8��'Q�Ev!�I�:��RQ[�Wj�mb1�7�%�L?��N�p���߆��$�,���1��G��,$�fc{-�o-"���k �mBr�����j�낶��gj�~�.��q��)nvɅ씭���].����dA��Z	 6Dou
[�~���jy��ll>	]�Λ��
�+o1*+�%YՌs���ʈi����'���`e��)��eC�81#��"ا�*>˙8�Ŋ�t���\}�2�ft)Q�r{-b�d�&��Z}q�{���TbX�|�R7�6�2e�?�4�Q��$�����V�81c�b�����_���B��H<X(U��oa|?��U������c "�^���wԣ���+C��J �9�+Ǆ��iI�&I���#��b=	�2x��*�w��*Ѳp��)U&�|&��,࢜�,�����$��)|�8�ʜ�|��Q���KK�42vq81$�痒�X�,i*�Q&c׊h
e�"�k�w���%J�.0Se2�U�h�Rԛ��")jB2S�.�k-�?qEQ��R�t�ߦ�MI־7�7-H��>���L]�@�%<uc�E�7�f�E���� ��r�J𹃣��NoDHS�%Q�ʫD�I0�|>���w.�6����dQ����.�?�QU!����3⁊�	�PѰl��շ�^Pn��{������m f��T �@��#���9��:������t�QY��`���&��Z�e��kI4|8�-P̖��W�T�#׺���RQx�������sք�9ws�t[ι�3�Z��@�2=}�@��>��|1��9�7���m���
6�f,uV}N �
"JKQʆ��HT��[�f�iĲ�>=���$#�/-���ʜ�7��{�6[�ѱf&���i��HC_���9��ǥ�ѕ�U���0�"zm$=�V�.���O�U,5�"2!����s%}���j۲r�0��~5-C?@���J�֓($^�.$m�?k&9�\R�>%Au���$^�
>�/7�����Ͷ�̨~:�O¡��F J��#D�Z�w�q�i��{�k���~-R-�l�p��mۡZ,&�S��)��_�]oP�$UM��\��Q����>'�T1�p�E�!츸�-��d!��Cm��y�t��w�Zv}�ԣ�:������x�f�	�v=��D�b�Ճ{҅�]�>S���}?}GHZ���� ��z���{Y���4�,&Z\��u���fV1�mJq��e�D���f���iXM碞mF�s#�S鮙(�׈�1�����Z ��p�Q��-м+�ޕ�"(��2c��%}s� ��{ҲC����(r�����q���{����=�YI��k��i~!�SS��#<>}p�u��4#�;�M��d��{YD"��W��|!�C˂R�f�̌�HfN[C���,
o� 569���^EĈ͜�V�Ip��앥�b&T9b;�a
��w�bX�4��0�<�L���&,i��ɱ�l�!&2�ܓ��0�N��s��c��N��P�g���-��ݪ�D�M��{�y\c��'��������L�0�2U��6}$���f�چa�-���͍�Νj�K�7���Ǒּ�TP����pc�YN�1 �B/�4f�w@X���.L|�jYש� n�
��Pٿs�=���g��>ǂc�� ��ڻ<rv�j�6е|.^UNtT�S��\m�Fl3n��g���r�C�\x=y�J|0R6���a��Vl�!"(�f� _63Yp�k[�u�g�v�'�cT 3�|ꑷX�/��4|B�O¡���xi$�z�xnU�H���U��sQw�M��t�������A�����㏯��,���^�g�uO`���
S�i7�8��U%���Kw��;�r���pgTp�_��d���I��fp�\���S��j��߹���WK�F|��^|Y�����ggI��n�C�+�Y��IC�a�aD�����\VD)�\FQ�^�Z�J�&��Q(�)ͯo�jp��4���Q��O�D*C�?�v¾��ڜ��:�1��g��Q�z�QF>�<�J!Y��xOC��X&^���8������[B=�O����삢fݳ�<��+#-eDdG��JW��z��p�u��#�z\s��� #B�=R��ņ:ec�|Q5#0��Z��vpʢ��0rOF۰��%j�.%��Q�V&l��/�������u���ޚ�`J��TPq��&�[�х�����0��wឩ�R�����P�#d&����T|���g���<����P]OB��Tq�qo�<��-/�ބ^V�[�h��0�M�
��og*ĥj��'X��G��7R��l�@<�q%��N�{!����� � �o��fX��ڈ:�I���� (����0<+@��Nc����M$���0����a��Ah{�ŋ�!_��v
wA��+�d�{��jjSa5J�ɂ��jR�??���?؊����Bǂ���,��|��c�n��ע�w�hѺ�l�N5d�N��_O����4|&���[�rw��T���)�h�=/u4p��i�=�8 (�����)��� �ɑԉ����b������B�<mo�4�������Q����I8t�D2���k�[d�;�����k������D�,d8@��V3e�Ez�^?�Z�}�/c�����>>���<�	��ڌ��n|[:�؍|�����{����<���o�bΈ�����e�(��� �!ka�;��.x��À���ia/��`P�mY&DR��nvWUV��7w���s�}/��hz#e���̌x��~�3~���4$�$s��`�Y,9h�r摣6L��*�� ��8���÷��sS��
��&c5�����HU�v���JP���C�@�2�+�H�z�ɋ��B�̽�_8 �$�g5�D�D(ȡi�Y�ś���u�X�(����p������v���fT��m������l��2�%f��Lo��=�u��Xzd Vb�Ҋro[�����0�s����L��	�@�9�Q5Z��[d��k�����<�,��YQ�6u+1���K�n�Ǌ�e���7�p��t~?50��b���h޶���,4`W<��>�#Z�(�����D��H�u@�:F���^�-���\	Ǿ������ �K���q>a���s�,�Gv�o<g��E���Z�j������dK�:����>�r��wq��d�����`W��BƷךmO�<��Y^^g�ꈂ�orVM�݁<�����%��[5���ٿ��{pit�X�w#9��SGξ��ج%M4�śu]�9zx_f�\�[��-�d!q�[��8���9�CiC����Ko�<3}N��X!�%ND�Z��T��l:�W�S����ز��V�T�;'K�C�1�k"��c-�7 ��;t˪5`*V\kTH�j�_ �*s��=�Id�;d�+��O��x����k��c�B���z(W7�$�ʱM��MV%Rh6�
6��@�]�U�U��j/Vy:+��4|"ҩ8>	��N��D��c#�V���J��ˠ9���V���p�S5�k��0��uz�sؗ��4�5��ʭF�;����������W�_���fD6�83����������!~�6
�ʙ�3���`��2/�oo4_��K��
/�Ucnկo^��HZF�x]Ve�,���V��\�QJx9���y���g�&�*�Txy�"<�Dcၕ��G�
���6��>���`Ca�#_���$3o�~.5�t.P�f#!�0[��T]��w~u%7�w���W�J�qL*-�eo�P�G�7�y��������8�@���4����q�k<֯����߉��E����
+s[�A�N3�֟��za�K�rC��&>�mX8e����8Z��ϏYcJ�K���h��D\FP�s&O  �������KoƐ���8؄Ff�,���LG|m��FD��+A 0���}q��y�Z��ںfr� N��������Gr���l�N:��qA����!ࣙ����xT`�E,o���8��*z�-�Y�E��[?�A���Wj�G�w���M̹D�>.������C>�|2�;��:�2 �����H5��˞�|���k��{�����ʍ�������qo�#��{�T;5Y\���j �Ԑ���1w퉬)�~G>y��c$w�W$�����y����_ߴ�hC�zqm�~��R�r1�e������ �W����x�8��u\Nl�~[��淋`Xq��1�z{E�g"V��ao=��b�(u{����G� ���k��g���T���<1�V�Mn~�/�Y��'��(�j�;>N۽�x�X���Q�5�g�	��C�� ?���ŸY$%Je���z����x.��M�G�(�܌)5�k�`�5J}��<���?ؓ���fkc9W�b�4i�'<_3Z%=%��1膠1ʬ����@2�ٰ��t���Aln���!ۜ\�ѿGњ
S�5���2J������@#X?ߑՖu���jH�L��޸l@se候n)��?���ʒ������Sn���`Tm �șlPf�x9+2.d�����?3.m��p^�O֐��[#��M Ԩ�0�u*����ls͜JW��J?o=��+}n����r���zn\��^���^�t� {A�gz��9��X�-H���X���ll�Q�N2�]^�'�Gj+�>y ��5�5�$J���^�͐,�N���2��oq�jIha�݋�z@W�C���>���bMc��4e�p_j����/�#c�+,�#K~d�|U��1���X {�,�z��mC�D�@�N����/�`5�o��0��g�>ݶ�ezc�8��0
�DVU)T�A����>K�Id�ZΞ�k ��P�G�!Y���g��Hj�ٚ�z+Ǔbcc8��>�A�+w`�Ű0�w<����O.����S�ەuB!��0k�g����J� s��1�!5o�k�-�g�[	k�.Y�8]X�m���p\7��P�,co�5�`2��k��wr�ྫྷ�>���2��c3��kT/�4]�w�;2�aOY��F^�+v�+bw��B��s�����c=�#���U樯g�|Y���nc�Е�I�JJ5�<��Ԗ�%3nأ��k��˯���g���u�T�>��  ���h[��q�w��_?x�������W��l�9������w����ɧr|�QY�鈒w5+�C�1��mI]�Z7�"�^ N��ֿ/ugb�v	 ����D���Ú-�~���E)ܡ�.�]��֓;͔)ZC��N�pt��^9����	���Q�N��rt���6�TǣW�qv�֗.J0�gx	]/Q�a�^����Ѧ�.������2���՗?+g�ˬ,�iY��Lx���Բ��绩�,Јb4U���od:�UYf���t�̀lX���#�F��Fջ]#������_7�0:-�y$U��$3�ln��g^�3�N�����q��J"nw\��QR깥�w<O�P�-B�LkP�:�6��1�}U����"bA��	�)l"B���p&�vW��"c��H�y�JR}-��5ҡؑW��amB�,Mqq���l�������C�IWDn_�ھC�Ye�b剪���!7K��QES���C@>sd�-�z��X��!��L�*胺a���P�-)*��v�"��d�Z@�[����ӽ�瀑�R$	=�f U�é��F� gV>f%g
qT!�����)�!x�,��Ae"B Vf�U��`CU�@Y[|(��	�t�贈�RXf��rߣt;������*#M$@`E[P�+�F������&�̖�C����m��f�9����R�XI�\jC`�=���~}��Q���F^�|\�>?�����,�
���C�y�ʣ��r˭:űѭצb��P�m?"��Z)'uX�ʍ�gˡ�'N�N;?��L� |�7-����Ky�����#�1cԐ���pak�D���������'���������;����������S:>	�.Lps*'x�֨8h�5Յ2G�6[ɢ�E7s�XK'�툌Rs��O�,Ԙh&�kJc�%'�JM3���}�\�������HG7N;ԥ��@H�M��\ qXs�
6�I����p,�
R�~r�?���%��ٻ�o�3��!�B��0ܟY��쓗�����߳:��*���R��ޢ^�2�Q���H^�⨪H�Ӕ�v�� 7FM�	`�I>r�O3���]�у����C�r$gN��{���0ov��{�^y��(�V����o!D-#����4�y���w;ƈ܆x"�ƂR�֘�tN��pP������hj�͞�G����[̨D��΢��wE#a�6+�̀����3zN�v;2�7������ ;��@�(19���5 ��kȜn3*��%�u펈��xI�G%!�����v���s��l��Ʋ����*�랴�T+$������;����wZ(�d����F��J���ē��p��RK�jdG�Cp=q�.%Z��;5w��V�!+OeV�3�^���Gg�����hD2BL�,�7���@Vdc�	�67:�\�f(����Na��t���j����?*s�L����-q �! ��**� P֜,*S�\��\_��2rT�8O49�`�90&�'0�=���˭f�cnyn:^�Fi܄�r)�`M��D^"ߋ$�	�
 ���hi ��h m��^��hiA���r0c��G��[����'cȲ�X�Ex��d_�Ft� �e6"D���Ec�������5�Dޞ*�?/���"e�M$�B�&���F���|8!fI= #V�����z�V��}����|�s���	��C��F�D0����.�����#­Lzs�5�
��]����̐��� ����eG���!ُv� ��N��F7*�(1��E�3�R���YL�Xf2�W�KS�hF �#A+55�P(�<�^���6��<r�_H�����@N�jlD��%a� ,7�>P�Dla�s�o���6=����a[�l(~��}�V���3/�{��3�,�2���|��`W�(���2Ǡ��~-��0�4puN4E��h��,V$�q�1�8C @��S�/�F���qY�R�8�@z1p�bP~�<"�Q�m�Ftʑ����,��d��5�@���3Y�G��n�-40���H4���:�mF6����ԉor:*�����c�F3
�
��pR���m�M��6$����>�<������Z1e[��Q��A�#s��S�λ��M��V�l�5�y������:!�����x��E)w4�I�m�*W6�Z�8Y�s�� ϒ�My�K��:�T�bC.�ˍ���s��|V#u�0�Ȉ��k�P�N8���D�E���އ���?&�����T�"��>F��P��g��t�lv�E5�a����+u�ׯ�@��4��	�zd;��� �4����PiI���`� Q��1� �e '=�kOV, X�������9 ~ge�mP-'��L6J��p��h�(ό�!����C��u0F�����H�؞k���b�x
�E��X&,�@��Z���U�օ@����$ЦĬQF~��$a|�w�z��N���FFw[��(�3��e���49���0{9��1(EW�j�R�?����^�V#���g_޿���~��{.���I8��%>�)u��\�wuq%��ʅ��-[=���z��h���0��4K�l1f�h����?��d)�gg2|~*�d%��#�f[��DF_��Dm5�uht�l�u1�M�,��Wj�IT+L�=��TBv�S$%�N:`վ���f=[�F��`�[�[�Ы��=�<��f��!��S��PC�H]����>2�y�^~&��u��}�})l����ӧ���	Z�!#:�:�bYp@���f���o�"s�`߇���`�M�os�6������P9bH�U7Ґ�9�2�@�^j�Yp6(�T�2T1J�Y(������Q��R���
���240?���Q0GͬJ] uɍeed|6�'�[iU38k�XK���ݥD`kS�*& 	:-8g���u>�uj�\���A�7���ԟ	�Cu�ٶ�j9 ���!P F��\.S���P_ �!ĵĄ������ %8�Օ�&�d� �|d���j�z�8"2g�`�^���9{� RH�f���Et��.6�ǀVO����2��ds����}�6��~�B�P��9]�Ń�&�DN
��Je�Ny���8���a�$�lkb$���T�����j���A�U��-ie#
\wO����K�2�ֆ���u=Yi�X��͛w���!S������%��J�%au1z=�M��@Y1�a�K0.	��c��5Ўŉzbb�f�|�D��P,h����}�]A{�NI_1u<��1�*}WH��r+��7~�ϞUTb��`{+�
 !V0cY��~J�zW��ŧ�j���$�.�����Pz/�Kx�����>ؓ�fu��$v����t!fp�����K)fwr��B���;]��/50hOs���ѱt4z���H��u�ęk9гy{�Vj�.!)Y,�h,����p�o��P^B`�h��8�3
v�(���c��u}'VĹ�s��q�����+䑕��A**����,�[�a =�ᢊ��#qJ�C�����0ud{�n�/�j��U���HD'��*��h�Yr��\�5��g�#>R��fF�C�f�a��1�KN�`'b��yUG9 ��|"��R��B���\]kFc!P�%�BJ���D&��Lf\Q�Կ��~���y���d(��qǯ�&P�Nt�����b}�R�E���hbhs2�٘���Y$���L����K���#��u`>�^�f�������ё���	[&g72)���(~ h ���$��\�_�X��D3ij��͒�qH���V�#Y���,�櫌#Iu��8�Q��C�#@��B*�@:T8h��U%��7��M,�� ��E�ebY�66h���n�d���c��8�p:7U;P���-.�S��Y�n�������Q�U�d-�:2=�kF6�7P��G�ljz"'>AK.<#S#���k� x�����~����G7RoY;h��y�=��S׿g���]I�[A�
��ب��`{ϑ[�[riX��Cp�ӽ1�/0���Ŵ�LOw�V{���,r,L�����Dj�S5H���i`��T��>�[��4X�=9����M���\^�c��8۫f3 �50J�����ߞ���?������B>���p�y�)�4�� �7t�)ɣ�Y��n,&��:�������Ǳ#��pl�,4rv]̠�K��G�eW3���7�C͂ j�l�H|1_��LMzu�2����)�W���t��9�M�y$F���a7�\�A ���UX�Y�#�I]jd�>� �WmW�*)T/S�5�-/Jp�l@rE�?���VN�G��2�ұ{����,������@��4�,��"�T��pf+�*�%^���D�!G<[}�%^7і3�<S$b��օ�0R�e-]Q��!�g���!��8�A�[��w#�Q^eA 2)�2�L��wwÊ������R��sV׫���I,��sC�����P��)���hx#+Lh���Lk>P&��	K�I���_��9�M��������-�3��j�{���;>���.�w�p_?��i �գ��F�͔x�D�g� �\}P��u�ز��x³֯B!� d`t܆���
Z� �&K����1.�3�Ȟ�W�ƶm����� �ҽ'+?�l-�2p*�a����F�S<��<�5US�-�Đg�Aj��s恕���Osk��R��F^�+ok�R�5���h�S�F1:]q��������%r����]
խ����}�"�1�N��2��*ȊN��V������*��"��5{R0�@V�1����Z�X'��o�v/���2P	JK�9�>B㠣�]ׄ� *5���x���ū�32�ȣǏ����ޛVG�S�z�/��k�;�����!��4�;�M�y��o���_���������[o�<>	���=5�
�іK����5��['���?�/� ���L��=~�X��G���?m��-��2_��G�3���.�������P��W_}��<%ب2�*A��t謺j�@�Qc��P��L�'a�~-�L��U�ޔ@�u�D��0��}�,*����l9�B��!�gurd�#M�x_Nu�>Ҿ)�}F�4�ۯ����1�A�Q�f8�0��H
�ۖ�����|��f�Y�w'nLtk�ڋ�g��{fN�eK���ym��˅
\7�4���9��U}vde�9.��@p�m�➾�!��=I�;4�S͊'�� �^/��x��S�
�B�#2)4����Ld�,AߔҢ��U�&��Y���*6n��_����b?y��r啤'�r���C};��m�D��F�����������;�%��5�{�P}��r�ꥬ�n��z?Fc��띨C%+Az��� ��<p>��&���#��5Y��@ J�ȉo�D�y�}��bm�тMRĹ��0�G�j�Q��� K��'�:�XPN�A��X̳jDf�;X�����
dVN�����b{��@�`K���RgFRC�Eq���@�®/�\V�XZ%+G1%��ɭt\X5�}zo�1��2 �
��1�D&��3n8u$X'_|����X�(ش���&1S��C[��Rr�	����g��@_ϣ��'36�o�b��)�<G��O5x^f�zX�-�k�Y��I���6BI��JG{V��ZM�7��F;�}M�:r��T?c�r��U[���=�j�m�c:����oj������?�'�����S�ĎO¡k�s)�,O�\sJD:�=!�yp,w����gg���L���K9;�A�-Gj<v�8� �RC�(�a:,�� �'����sp(χ����_��1�"J���4�ˡ�g��a,�Z���F���"�C�A�-�PS}�12Du��B�ԍ	�;2TKN���p���Cߞ�.<��������y}�K���q�E1��������ۯ�l���fZ���}jO���M�#v~���s(�jJ�M�ˇ�B�[Ubk��0���	Ø�:��� �I�^ZX?��>�O0M�h����+B�������pM�L��i �2J�di�>^�TeF���B�'2�& ��!v	ԁa�$D"6�[��Pg��L�d�s��f��E��233bjB�n��v�$aTJ,#�p������o��D���@�PEu�`
�������|�t�Ⱥ�X������\���hB�.�E��������}��ߓN�Cm�����u�A���+�%-.g�R�t��w��-@s���Hy@��j4�"Y)�Yqx{�~|m՝��mͦM#�J�tq9>Y��Z*j$s-�T�z���i��+'"&��uGJ�ܘ�hCBr�20�3��w����F�ya����DO�i�Ȱ+�n99 ��/��H����u��q�� hm=v
E�9�˓Ϟ�U�TF�!+$Ë�(�����x9��=�pX��ģh �����:p4[ܳ )�ڃ=U4L���)�BL�XF���T���83|��zb8p�����MXa�-������l���ܓ ��1��'�_�A�����n��/�����������C[�Ώ��$z��I9�����`��l	N^�h7���id�#��H&j|�.o���N��}�h�[�' �X ��(�o�}^�VO���q|yu'w���ӟw��.5c���y���ʾ��D%������RntsO1�BR��.�&?�:﹕���1�5QT�Vq��|���aql;�ʁG�{A ��=�^��B��?K��_��7��լ�ͅ�C-3Z�$߈�l��)���3F+��#�@-����=�pE��O��ͣ�=`b�F1Ia�� [�ݮ�?z���nv5���vV��İ�N����N#[k������v���Y�KN�$�CP�G��h��M@�(6�.�س $�ѱz�~�`���e:}$YH�����'j���'�`7��{]�銣�H�w��*�j�:z-�Nd_�{t�/d=�Tu}�z�N���;�ta����}|*��}��3?H���,t��Tg:ø�¤f5(����8���%�~�~|��c�,��m�%�IǍ��'�T@��K/d�ԧ��~�
%�g�c��rrL�m�{�l0�6�2���y�%pR,�%�Y?���~yQLY����v�.��"�M�xJl�DH/�q<��Ya���.��(y	��5x�B��i�\���dbO.0Q���ֹh& "<��޺g�����l�U�жncױ��U�s��"�Y)���X��2xنP�D�KN�md?�þ]�x�J���.V~������#�:{'C�=KN�tyOG�k:��~^-�خ#,��1�8f���d$�/_�����b[������e�$�:-Zs�]�I����׋h�H�v/gwա�t��/�so��6e���Z��N5����Ũ�B�,_�l�ᵛm�ٚt���$�ر���< i�$� �IM���Qs����, ך.	�[rQ��Nb���
�%R���`�R���̿G>��8'�a�,V�*���3���7T�ZlJ��%}3
����^��K�D��7���a�ѶP��N$���s�	,�%I�!�t�B�-2��M�ͬ>�a�	G���y�(}�ػf�����\7n��xō�R�R���K��^޵%��Kr<}]��3IO*̩�l78v���*{�K�X{@��(��!@0	f���@a�-��/�\j5O���Q3���[*5�	6� ����� ����|�$��k�������~9=�Y*�ATo��HmOX�z��w���/��?�0�Бu�9Lש\i�<o�:���C�� ew�|sc��8"B|_
�*�َH��3
��bmp����@�l]Q6	ִA���v�k~6� r��V�e�� ��Rh�5�K�h�F� n�Z�3��y�e��} 	f,��aRa��)P���)�F���.�6œX�j��ﷸ��E�e�?��-�Z�ؓ�@�TU;��Q��s�)�����HK��^wTS0��Ց�����m�U�!p�ZK)w2���y@ 
��<�sG�E�1G�<3'�ŗr��Tq!iQ� �V�
���U����х�50_`<�9cUl9������8756�C���
iVKIF�D05����Wѻ���р�?.�?���g�}2��C/�������d����k ��zB�ۑ.�;uȋۡ>�f�5�D|BJ҄J��u)_���X�R�>#�%�ܒ����78����{���ƺ1�,��g^���1Ѣ�کGҋ��C�P#Bv���.��	@!u���td��0�X��$()J�ss���:��}�JbЅ�fYO�M|�1{��	C��<E�(K��	&w�jF���t�Y�5�J�L�[�MaΘ�݅�IML�;�,	#HJ�QzVNu��qSX?��a�HC`�1vzU����Wd$3�!�Z��)�
W��%�e��PP��
A�ls ���Z�gs�I�7��@@�����
�[���BF�+��d|�6`�"c����k&Ӓ�N����ݭ��H��:u���ԵQ�V��͉Et�s��-���c'�	X��Ss�\;�R�#Hl����0�[�VITI��bW4�����1���\#�z�#��9w�����L�XB�F=i�B��y�w|�'�˽'���#�=< *�vr+�߾�ōRv��u;7�^�B�5�A/��z����&s�� �Չ7酄���.�wP��糥��-�7�B�>�/��C��"�z& ���t8:�N�;���W����B�58�11[�����сF}u9���j���� !	����(,WDO���o4#���kя1DP��u1�����x�\J9�VЏ[��:X�j 8���dJ�{Њs���8��ԀW�U���*I��|`+���4h�B����(����![e�sK�/36�Q"&Q�e��?״j{Q�8P�Y& ��$7�V?�@���9]�p�gu�3���:G��5�B���lS%hC�*hR�~RC��^��5)��V�Jj�k�Uh��Oh4���'�j�����G����?���w~g+"�8��Ρ�Ê޼yӸ=��`1���?����d�[�f;ā`���ꎛK��}qq*�'$��\�F��d�Ht��e�j�r����i1���%�t{/����e��;��!���������<�6aMѬQ�QxPC�\-O-��Id�y���@idY3F�<+��J�`�^U�ܥ����?h�v�HW����4��G?�y��U����D!����4v�Y�X�͖s��DaӨ%"�D3w�
vQ~n��s�r�Rͬ�g-��y���9��h]aHZM�~[�2�i ��� ��'�pb^w�-�K�����e:���k���এ�*�����,�����ul�2Ku6��kƊRF� ��~W��ZN߼�����������Su��,���ծ�z�n�-���g���@�'�dO�ju�W�D�:���3M+�r�X6e��7=/Hɭ�9J�k����:��ٜW'|�QJ���ẕ3qq\�C3����fЗ�No�5P4,������M9���w���`oG��$Ξ���/�����t����=�;���1���u�bb((K@����z u9W';��|t��~er���{��ٵ i����7/ə�R��=��w��K�]"�"`{,E�!̗r������Oexv!�o��Tx������������5���w����M�l���Z��]�ݓ�^�؝�s�R/�6���AbӟC�++�e���=�A�R.t�,��$�[(�g<ZEb�+��T@$)1+��`�� }X�.޼c����������>̠�R���2K/e�����>!M� ?�*�x+�9(6��tNnt�6�[�B"�maW]�J6w�;��q�^n��8�6��X�����u���D.p?���j�O�������M}�?0���Q9t�a����~��߽9?�צ���t9�����[5��f?���MI�A����_L4�K1��18�Z�c�9�4�e��0&Ȏ%�~�@7c��'��-�/��y,s]8�áF���r�r 7B�>2�j'���(B��*�@n	bu�K�sK�:�p�"
%�qy�%���l@���;�]�?y�Y�14����7�2�<����%;G�e��!�	y�S����Y��F����������W�6m���nb�����\�l�U�����4h�j�U�[�b������յ��9�tqE��C�
�O�q�^jN�ƙl�����d�,���i�li�_��D2J�A�)0��~1���#h��.d��2�����:�O2Fp踠��������Dv�١C�(V�9���Z2��%=�,#xf�ѵ<�Ɉo�C�e�-P��^|��L��3�Ih#DD9H�Ͻے|Ж��^� N0�]�zK����]Τ0�������[������ky���7_}�}�����@�X���y�Z��B��*���9����]�7�{�J��7r����1�@!kW��wKo����t�y���
������ĝ���<�H�D���+ ��y���{(W�?p���t,�ߗ�����_�
Ǡ��
�(���{�TXl�8��/W���W]�F�xrK}��W��G��M��.���w�]y/��K|?a����z�DeK���%���j�*�R9ёu.n�u�w}�R�������Y��=8�����;�(��-@e܈D[�(A�[m&*\iM�~ 1��\sѺV��X�]CLL���+S�l��0�N
$���;�M3���
��Uv�F63���WQ,��8?���}���v��N��~� ��ơ�
Ϟ=��޼y�߼~���n�����9�#Q��}������9Ӓ���Vsc6By��;X
M������k��s�����UG�PCߕ���(a����h���oLQ� m0h�^g��g�=+�x�ɢ���ys��<�k~�/�����P��ˣ�^��?��vҎ�G/dz}E|��c|��X��5���{�$`�~�̇����pP�m�؛wbeEd��͊65K �����XO��]=���f\��F�@xr�����N�G�f 稁��k�lj����{j�Y��2p�)L�$W"�����]�鳸>}+u��1h� ��bRk�58�r�
���xV`��%��
��T��#����2+��������FVөtbu:��l잙,m��O��wۣ���߷�����������/�7�,W@K�0��z9�,wG��Rc�z_�C}��/�����}�H��do����ٹ�?{.��su�/�1_KC?��D
�	�;fӇ�2=?g���9jG�  ��IDAT��u��{��Swu>Ԭ��AŮ:������A������+��N�� ���+r��o�r�~��7&�k��o�d9�����g�cm$�S�C�c�h�eO]��9z��:�����Y���&R��/2U3bDD8�s���׃'���^k�w�6O��V*z��,��,h���Y��r����m�S�g��y�tԏ1Ε�������=��E�΂S�nٗԪ�&�۽�ߏ݆��g3��X�_6���l���,�8�dթ��+B\9q)B�-��]���8�^�6�q5En�����ʩ;��Y"s
#G�����Y��'�׊4���7w�C����=�()b?���ŋ����߹���b�L����%�d��7�%�9P��\R@c	�)9yj%wqd��2d=i.��V�|2�86;�l������h&��+��@;�:���C�� 6J�0�;��]dnl�4�Б�0���=g�>��m�PD��.#T�՛�<�ɴF[ݢ������Fr�o�`O�vv�	5*�>hm#C�g2����|�]9���K�7�8Cقf<^l�0*�`���Mf3���:�4zق#W����A0i�%��A3׺�C�w:��@���j-͒��X����3W�N��z5��NG�D�q������� 3��U �~�X�o���z_�!��m�5�Y�렵+�*���F�˕L/@�����D�i!�G���+�����U���k��ω𾸸 qK����^7q��4��s�����e+����떣�UG�^���|����v��0tP5����<u�Gr��#u�=DFDM��ݥܪS?�k||�Y��eh��o_��ӟ�\.~�L�g�-�����a�S%0/_��}}y!�~�Sy��?��=d�POk��r���?Ҍ��#iI_�;��7�2�d{h y�nJ���@2u��Vp�fh���ݩ���k��[rܣ�*f�h�`� �D��w��{�P:J����K!�$�Yr$A&&7�y Z�z�kG�p�����+�FS����RTѐ��O�g�Q�Ԝ��1&�;hEj�~�#bhz���YFr�AQ��@�f��M��
/!�#o�"	�g�m>NZ�
�N���H,�gG��^	�ň�:K@��e��uk%���Ʃ�5��87^��Fܑ��y�ث
��j��3�JQ���c�Yg�ľs?�湷�ݹ��<C�e�1^y��W��������v>��������7~�7V��C�����_N��W�<��vB�"��4�b�ɊR��Pб�*�Ը��r��E]���ɀhF9-%M�?tL��Z�L���lԚ6��O���"�C��H�x�i�>�Ȓ�\����E�`�3Mb�hS/+�b�>�Zw�"GnG�8Uf��u�X�ư�(x8��ܲB+'���H�PJ�km��f��$kV�����q��xߝl��5����a�%��	�t�����9�|���	�Fro�չ�{]
���%Zl�$5,�D�~����up20���Iޒ�3~�$M_<v�cp��$)E@�k�m��@�F5�2�d<�'��l�}7S]s�=LJ�zD�J\7�W��^f4��b-K���13;ӠdZM(�i����"#T,�(!�Co�\�_r��������*tZ?1� A1	����E��D�_��:�vo��z��i�f����<|�T����˺۠�ե:���<��W/e1������a�RH
R��{۝%���7�̌�LrHk����ñ�@���'���F�%��C���IC�mvw���������:� *�޹:�O˃�~�{{=���s�j��
��`z��j`af��4p}��@?���C�)�ɛg����J.N��f�"�*�Ys!�d&��r�셮g+�B��ZL�@U���?<����a���������3v:��`�Ds��g<LH��g5�Y&��G�8ɒecb�G!��@h�϶`��@B�)� ���b�)nպ����6��_f�~2F3Q��
ERY��o �G��K<01�߂� ������2�
�PX% a�U?�9Q5M��r��H.��Nf�Y�6J�����?_����(���8�ɤ�V�Ɗ�ZJ���`�� ���e���eἾ�U]rV�%R��"��`�e��yG,�`�k�B�&B&���o���X�r˨�Հq	��rm�N�k��i��l����YȎQ��A	����2ZλcA-����{$Ռ'Uɜ~��P���Rˈ�%�� ��-u<u͚z�`�-
�����rtا�Y�nY�X,'�*@��{�V�*����n��q	��lf���ׁ��@�3�M��a�D1�3��# �nndJ]����q��P^J��c�~�V�dl_K��@����#���)Q��It��4���HsN@DgdY5�RmjU�ZҐ��Up���:�}0�Erx�����L3�KJ�.��������QrN`#��	�?�盝�U�
�����y^>�������o�hK2"��qVZ���CS��cu����!�h�^�f������r��#)Zu�˫Ky�򵮛��v���q����1����҄ib�N �eri���hcL+YV��ߙ�/�E�p�hTN��:�j��B�}���$h ��t�,��&g�k;m��̦��B7Q�ְj�J�E���]���}�	L����ϸ��![lC���3:��"����@=��h*�~���og\c����/7Nxlb1�����:�����(�����m����m�,�}b86;�y�6d3�$x��V���f���yU�.+W�	����37���J���2h����W�N�k��}����Y2��512)��ϫV���c�6�K�Y�[�=�*��T�yy��80���Ȧ�RJܨx48���� �n�77���gO��(�п�P��Y4���yi]'`+g	��QK͘�*EU��F���r�`Y���8'�F��`� �z�&P<�P� ���L͜?�f�	G!�Ο\1��!Bb4��š]]��2-5��KaF���z遣R�2��1�</�OCy�gQlz���M�h���j���@��.lC��Z�G[�x�a��%����ў���`�L�����.�nS�~xlGކe5���t�i�4��ԉ��5���d�Fs�E���cGϵ8��:`��hDr��3�z�; (i��9p(���L,��u�@��+�[@�a�D?�!��xi�۟�ĩo4�����/9θ�ٿ�)Ja�,'j7E!���h�@��៱TFm�^~�}.��z�~��[u��z��D,�\-SGGkЧ�p��H�>�X��:�뛡��z�'��}2bo/����R�h}�ﷸI�ZБ��\���ӬZ�E�0�Y�xa(i�8�zCZ}�>zp>$:�
f���9��¹ɱ�ж��`@��L}y܆VG��<�=]T#t�4 �L�s�� ��Y�9����9���;]9�챌�#�Ӏ�ju�m�b~�6��t;m��ԁ_�=e�=F�vQQ�6�;��eC 
��ܪ%IaԼtڶ<,Wɷ�gU7��p#����
f�Q�?����R����m�U�LUГ��>�t���B�\�~������M�p�t^�R�-���dS>��&�����I;*]L���r��"�APp����(�~���^V�y�5u˅ώ�lS�m"��AA̟k�3K~�h�F�����A��������q�=�..X.EO}�ӢyY'��.�U��c��Z� h�Jp��>���lKu����)���C�ԍ	�5ʌ�I�X@u����jx�RYA
׵�����]�o��`t��i��9Ɓ0���:ΞfnPU�\_��J�n,��Y2::1v9R3��A��ˊk�t���n@_������ �X��RW��֠/�nC�! �kʊ,V����5��b,Q�ə�)*��m0ަ��~���Xm�mvY�]�lYN�lBn�hD�SW��<�B��X��p^z���� ǉ,Y�l�UYƇ�!��H_���>�JxuVB�����#�X��A[�*�/odzv&2�;��2h66�d��*�k�ӱ��Ȅ={�W��ݨ3@�Q����Ǝ�<fF>+�Ί��E�Ȉt��AU�?K���C"����J�8"7d�QTF{��5�Cd�9��ݎ�|��t�\e5��Xbd�w�~G��B�ߜr�~�7����1h9{�J� ����GJ*��z�%OND����q�:=|�@zP������c��)�Y���e �s�21y�3C�cm��� /t��A����=8�\(�Fd����t/ ��֕��b��������+9:�'�O��ð�x�)?��q��vd������[@��B��#V�V�5�+��]9U�y ��� *.� P��x��Y����� ��e��Y��D�)#kۚv�,���HV�Qrz�Ϡ �6Yp�daM����|�|kd�Ė@�Ƒ_���h8�{�g���֢ۊ2�/K��.I�DX=S��F�\���Rqm���.��ϑ����(,Av Q�쁅��e9WF�`��Q���ՐR��80�����x6��ś�_��9t�5B��5�Bf���L,�D��<�����L��*v�W�g����X��z�QEt�B�2҆�P����bE�����2Q�f����}J͞��t � T�2=�f�p	'I}�~k\�UuUϨ�X����Z�Q�PJ&�νP�;T����LY�^�a��{��ԩ�G;2���I����˨�KI��_��Vs�����ݻ����(A(ޛ�B�
;>�1Z��B[���+u(��c6bY�x�^��]� :}������Uǌ�
Փ�dJ��=n �Z�ǯ�0�5&?��ϼ�\��3Y\���C`d�y��}���s�j2� K���1w�gά�Ԯm�����i�f�,r��o���@j�˽��aB�,��s��cͲ�G��ato���Z:\P�&�d>f���/^@3U4 �w|_��q	흁_��$�~��2C�c�z_��iG�+4+��+=������Su�G�tB�{��΀�l��暙��0*S���Յ3�:OW������;X�i`��J �f�)V	�B94��%i`[о����A�/�~�3y�_HP;����#�}�Tvwz�3���_��ߐ~��1m�$���ޯ����Wg��(䃱��\�vΔONҊx�Di��b��Hx���sJ�����K�ء�@�B� �=�
\V�lg�>��������e�L�]��3[Mrc�*{�y����+�vlg�e����wə�Η��M!�Y7�M����a=���+'Lj�3^e�m��׺fYΨ|lծ��"�H\r9D���2�/��Q1��^e��l�1��z_��C��C]�>�"]q��z�/�|��9�ɒ��0n�='���D7<R��:JHi�������%��&�Ջ�r���ݘ�W[�D�@Ҷ;�,�Xr����X���J�G�@58[[��D6��\�r�]�aA
%������ V�3T=*�Q�5)��0.'��_+j�����::P�rbd��z�X�G���o�X��tBC�QKn�\�t���e��C���l�%Ͽ�wsl�x&ؔ<����`�� ��� �1_�s�D�?�����-��-4�M�@�>��)�(}�P�!uJ�1�5ؚ��K��A�lT ����kH�Z��x����Tq�Ue^���ێ�pc�LՓ�l;�@������ʍ���mbQ��ۿ��,��S^��/x��{���vk�@���O>��<��j�1������_�O�'�9�ӆ�g$b��uY���K��@��?���otݯ�-�a�֪#5���Y��1 �H!�N3���fC�jr{v)�᝜�{#�}#����!��RzZ�5�!��3<(�ì�t߀�ջw�qJ;��e��U8x��X�+�ϗ_#mu����G2~�V���GC0q��'{ ���`J<@��v������ip��od�S؀�7Zu�t#�[��}b�{�)o� cc�<)��������C��KZ��)+NN���[;��@_�O�p�g���G�\b�2Br�zͿ\�e`P�Ըo���ꊿ\U�p�n��y��^�L#�3q�#;��}&��+L%�	�d���QgЉ�]��qB�Q����>y*��O5P��b
k?��[��I$�9��6��{���Q���Lߒ�b<��_�*��<>��z���E�&v@���f����*-tW�����		�:Hd�
���!��+.4�_��޽���ϹY��\���˳35(��y!
o�w[6Ρ��(��_Ĭ�������S'r�lN�S�- ����eǘ
����ii��L��~�L���7Y��$��ޡ�� ���0A3�5�}�~[���w�oe � �P2�si��o96���k�����~�J���Ƽդw��v���Kp����D �B��T&��LF2�l������� ��g���_�����x��Hl�w#�i���`0�D���H\V2��n�*99fz���%�0+&�.7�X�Q����7�AOV��/�+qQ��2�o1	����Gi�yQe�-Ѫ7	#m��B1��݁fǏ����N�2����y����;{r<PǦ����:~8�I�ے���������2���N���㌥�ȳ���7w���;}}�������r5��t*������gt��l(��A_��&B8�=m
j�o��!�&��J�w����Dn_��>~/8��f�9�-*+(�C�!�{����7�,�?�޽�o�������)�� 1J]8�'�˓'O���>��kr0��0�\���
}���n�o}=�s���|U�/�t�El�a�n�so�������6�����+�š�Q�Ի�(|������T���q9�\|F9�I:����¨�%߀��m�;�[ʑbk+`�?9�{��C�a7�����;�@���[N�U�����5]7�Ƶ;��4��1m��D?v~=$���vn�+L����&��H�� ����t��)��sF�¯�	>��q�Y�i#Z]3��7�� ���3]��7�@Ґ��p��qCWF��t9��]*��=2aq[�kD��Z��X�d��u5j�#�:��s�ʊ�U�e6�*�oD��4K�.�Z��%2�P��Y=4���c|��J��o)3��]�3��e/+[Z���g@V�5���G�z�$�k0���R����4��!#.w4��{����e�8d�/�6N��>����|�X`s1���9�m#u� �JW�vK�./��抔�<@ �>נ����c`;ݎ��S5�u�=��h��R��@��XL���Z&�D�d��/�����J�������r��Kd�j�Ni)�7m�|��
&c�� ����
�{���r��G����eп����G����	��o�����H�P+��}9���ޞ̠p��>��Y�-�LR���e��o��P���7FUY�Ѿ���3�ݏ�ø&������������?cƍl���C��4����9Z[P�Moe�ε�Ϫ�/�p�^c������ �v�<�d��kX���K4�k�|�>1g��:�zZ��%YM,�ڊ�^��Pn5����<O*Y�C;� =8M8��ɥ&Ky����{��iz:���c�5j5����9	����c��3@s�`J�Æ
Ikvi{0��R�@�����Tn 5;�YB�m���8e��F��>p���Q�@�PW�� �-U�#�>�Q�-İ��+"�r��$�E��2��=��|����_��/�=���nk��B|��g`�	bU��d����|�j��g����|�U�kϫ�5V
|��:���fhZ�,W5{]����_p��Rz��]�4�X��-L[i
SF¸�p���~\+4�ep���ǜ8��Xg��4�fЀ�U c+Y��Vǁ�"^K=��r٫�ľ\U���(������C��l�6p�b�Մ�@]@�� ��F���%��H��s�Gvn%�>+l�-!6B��B�'���⌼��V]�fd�=�U3��%�o:�˝�<�O��d,�(�e���9���l���ͩa�J0t�����5q�f��\4[[B0A�>�^�k3�z?�	~�s@�Ͻ�}����g�����J�ڸa`�",�# N�f�)�t!g�_��p"{7c� ���8:�*Wo_�6�U\4�,���s��ĺ������ґV�cS��|���ۑYϬ���/T�;�[��o��t~*c�W ����ddѢ@�.4����+_�6��k�S�~�=U�C��J[�R'���a>�#����1)��Wo��@{� �X��~�7���H��������;�]��2ۨ�p�����E�0
H���*,��ehgA[}��������qr�E�i�F�I��ب��t�)�}���>_]��o��~{G�9��z/�=�R�I^�~wdշ�:��<���lY\�|%�_=���5��jaX�²�C}����?>��i]�R��d4&��� �!PO؆vo|��[��0ެ���B��xO]*4�{cT�~�3+��ʇ	k�枙��a{��mO�A M�(<>��>���̷�u�a��R����$�uO�OQ����G���@���w��kX��Q�l B�o�Z(|?�Cg��ܛ�d5�{��sM�����G��c�'E��5�}�\R�c��`�Y/P�X�q�eer]	���OtP@*b")+����"6*�����ꝭ�2'!��b5_���e8� c�C�;�ll}}�ɁC}�΢��s�|�Һ���3�a�'�������cP���Y��ݙ[��;��+������t6��Z����w�2�l���
�ь�5������#ɍ#A+Н�^'�ra��(M	�������ۗ��b���bY[���D��E�zmK�qc��ɛ�S�����$��/E3�&�b�F�A޷�~J��O�#��&^n'yuq.��h/�����z���c��\į��k�r����/Q�F�#��7v@��*�l�W���۰�v��5�_��.���,�[B�Z�̉�h',k�Sg�&8�`��5� �,�7ᘂ��udK-�kw�]�v� ������6��Y<�8Q����}�.���,�ԡ�P7��Ǘg�63VV�9	˒<��X�U�N�;8���jv�d�k#�G�Ѩ�lS!	�}�G��& ��5*4�g�L�QH��ᘡֆ~{��6	Xd�kbf��G6��\I��'m�R퉮�ݮtIG����N�+z�$tj1�Xs���
��}��{�{�wt@p�����Y�&�b�2�󰊝��Y�ߪ՟E�V�����k���D<�*�* ���[��n��PyT � ���3�_d��'�Og2� �T�����~�o���i�7�[���S;^���ʕ���ծ��l��;]�eW?���r���RjC�rYf�M�F���B5��3�)C���%y�W��?7�q��$���Q&'��v�5����3v߆��nH��V^~E	�X�Ɔ��}O0�F�(g���k/gSfҽv���-�ðȦ�y 19����%��y��#I�/�s�������J�)I[X�L� 2
G�H���>�Ȍ������fi�m��*���>Og2� &����x-�9�HG#��� ��8��u+K��L�&�/�Ӽ�B}z�vk3���������,fF��`��|��\���L�~!�Ԯt���"%�� �{��S��#��:�4�X��� ��0�$\�F|���9g�k�%�U��B��V�m��� �g��K���>y�0�Q�*��Kረ�D�Μ�<�}*���Lg[���,=����Ab��j��+ �w�]�����1�9���(o4���=#�t��G��0���u��7��u�zw ;�����=ͦ�YS'�#��.�N3�/Gz)��Fhs*j�m�C̼�;���$Ӡ���Ci��r��F�Q�� ����Ҁ;����`C� 9�$��~��z�=9x�P:�@�{U��g��l��b�rb�sjV5 �k�b�;kJ�b8���ȕ�_F� ��p�,��&�B��7�etĘ�ii6��|8�%3�q ���P�I��7���F���1��w5��ʛׯ9�:�L5(�iO2�Ƿ�����	��%��ý_��U'W�c`_X��
���=���~���X��¦�Y%g���!��dn!�z~!�z��2�5���o��?��t�:L�/�j22�\1�/�<e>o�T6A�������p �mNv!.%X����=�ez�o�r��1��Z��Շ�7��S�hz-4	�C��$Ohح\ �C�/�;������;����0�JP��G'I��m�p���Y�u�:@��%a%�N��FĻ�{��۬���"��L�)0g��r��+yR�9�D��S.)x�K	2"�z�Ñ���2��fR������8[�<���/4Q�F�P�σ���d���\�
��ld� �Y�����_}C�@C��wI�� </��W&X�����I�mc���x	�-�ׯ�p�̡���˅^/�"{'���T��2��||�X��s��ݑ�]4`*qT��Y��;�~l��k�h�ς����A��v�ѫAQG�j
���V��&��$������mD�(��>���x���e���eV�LU�(4e���ǁCN,d��e�`���qc�(�1{�%6�t�px��<����s�Ou ���D��<��?���f�A�q[����C��Q��|����KIo'�O}�.�:�ӥ�k�`Ov�S���N�c_�u:r� �f ��AUg<ɻ��T�}!]u�Q�'z^{G��p��kd���LV���K��&�P�@�©���!�z��n+���P�|
�0�5��:�R��P9c۬�A��2<d�(N��?������n*rv*�w�kڭ�A���"��.��I7[��ڏ�<���H��K�vV2|y&ӻ�t��xr$ǿ��|.Xǫ�/�v2����gҍ���H����T~������7r�,�C(��^�K0����1���l��EYY�2��������" L"�0�o�U�A��)zϙ	O��CPp�Po*���,0R����
}���_���r��sr~�~�{�A��Grp��׷rs��f�6d��V#���W3i&m��w��܉c#L)���}ʪ�iZ��@���� �7үh]�۔Ep��&,P���)D�3����ơ�(����pla9_�a��`�R�7�H�}�tds6�d��-PŶ�]ң��}{{#/�yƬrG��r1�!pgo���`0��ZY�QZ�$��?�Ggb�F!W
)�@$+ �P]#ʧ��.����>���i$7 ��m�v�O2��\;�)���	gX%(�^鶠:��65$ �:]٫u���Xz��fc+����zk�����&K�\ǖ����s�9!�	� ������-��ڴ�Ho��sj������/Ԣ���c=� $�1y�ϣ���sT��G2A�*0J0�6ܫ��sp�'e�qKl���#�L��A��y��@8��,�_)7AB�0�Z�m�7�V_�����Ƞ��յ��2MNS/�������&�`��U_�'�mE�	[K9	��<䪡��H���4�+2�FƁ��k����˗rPWO��GZ���Y/b����k�7�n��GSAy51^��#[�GAr�UhZ#��/����{��)�196��;֬���!�����y �99?���������)N��t|��}9�FF�o��E�u6��������i�y'���e|s#�{Oc��V��lڹ�j������Ͽ'��?��'[0su��|��ߩ����?#��<A�2��ū琲d	3�ɟ�������$g�.O��_<z"-u� Ħ1cM�Vv��;��HZ�w���"A�B�{�	�Ց�A������ϥ���}�譣?���ը��]q�3��B��#J����z��tO���*R%�>F�ȓad3,�R�rƳ�yPV2#�'r��ˢ�8�E��{9�G#ڪ|��3R�Ʊ@����2&�73	ަ3څ��؉�7V�B�����
��������͝��N�K ̐�=�gOu��Ȋ�k�`#��5;��Рs����{�����������Z V
f�sI���{��Q-Lk��_'���:
ؚ��6cl������Qw:4���@0�2�7%V�!y�.�M�����rz_��z�3�+/�L-�xf\�}u�����P��bDf�^���!IӦ4��0s��D�@�c� �] ��)���u��|n�c��5�'x<��E{(y_��UK�X�R�є�<�|K�9v�A���V_�~�BV��e]y���\�|%��ȏo�)"E{ �gO�����A����R�������p:�p��7I�$�IX&Gy�lx��˒�j6[�kҎ��������P����3jwZ��k���zK��I3F�^0 �~&�|ӝ9���kڡܮ���מ3�>�u�2d�Gu�ƇʹX�}�#��#�����j��5���1�΍%�[N1��К$^:����=�@^�t�/�$���\�t)��?�Jbkc��L��Z�h`��%)y����x�Fo����X���ou�t���Q��fA1��͵L5�MW3ή߾{�ײ�����0��v�R��f$� �w~&���t�X�R"z�7�{����D���ȵ��.�{������^Ky��RjD��*�&[(
*^�Ad���&��2G�3Kc#~O6�8�F��6��ܭ,iwR���B��ITĐɣ��ҮG��zlO�찐��"?>��Q���"��f���=a�`�"#jm�J!!�mc��t�A<#�f�X�;���Ծ.��<��E>�|�g�F�GI�`��ޚ39�}K.e��aDۀ5%V�lm��އFh���5��q����{A�Y��ep�0�����^�Z�k����_�����WR�;��w�je�=�����\?<[Xic��{;E�������C��ӛT��և��j��![QSv"8h��tIT���3��@SD���X�U��t���+�*Bƾ"��,Fu>�ؠ<�$���)!D(�	@R���E��`�u��)zkj�&��zWi�����3�~'@y0������	�{����Y�r����Ⱥ�c���k< EIɋ�S�N�e���T��� ���I���ё�^����sz�~�)�f����f�8��k10a�\,�[`f���)=�  �)'q ��#��)��[��M0��Q�Ƒ����[t6_�i�g�&qf5��D���A����e����kJ-Ym�Ҿƞ�	ôlnB"���d�<�&�rb�X����l4�?���O�����oٟ�#��K����(��ũ���$� ��Y��/e�u�P��^��s��￑��-���z�S���r
�f���=g���8���������ˑ�gKi���g���j� '���v����d��DC ����V0��p���2X��ؓ��=	��Ɲ
(|I!�
c��%�aX��x�h��4�%�;�VR�I�ʡ3gOs�b~=��d,���&�!�Q�5�9뇧mݯm����&���J��9J�z-���8	����ف�؁�d�-c	<m�Z�@ú���&���e���\���_k�%Ϛ���ж�a�2��@�Q�4��ϑ5����6z���x/��A��Z�k�k�}HfP�{8�_Uؗ��@�d�2a�i���&�榑z����RG��5¬��-�{Fŝ_���+�?��d:��#L�j�6f,�G>�Cђ�d6��C��w����&7�U '1zj��PF�nf�;�,�f�g�2K�遦/oj�8.R',HĹ�Я�\gZ�r�Ty�_#�/g��.��S5�~��/��V4`Pϼ��0z �	�9�Ҏ���l5�AvQ-gYRk2������s:S���_QF�����L�=0��yo�Ցi���-Źm��څY�=���b$���R�_e&*��(��cqx�T�Kl� �&c|�W�n��[r>�	J�cU�����
,r�,���l��e!X��5��s��#�_b���tѼ5ҕ�3��a�o��Tz0��V~�̼�}9~������6�*�Z�k�}��R� �h�6z�zo�s�rlɾ��.4�}��/�q=�g�>����L_}If7��k"��	��c���t�cA���s�OK�|��0�~��~/G�P�TG��<�@@��"��b�]��M�4�HN�1�l��1��!��,��$nr�vL�l#�a�Tb���SD��������Q����� ����/�?{���˻;��=���"�N^�䏿;�������H�2������4�>d��1�7˟d�X����;Z@x^�
ͩ���@3�w���%tlI*{�\��U�*s���#���w+:W���?�L�V���&q-�.�Yr��-.5��`k� �V-�u�6�<��KZY�`�:q��2c�
�i VZr��
��g������r���ĵ� �q'��$�ɋ<�K��_J��0�r+�"Cg&�����G�	\h��ߦ��#ܣ�\ȣ�L�	
<l��ax8u̱3bM}��Ll;?���#9ctW��c��N��2�%�V�ER�yaA���>Ey��(�������Pj�H��{
@t����3��aܲ���z�Wz��b��Q��p�U7����u�C:���T�
�D�~��^?d	�p�&���%y���矱K+��;P�`ê��9�W����wҴ��Nހ����g�3J]	3���P��}- Y�mIְ6ެ�2u������#q�x�"�;sUa?܂u�=�����o���W����ʑ�_���A�4������͛,�5B�0�{�!>�@�̀�����H��Dn���H������J@;���C��b���e]�3�?�:FC��YՖ�3�Xd�1�b��)��}��z�ې�#��0_1�'y�>{���/�reń�|����>�$$�D@(�������@�60���剭Tw0![t1h�)
sj$�b��9�p���]]���?���F��n�l:Y΀4�ۖ�l�V���P��8�� '77l��?���teq?a�C;p�F(m��}�+*m@�ly!�N<��ځ��8��	,�� 8:����b\�r�62kX�fM�Xq[�q	�F�L�R��9�@Gᙚ��y�}�X�o�9�#0�������&� W�7�x��ҫ��'�wn�"��_���G���OΩ2]�p�N/��P�
>����;l'����(�C� =����e��|��[w��������:�7����(�Q���r� �h0���&�M���l��tJ'�f`�t�,X���tQ�B�ܵ��mhQRb/���&�;�4��3�
�=s�5��{�ސ|���َ{^���ՙ����}��J;X�?K�ht�8(Wс�+��8�E�	���ѫ��� Hh"^�ۗ��:�r�X���̑S�����(���|(�n�_�D&}j��4��m�A�.�hq1��dY+�h �K�SL�������Xz��`�
MԀ�fMx�������D`F�if�F�$R�3�ި�N���C���`��L
�w��dA3̵�hC p�?\����wt�3u�G�A���eŨ{�'����_���5ȇ=JZ�@���b�h��,h��R��n��Ub�;�!ة���p�kFB �e½���6s� �5 �t���RigI�(�#.݊l8��dv=��Φ2߳�;�X*��0[AxZi�m��Tڦ��r��wr��;�� ��e�ڵt��؃?� 3u�ؿ��{٪c����oGF��}��-Z#�O�*0��oץL3��Wt�M�(���ƌуD����H-P�*Pǀ,k`[d�m 5;(@t�y��� 1�FZ&�-K|D��q�:Nu���4��z�C�xTȠd�.$���&��&�"	���}S}�y�FY�>�D�A|Сό�/
��e���W�+����0YI�&��4ie>!��^�:����r��2r)6Yzmq��7�%ggg��"�?��4��@3���;�
s�p�eZ#�:���=c��h�mt�F��W0h|PaHYf't�2"
�h`T�z^Cu��y���g��h���Vu� ��R�N�:�`��p�| ;�B��Y��n����8�;��Ki=ک3�d��OPf���l��ux�x�j !��1�G�It.�����l%Q�5q��@�*E*���>�<���zt�46�Ęј�g~�;2�q������X��Z�s@/Ϙ�0�=V����8D�4k!�r����v^�?�f�#x�P��keQ��P!�΅� �5l��7�����2q���8�� ���f=��s��I��^����}#���Fs��fr<���g#Y���fG)z}�����G�}p���
��=� ,�)����fu!�`z�RNO��T�Im
5�]؃j�)��l ���q[���l�G������0[`Et?m�e�l���F�����\d� ���v����,''"z��^ۜs0`fNuBk�����F����du}K��D�T�9����*��[d�oՁOA:�%��C����+�{��=�t�������f3`�݊Hl��t't �fv�$s�=�R ���V�����D�O�sݶ�K�.M����-�ڀ#�'�k"Ϊ,��MǱ���栭EE��C8ZΩ()&��K�m��>� <��U��!o�p� ��� �9w�ZK��@��P��}�C0���l@Ԏ?���
h��|�a��p/5�?��dz�n��j��A���4Kl�3<(
��m�EJP*Æ���pX Ps=r|�}�:.�v��q/�n93�)d18��S:�bu���tT�rS������r�fE'җh+	l��L3�#�^��u�>ü,J�E[����%���F�!Ji���l�YԠӕVok�����,m�^T-��#u�00z)��T�gR5@�x���k9Wֲ��/xx&���F7ƻ�,;���;A �MN�Ǻ�s�C�ԉv~���m�f��㸎�_�:�I��hax�2�t�����=���P���61���u���(A�i]e��U{�ˏ6Q�b�T�qdq�%�*�sV'^]19Q[3��! ��"*IȊֳ�;���I�R���/2�fd~��*��E�Cg�#H�$8Qi��#,�r�!�>�3��f���@�]�ː��d^_�ۑf����\��Sf����P�8g�0-�&6�vK�ɓ'q^���g�/�2��,�_��~��l �A�%q�+2إ�E��*��ۉ�&����N�����g��Jju^������z:�>����#(�l�f\����$�.��	�K�`�2�'�0ʆv��[��[�O��ו�f�}}�p:����D:�ݤ�89b�QL��0���J�Qb1�_��h���		'h�h�JS�(mwZ������m=���]oP�[��O?J������:����+��1P�h�j���F��\΋��l�aOJL"�=�.k:�1X�4ؙ�5ߨ}~�i	F�۾\1��|yf|��)�����B��_ب_������:���6e�^�|m�����D�x��,�~�(��u�������x�5���	�~��k�ܢ������J:��8�l!�#��f��%�����MY�><"❽Ϊj�	��Vj Jg&�bs� ���:����6g��R�}[Y�����S-�q��0Kڀ�2�\�SU��a9��4�X3+Y��]���&��k�G��Y��F�w���$i���|c_>�yG0�g�o��
�c>���3��J�t�0�h`}0
���F��uS[k�G�c�6���6�C�m�7�R����@g�K��@��r���֣��+�*�H�X&@�v�xv���rt/�?�C�*[2ysmI��/��I�g�����%^��c���mMU��J�aUޅ�Lٳ�f� �Ķ�zd}�YQ�Y6�r��}$[]#��1	gΞ�$���ƽBKC_��koF�Z&惲;�"��T�ЂI��>�&3Lނʉ]�kl�>�g����2��P�x��.8j,-t�X%���� �}DA�)!�����~�4���p����V���u���<�8���?���������zd���ڮb�r�/c*��F+�4�5�����ldo����*��1DGV���E0·-�h5�EK�a$G�m���5��A&�Ouy{CY��b�kjE�*�W���C�s���;��T]o�N"xI5��G��7_K��T���o(C��Zh���۟���^n����I���ۏZk��%�sN={�H�?z���\��;�L��t�#�-|�\��g���}����O��d:��3��gı/,�
Gp�7��(�#�����9��v��	�@)5�}~2���Ƣ� ���[Jq&.�]i�I1����"e���4� �F�� ������r�A�62il��R6��з%7���#]�$^nShJq&�J�g�G��lxvj�X�C�07�'���@n��<�D�>����#W��V��F�3����o|�-?�K߬�ۃ��/��g^>(�Q��dgF�<H�!͒��qX�������x��w�Bm�s�|U�9�|	�5�w�yϐ�QpF�+��Х�`�#2lϠ�G�̮���^�����r��j2c`�A� �._�e��A�6�g�8�в���2=�8��^��� ��vz��d$��_�����ʘ��6���`HQ�^� =잜������-}�ǝu�_��\v=b[9���}T�<���-�in�!�sٱB�����1���X��^�_�wCE)���ަ�H[̾���5����:������<�z����"dŁ��n73��m	׊9Z��A~�AS$ua���_'ܓ������9��kY��й�ձ����F#���O��`��Y���T<�bk�����������S�F��7���}u�)T$�G$��{�	��9�Cڌ�53u��j��X�U���}���
mk��NlPm���f�p};���'��:�Ͼz-+]��7����2�Ͼ��'�������L[Aо"� C���!h�nc=��8?��|�k���_��ﾕ��FƗ5�P��R%��-�U�}B�]��C�k�:�W�;$�/���۾�-�)[ɯ��;ˠ�J,�iC0��z9U����Yo��0��%p����2Iy�����D�gD\��Q��֩q=c����d`z�b_��K��OS+�C�P����Jf��P��PL��~2���z1�LL��p�
Yi�	M�pPj�rS���*���؟�y���i�,f���@�&��>�rwD��< ���������:쵛�����q��tO���c��Sc�
M[e�<w�T��{�!��u!���1�Įp�av�`vwO�@�Gk?�B(�mm���Z�!��w.ȃ���V���F�S�(g����Y��U]�A>Xji�}����1so4����ZIk��3@�?�J@����\�]K3­9�Ǐd�)��>����V�g+�M�X�'��̸ p��![�LF���,�xVy�!X����X�B��RB/�)�����~B�=��cۥ� ��u R׮��eՠD��&�ܲ�X��:#`�"�{��d@��	���b(��`?C4��Z�03����L���k�h�Q����y0���)��|�w2u؋�p�V`���
z�5 h�Hn�}���܁�H���H�6pP�f}�:��<�&(�����(��%A���@'	p󅜡MC� ����YL�pt�m2}���Q'>�HJ�ڀ��rB��A�%O���峧����g?o�H3�N���L�Ў�gb��7`^�����z�f�CT�4�C�e�C���z����	��c]��G�I^�����G��Ѩp6_����
��̮j��}H���lOW������<�)Nb ��P���?8��M�> �{�F '�Nb����JCh2.252JU\��=%��Y�2S�.���[jv{�`M�	#7���'���Z\ȉS#��������ʩ}��Տ���~�͜��˚���t�����_I�w�"Aƽ8��&M?�@c%��yπ�@����߹ną�Cd�7�޼`b�=V���WW3�ǯ^��1E����K���c:ь#9���Y�JN1��5:7�����ft+��T�ܜU!J�jF��� ���}�$i�m�Y���
<��<��]|�~�6��Bm�1R���-g����ԙ�A���J�v�ӗ��\S�i��3u��z@5�$lc��|{�)�{���ܶ]�b� �=[�E���b�u�o"���!X���k˚���'���Z ��2`X�X���oI-��ɡ��=��D�B'��ql��ј6��1�E���j�ez��� ���Қ��vjZ��N�Y�^]˲W�`	�~�6`w{Ǟ=���]�Wr�.F�j�bƩN�؜{�bHPj���ğԜAP��4��������ڝ��k��w��u�%-�<�z�ПQ�6i���nM��1�'7��~Ʒ�x�gY��F���j�vw<#Mv����o��epr"}0�á���[�iӊ�|�� �9�-}��\hPm������:L��3�dq��J����ǜ|�UbR	���	9�:hD]��!�3��`8b)���~.7�Ñ�]�����G:��x�z!�=�쇟�y�N.�F�0�\GڽB��u���8"m�����:��`�ι���K�
ƽL%#3��VzO�0�w&4�o��9���5�<���d ���f���H%J띂<��m�2��p�@�R�$����/j����ݗ����9�\�xUZ��OL_8����Ơe�޺�H���ț�7{hbf<�L�=�/��[�ЎF?z�Kqdu$�����u��gf
�P�gi]��O1�/ �{'Gd	�^���vIgxR<���t�mu�^W�jL�1^S��}�w
m6Pޱ�ʝ䅍�@y��~<�	��S���x�̼ZI��Rh�wX��(�xV�Th���6�}��B"�L�W��:�^�M!̇#��!�O'2�O��^��~�N�5���V[6����ɝ$����U��3���^�%VTRg)s���Q犊ZЀ"u�S���{��R
=p��`��גiP�w�tB=Lg&�x���19��=�p��|��]KV�8�ad�m8��J��A�>�_��5�xO �iE���V��S���A��m?R�<q��%6A�޹U�,6�>�gQ9*I�1t���>�%��lt鐹ct@����}��������L��р�C� ڒ �����	���O��F��{�֘����)�H�2hbd!3��2V;)��������o����!�	��}�__�z>���w�.Z��'-��6������Rnn~���C�h�;0C{iJ�̱.����B�{88jF~"�;��=�Ƞ�.���ڸ����w��(�&d�����G|H�ɜ�tfd-*��joEH)>�ǈG�ӢRZ���3��wD�g޳j>'��0Jq��nh4�ݬF�����u��}��+� #$ �HZ��1���j$n���R��Y��n;
�*U��,����a��wgN�tWw*IOZ�n�J8�C�`�;f�V��q������ELU��`9� �ؼvD��q0�k���+Bee#����MQ�U�0��^-d��!�ݳc�,7j�PRD˃�b(5�GB� ���F��E�v�`::�?�vMɕ�+��I���ݗ�P����^����9�k^�E�^y�Db�đ�Đ�l�[XБ��i7��o��L�®�h�,W�,��6z_6�^����j�T�Q'ҕ��ф��R�;�DM�'Č�=m�ٺ�9�)�6� �0����tƠ����9�Ǘsu苙t�\{E�&�y��J�&N|G`�g�b�8��yj&p.bs����Ykr��:���W�5_Od�{z����Kف��(�ڢ�m9։�0�`��s���O�(�ӌk�㜑G��.�3��P_N"���)T�R��'��-����f{}f�mjX�8���hQFҭ�Q`6�dS�l��/e<����N�ɂ3��څr[IO��q�/�\�6|;]H� �Z7�L���6�L�K���*\��Soo�*v���w�����R>��q��jP���鞇�r���R����)��W�U�Ń�<�0mQ�`��˵F姧��k,�=�t�$� �d�ł2�N������ei����4��e���xm(��&�ۑ�MD�c"-�@=G��Ԇ���F������i^�mp�К�9Ge N��AJbcb$�P�4Q�q�iʎ=[5���n+��qь�l."��{�1�8��/D�������lgV&Lxm���Ԝj�sU�:d�b�0��X>޳��+1C�)�r���U�,miS��Y'����@$by����F\���X�[h������{�܌�0����k9R��^�SE�܌-f��Ѫ��1��{:m�
�.Υ���+�f��  
�C�;���i��)e/�X�C��Iڂ���J�|�7@�s3=�_Ӭ� @�K�"��S6��$���/�nd�����cl�vF�C��"D�c^XI�を� f�p/�Cd��{�Y����:��d�- �C�k h1�Yv�n�z�W R��1�ŞR�S����L�pꛍ]��:7�X`jօ^#��%����`���=�99]�l��������{(R#��4Z>r[?��b��@I'ao�9 �ٻ�9,��FO�Yc���(�pA����0�
BU�E[h�z�'q7~h$eq_1��Y�����g)3{�v��_6��Ʒ��n��N�N�h*�%�K[�B�f��nbdJ��U`�������R�r��tV㊎�n�Aڴ%	-�M@����d�?w`b#)��� 
A��D(-A��FC��^���{`z�Y��w?���S���X��E 9QH��ա#j� P�ù���j�MQl�>��h��`s�q�2�����J�,�f�f��2�c<d&r]o=���	+`�{�#8,�G��g��]�s��"��[�Ut����W.8�6��b���T�q�Hv8��f�l@��Ү��
 pR��$�ш� Ep���k�>7#��½�rUj"��bMd�b�n� ��QzL����w>�
�^���(��|(Z�$��*�O��ab�,�^,ث�lY�	'��������f���yp*�y:B<ô��j~�ja6��h|u#��{�߹G���N�]JW��]"��;]Ow��6|����ɹ\�x!=�6�\��|#u�(�"���sO��e��Rz��Glbd�v�2d��-��}�4)8�{"�w����&� �(V���ǘx���������%��s�D�:�z#	�~���տ��(ͼ�X��k&��~�l�^��U��W_1��sO�+�ee�m���� x��X�����ͪ!���I�ԪfIE�v��^<y.��+a"8������RSg9l�gQ8(wNwT���W/�DfNbT�z����m/��ץ܏&zz�,5��.�R�Sq����P{�����\�[/{-`�Z��R���G�2o1���jQ�7 �AU��1��^$�-+G%�,�E;�m��*�O�9���Y� �;���`�&qQ�z��<���{=��ڄ`L�3����t�c���J��D�e��X�	��G�ST�>е�qQ�e� 2��x"���S��ʆ�Sp���v�$d>L����C]�/Aa��0��!"��*�0񨊋���zC4D�t������X��߰ߕ��ǜ���X�Y�����|Ε:������(}n�-���b &2q�.�0��3�z�z ����82��=��˹f�+�q���h=����9��KY���\<{&GO.$�s�NZ���.N%]o�{<��g�IG�Tm��J�q�Hv=��Oz7[H5Nx��b�����a{G����Sk��Fרe!.�N[���@�.�L��Ď$O��({��;�fЩ�v���dN���'�)�s���E\H��r?G_P��$Nd� ���NQT�L9O��x�t���߃�l��&�z5���J���TF��!HBI0��
�PW]���_�����e=,d��nt��~&��X��5���ez}�$&3S��9�̊F4�z���Ǹ��i�������ZڿcP1���A�#p�HjҴ�ȎbO`������L�hT��	���uǃ�o�l�C�u��נ����f��+�ٍ��f-�W#���@��"Q�9��؆5�XP��VQ�	��ǜ����k�@��s H��y(��R��D�K��O�l����}.�u��pJ@��\k�焾vɪ�&,[���n�gM���-��<Q���*Kb=D�p(�>3�	l��Jj�ƒ�xB;��}ꠀ�����; ���y��`�������q�cr��{��ƒ/�ޏ�bb��yp� >ѐ��n$��s�{jc�XpX�0jH0���B�T��A��$dA�b]"F(�qG�1{ű@�4M�Oׅ>�P���75V+|^�9JG`��,9�	�����@��C'�R�pQpI��14�A����gr~<Јw���J_�}9Sg�a��|,��fc�ހ���Ԉ����^�ڌzƇ�F��.!p�El.�;)X�`&�(��zr�A��D�b��W���D�r#�02�v#���AR�?�\ɽF�A��W��I��c֔(Ϟ�꾒�ɭ�8k��2��&�H6z`Wjg����M�2q��C�(A�6�|!�$�����	QX�k�I;ۂ�~f���Z������Q ء|�m؃��D�@m=M�-�
�z.����α�>荙S�^b��2�G��#*<sJ��ٺ�S'�_������#}q�\�~�J�_|F��
:�+�����HG���D�N*�ѩf�k��|S�L��d�������G���3��dԡD�C��奌����5*&n[y��C��s�1�~���I��u�ܳ}�/~S�"ܩ�R�k�#c�r?`�ِ97�~ł��UHKZ�����; H�/�#��B,@bF4����˶��7E�Z��X�w^& *p�o5xȑՋ;8<?1V�(��#��!���m��bG#�ؾ@�ZY��\��&n�0��������ı�����A"�]�\y�N	b1���V�j;o@�1���e��c+�܃�H�2q$���Yݻ;����z$�v ',��x*��t8:������I�1�D����X�� 1���:�3�y�5���Hr���B�o�Ae:���!a� �� ,�V<���L̂ۈ��^o�y����� 5���Ej��O��t�p�rd`�H����FX��C0Q8y���\X���n\��zO:pb�lԡ#���ry��TN@6��46>@ZX ��:��.$�M7�19�����3 �Şt��G�� cH� L&�á�x�D�P�z�РO"��u!�(�MX�q]l����>2��`(.cd���5�4�N��*+g��Tۦ�@!��D�Q�H�_�hUj�`�a�l%,��r�QW_ҙ�$�(=a��:j#z��i��fN9��񦟛Z<��K�| ������vP�%�A�������7��g!��%w��Ѷh�;N���|�d oO�]�ڡ'}7R��� ���wd$��)Q�E���*I�m��uPb�_�����N���������w�@��U�=���Y![�zH��1�A�3��Zޙ�$�e{N��ǱRP���a����+0��I�Q���֐�/��D���ٿ����:{���vI���.D�Ǿ,�jG�d@��[��7�Ld�&��I��� W�iV�ں�pU�Hb^��g�lQ�U=��z� 	I�۸X�y�^_*]C`.[�����&^u#�"�9o޻�(w��<O6�d0>����g-�R��m��uJ#�I)lR���ü�z%[�\]�L�棱&;V����;ŏ覲?i �Ĭ$�Arh�Y��ǣ�VD<����FXf���XۤB�ϸ����ܹY2a[�2B��H��RUO"�8��g�?ך���v���P��^��'�����CF��xpV[>��$2��P�ψ�v��
�M��R��U|�)���f$t�f�"���aW���f?{+��[�q~��2��ve�м�Jy�-{�hr��`f�J���|�>�`��`e��ʚ�{G<���x�̇���57J[� z̷��r���⳧�ż��5�!��K�=���r��`ÏGt�y�C�3��b� ټ-����o��Һ1켽"p��4����?�s<�IOS�3c���g,�%�EQ�`�R�W	Q��C����C�~���Pe�u�^�˦FfJmBX��~/*<����Ȏ�K��!/G����)eˍ7%G}?�z����ߏ���5��^����+�=��=	������T�(I�Vǧ���P�>��r$w�[:���Ȏ��g�֚o:�S�	���cI'/��!��/�_d?~�C1*�$�&6�R7��Q1�2&+Z�W�`lmf���sfV�j�X�� �cy������U�}�4�^�����9˜���6a�u�Ħ���@b+US����Nxfs�,�RM�'h�ٯ�,�a~�w9�-ܯ=��ܙ'^�7涚6%�޻J��_&X�h���i.]�(�*�#�5'��%�������ȸ; 0p�$���<� (}2s�y���Rڰ	 �����l"˛k�_��5�4���84�e�6��C�8V���zk/V<8��f=6�9be{V;c��V�I�q	��Q�<�8xɠ��Uf��)[C^
��-���?�mڃ��4���~����x������'p|2%w�rCAf���D��d���6cb���*�e5����m�g9��l�d�aLD���~��35�fP��>Ǉf����2���Cp^�D��������=[T�_��G�Q�+&������ё���ʰ?��,�[�ʕ�mȘ�ʥ7� ����??SG=���Ϟ�FX�I����Hn��,�G3x�~�5��m��L<���#Ә��`��q��E��ɳ����#jk�߽���l��]��jC�7��V�bY� ��ˇ�D|��Igf��p���d���&MI�~��jd$�?$�y	2�6.��2sZ��F��_����,�#�-WLe�����k��[n���J����{P�ơ�`uzU�.H�/�~wM8��"9����{#N�_/�TIv$*1ǘa�L�aMg7h��D/��d���6�����l21��-eF��"s.�8��h��
J��t��=þ��uP�<�h��/�8[�yOu3գ��,�$�Rqߦ���F��@�ΪR�|�����,RW��.��
���g��g��uK��������K�8pꣂ="�f=�Vmƻ��ޱ�s�j�_'���4*�л۝�0A����C]�]������F��F�ņ���G�Sn���g�I�O��x^܏"�$p\c��"���c��<���-���zں��.P_!!�d�$#���V�;�=i�z�;�ڵ�/�H��n�3�W1�0�BN<�*��蟎C�3_�Jͭ'��X���9����M���S�ͯ�b�63L��d��V��G���t�ь3�Ȍ0l���=�<(=�K'n���6%.,�H�o� c�/��xH,e��=����e��v1�������A_��:��>��!N��a��.�g �K��^�'�̈́r��ɉA������ә����>�w���t�Η�!"gR�]� S_� |x~z*O�O��l(���e�#zUVs�nɂ��"����lkN�b�����R{����f����m��S(���T��G�T�aY=4�kV9h����÷>����A�tX�Ј� ߁V��c�; �9�3��a������#�����D�FPä���"C ����9�`��%�4,4����c��pf�o�����%F�`�F��q.I���1ʵ�k�S��������C��<����a�����{�辭8F��\ϲW5��Y�9~��Lp�A�����!�Vn�X�I�pT���<���i\O��`�jq�4�,���J���}Xz��#��!j�\8�f�>�M�-i��!a�=@.��gѮ�()�9>,p[HH��)Sg�sMpؒJҭ���$�ɍ����zCz"�@%	r��在v�`� ���t,����4�i����˼�+[q�6��Z��dK2IyX�8�� ��t���N�_��VőU�Ɉ�R&�JU=�9��b�<�AG�^hL�bb�� ��^�"�<�M����-�_�������m�|��<����f�v�r���/��NU�S'�H�_<�D�ʚ�������&Hc�t�h|O-k����f�kR.F����ix�<�>�[5���)�	)/��8bH˹f�s���ù����.$>�����k ����,�L-3ݬ�; �"�6�Ybn�E��P9i��q��sTt$;�Y��h��,���Yɬ�4s٩��Р�&a�\������L./s�����г=
6�PeV�gT�T��hm�Ȓ�Ԕ�`�r�����z♕7!��TH� �k�ײ/+c����uR�����5q�f<s��Kk�@���рi��=I��Z6r$dk���Yʻ����n����x� J�+��k�e��B�:�a:� ��8�|f%]T�H<=�4�X<,e:�u�l�!�}��[+��Q)�A� �V����eX���[�j.ٛ�M(cgҭh�,�������K=��ɔ���xWN��{��2v�(����f��sF����}�A6�s���I��s��b*d�1S'��%q`d�
b%�ㄞ��S�¡�`��T;2YMe���!v6�78{�����z��x��9����Ef�d�6����W�����_��{�ٔ���-uߢ�V��F�*���N�b��z\1��b��I>��	z)h�r��޶�]����S]�F{������/ɼ�j&nS-b�ǥif๞��8���Y�)�`�r��p�5�7��1�|03V��E�sY8���� (������Cׇ�̗j���Lg����=�:�.sU��=[,`;��`�52!���kA���&�rO�b�q2��m֥�i���U}�(ڝ�p��Ac%qn�҈T���z���bI$�a��WA)�jn$8���4{����z'S='̯�a��~n�ȿ���C�=���S�r��l�������7����ޔ�]���N����6smR�V�2���F��~j��U�G'g
�����l� �is�7Yk����x5�5��i�[�DX������Zil���K��i(Y!�=�j�K�b-�����AG�����c,�Ͼ'�ݜZ�F,����,C�L��n�&J���:�^K��L�R�����T��+K`"�9�	,�&���zc|� ]�݇B��s�2��~�i������%T~��6��)�n���Á�<~,G��t�u?:=�w�?��O�h [�	q0�� G�?�4�Q=����X�)�¨�} �?>W\};#>��"#0q������kɚgg�~�2�����gx?8�ʫ9�v�HHT�/H�Z�%������Xn�����wk��\m�
�� �AmM�;z�u�`4dD���ĳ����?9��d�57��4�^I�%�Z7՚6$��K�����2�P�
4V�Wƀ��m�W�U�+\���209\�����뫭�C�e댂h)F�iq���������&��IH(�g��	I諗�9[�ļ��+��9��j���l��e��ȿ��e=����W�� � ث�9`߃'κ�f���ߪ��:�>_��&���(��)JZ����̣!o�\��'����:܎�a��X/�jdBPU�!�7s�f�1n�����9��n�e�;;R$��#঄���n��N̵����6zC�E�XG�9�K�k�ɶ)���w�b>��P>�Ej6���7kc�YT72mN�Rs�;�̪n����Y��=xQaw+;�>Rg�Q"n��"���ٔlz� 1;�r]�+3��y�1ζ��4�rDؒ�H�Q.��������g���m��5��@cg�����i�}�$.A�L��"�)����I԰���eGL"����1����"�Un�:K"v�&�zŁF������y|�ch���|���yiߪ�(��S	�=���W
2���mX�AP�~oI"#��}]q4�Hq��R�_+�^[���놁[��	gs\c���<��_|!�Ʒ�W2�NY����s����[t��ZRǼ%��c��kG���4{� Ȇ{�Y����5uURX�z�9 (Qف�![�u9N�����=ӄ�P�7&��y�ppJ�>���C������.�s`��<z�k)�?��}M�VM�8~6ڂyj�y|Fo �ֵ����$>��i�_g�7� �:�����+:�3�ד)�P�3�� Du��%(41�h}��J<ƅ�gȼ	�0�fp"��밶ՖltݠZ���y��jG�r{}C�
9]V�t�ZCFI�h�&>g�Z-�9H�&��U5��Ցo�g���BW���t�O��Xc�α1�B-�OR����mY`��+��em9����@��|ɀ�K h9`�D����G�۫�L��� �z�@ớ��j�%}�I�?!��Nw����鄣T XdD=WT���T�An���> '��B�h�ܸG�ߓ���E�������I#3���᎗�S#N���\$3�4��kVYR��rd�;���
�qd�$�� �6�(��$��̀iD�C�Y7�C�1!�7�2S�s��gh���-q�<����o���^��`C�g�e�3�&H��񍤹w�U|�LY�wҥ�U��a鹫sm�-��������|���)�i�BRrZ!!�t��9�q*�!՚�x*��9)���Q7�D;�;�MG �E~|ޗ}������� �|е�=��;o��S�����Xňs�|�����;ꀈqBv���c�����0#i	�0��XK!�ml�B$�͖� �(���=��:��Q"���؉��5>��(b�B5@2/�nP�i;���"�ɉ���l��c�I�8����&ȷ��WTVi3���~/�U�抡��85�Q������Ed����M�dA���),[���@� !T�!��>V�V��{�8yV�<�l�8	R �'4��+a͊~"K�] ���N&]�7�w��QUS��9J�&��D��D��X�,m˲N�J���:C�M��4�Xj?x�`.9x��r�I��\f|�t��#*Q���T��}�HF`�C�EϷt=���AW��J���)[hx����۷�H��>�*�bسuK���^�Q����L���׵Ug�5y��h���#bUvD���?q"�-�� )@UkЕG����[2�ұV���0����+�ǧ\k �Y�����v�U�V���>I���8�gϞ-_�z��u��o��w��ֆ�Q���2c�`#	�&o�gR˱|'I�f��Ґ�g|k����bi�n9�B���V�-*��6`���Ш.1�hQ.z���E����gγl�	��6��އG�+��bF&�T�e�,�\�s3҈���iS]��N��q6�A8��O�y�ME"5�;�'s����!t��(o[�;K��s��!��3i�$�IA�1E�}�
d�F�=�V��w3�0�XZ�*A9��U�<� 4�z뀗���P��10Ì7�0Udۚ+]-���W����d���0���X�; $��p!�A�VD2��mY��e�˱*G��ܴ�Bhf�P�|���`H�,5�N�]��g��\Ǭ�`�	D=����)�Qp�8>���o����_8�'K@�g�F��/�`R������#ـXG��x�y����xh���zt������ŉ�����U�"��h�'?�9J����1�QqU��:T��RbU#rx��*3��J�ȕ�8U�Q췳�G� B7����@ɚZ+s�U�+�<��x��Zh��� uC������8���H3kϹtW
�I��e�����o��D$��s�#z�6+�Wj�o��gsc�Ipn����?������c��Ao��  ��;�dGx��f�K�-$(��Ԧ��V`�<?��pH[��7���[��Z�Ԩ+�=���S�ࣻ�H�Y�<J�F������5
,k@�?��|��j�2�]�n3	��Ak��i��o����!L[��?Yk��+X�9~�#pI����q�'�ɔl��鷬:։=����%˶�	��C��/���?�����dxs7��a�|�N⹬��$�W(��L��2T'TtZ�<ȖU;�\�� 31PDJŝ��iV�Ϫ����%m+�'0 ]] �C�^�JX����D&��\�9@9$w��2:�T܈��@OD��L'�\|GYΊYSe�4� ����?�@�t?�i���g��sU�7읓]����K��\��H�����}�?����EW�Ot���=�L73X�-��
(F�d���r6g�+���8N�p>�=?���Fȕ�܎��O�2_,�ZL�m�B7+�S>{|!��=f����\��˚dNB�Z�QБs����9O��rws'�Iuc#��B�9���"���BQ</NYx%
[����/I\g��֌HC�����w��ޟ��a�l�e�ί> �I���	Ugj�Z
>��_`�c6�gϠ�n�}�=�A��.�`H���Q�Mu?�'z/5�Z�z6V�=0�jfdEh% ��IRt��p����03�UYƃ�g�C֛���_f�w��	��R��L���@�q�2[x�J��:��f�Y �}����,�/��B�P�t�'՟M�G)��z�⎊ל�xu���Ϳ}�B���4�����^C�d ��y,����d����@�ܖ[�u�Ff���
�'��LzE� ra�J�4�}m����7#���J��o�wD�#h.����n�i{�Cjel�E��'v�1w�1�.!������X)��H�V���]y������Z&!��G�hF��x<�n�/}8q0�a�x���\�|%��9�)�����4�\�>_z���iq��2V�����dZ�
��Q��6!�e{��9�~�Z���ӥ|��'��q����I��t}���I��ϫ����}���_�?Y܍�W�ܥ�aa�{r,]��|��%��+3��՚���R#E-�fM��z���R�P�Gg�tR2�����J6���q�%���f�Qއ[,눟2`ʮp^0��I�L*x��)9�촩L����]7���5A#y�a��_9�)�oK-�����)���z�����(dR)F�c@��'� ��}z,�Ԩ3��ʇ]y񛯥�������ٗڦz�v�l����E�)t�5xѿy���N����'���Y�C��;Y��� ~	��y;�G�����^�o�k���9����y�	Xэ�����/_|�\^�~�,�'�+� �Y��a�C %JQ�F�,����S��+�t�v�0qA3nr^�`f {�:7��&����fiHh�j8�\������j�5��F`PC� q�0���9������ܸ���ۇ}���>��}X*NM(�y��I<G���#B@�'��huZ4���#*N��T5ǱZ Ɓ�+7�!�i�����*1G���
�S�-@�`�2@('1*��ZX�~��Q��5��wpr�=��7���;F������L�N�����AXVZ��MaЪ&֮O��(���xF�����@�ʸܫ&8��b��ݝ�`��L�E�f�5@����u�0��6/ML��
N���<}xx����ϝ���V���%�"f���޿��;��2��I���[@.v'��#���� ���k�l�>�s8??��f��_G�kR��P���ׯ�ݛ��۷��od��I��I�I�r�sc��Cdk'Ë3y��� ��§�V�����dC^��\]_����|��7 k�*�� �7���,�[�-�Kb�`��g�k���J��B>��r�8���k�o�5����L�_e����Knr�� ����]-�>-��[��oF#AIl6�K}3]t]�����>�/:N֒��}��$���ׯ�����4*<{�^^�ß���ŵ��ȉ�D�� >=�4#2�S�`�#�想]9�6��PVĜ,�y0�u��~��G%�`ԐA�C��t�!(���kB�l���˩� ��+�C��Uz-�̽!I�s-�<��8�����$#�o�>�yt-�c͆GsLWҾ��^���:��=����eΆr�J�_�Ѡ�l���B(*M�ך��^^ 5X]uj����DГ+�E�JLj}�^ԏ]9Ѭ��������/��w�pz���ץ(�ΐ٠�	�3�,�}�O�6>`Ы����^m7��1{��w��ϟ?���a2C�2���L6����c�	�=s$���eI0�-fKYk�3��:Q�ZI�{��</�G<�ϊ��Cp������@�Դ�����;L( `	�l}Nk`,w��e��?��j�(�w�R��ɉ����iS*
��x�Ӏ�o'��E®��0`��~)�'H�T�᣽t3���]d�1C�]��z�Y�l�h����p+oSFՆ�r�σ�9>��޾�$��4�����i:$Xqn�	X?��^�1�E�F�tma¥E�7!TG��*8�>�K���\�J �T�P�J� %��5���%@��]��{�s����a�xp�6%3�"�d�>���[�ߡ���s�}^c�,thg�݃G���Jj2�X?���ޗ&�bא�����g~.������Z��Sf�d�D]Am�?}��BY���l���y��m�PM��[f�k@�Z�_E�g����^�noe9��=����A� �]��>ħ2]u:�����8vg�Tcx��Zku�)���(0�/���r�F�ɣ��g��)iF�ys��hDG��#����A�7��@���!�H��/?%�^!?ޏ��=Ɇ�⦣���Uþ�if�R����u�(cLh`tBЁ,�=�ܐP�6b	̾g�B�l	R�k�vk�^��ks�	A1;70��������O�9 � ��21רj�gw13�:�fյ����	�V Ŕ功�jzw���F��B7�>����\�_��K���z!@�񮆸���:�S�"�P��f�G���#����U��v	���+S9�z���j�N�';U��T�����������} -���@�x�\n�+��Fg�����޶9��h��cr���4���`Ʋ,��48����f�в�3�������@���Wz�gr=�Hy3����LJ�D2���x V����O_|&g�_
V��f3��Hż\���n�l�Z���җ7�<���ulip�'��u���zl�O�*h��p�&!hH,�����@Q���zZ-�7Q��e��+�(n�w.[S������>u m��$��:�T%u�����E��s�-*(9�e혡��A2��r9gy||Ld6^.d�vm\��{�)���E���H��Qz6�
O��4QM��-!z5�SR�|�-��Ҧ=�P���>�
��;`@������ct���Ȭ�b{�"">4 :��Q�ПBv�Ѭ��|;��q�l�xj��#6��1*�@�k6��=�釢[4��^���%跱n��z���tϏ58�m��&��d.��Ff�EC짧�������ז�bf��Y����=:=���#hs�%�s�뾻���� ]���:���2�ܱ���k<�g0P[�J��V�|U%I]~X��$�Oڡ��U{=]lG�es����Ӎfy��Bҳ�G�F�����4ʾ���hC�TN��d���?ֿ�
��Q�lk�6��Ṝ�8Ѭs��#S���1�l>ׅ��Kz7kK~7�!��8�]q�b�_ �$��^P�I3 Dx�b�fS`N?�D����\3 �Z�iNr�3o+�t�'1D�`�t ���_2��JY�j��ߏ2k����#�8��͚�>��߰����(���Q-"��l�e�;�#sݕS5���/ü+��|w���n���9�A�:{,Ǻ�.tCw�z�ר����8>|.�Ϟit�d�H�e��Zn�\�fls���9�O����������-�-�� �i��)t�,?�\Fb����R�	����x�Y�l��67p�X���T�F�v֚�����pl*�^~�ՠj#'�����ic�H��}y/�M�A^ƾ2�<�!P��L^Vk��S9~�������͍fS����[;�Ej�}|�n*�OZ1��Qd_r�L��9������)�X1K�?nއ��b�xQ/���F���
���v�ऺ�)�{�&���څ��^)#�) u����W'4h[ Sm��i�����> (���yH�~o�P��zA���	�86�������fo�'N���=�+�M�ݘaO�5��nzi���eȸ}pl %�$����κƱw㨣9��l����)�����u/����3[��Z˚�f��+RC����j����M�� x���ö]�8#hgp�6�A��G��<}�TN�>������V�=&_��k��iPz{})����G����?|�5��ݏrs=2����^N��$ �P�����M&����w�>>��ׯ5��\���k�R�|s}�g�_ߛF9�Fw�a��� ��6N��D�~�%�ל��ӷ�ʷ߾�������|>���ڱ��!|�A@�Gjz �Rېc�-��'�+�i;�d�-S�5��<�� X�YU�@���)u�\�-Ͳ�u��øwKR��:SMT&�.�'�#;kq�h�=7�H�n�Z�̷��{b��jp{�1�Є&�y�HI�7�V�D���jH0ϛ��Ĝ&�$���]],1�8)��:#����X�2w����{�9+w�8�c�93H�.�r�+-Cw ��cN2"�A��,�Y�5x8����r��&�$Y�ts�ՠ�*�>��(��^"��j�y}y��d;��{��S�����H.��`mu�1���U#�6xO1C�`��R�A5��4�A��0��0���g��=�+���@�FL->�#2�T��4���56�/*9~�x�F򽎌����:�9���g�$ّ$h�I�OZ��A8̜���9�?��`vnvf���J�;;S��<"vvjE@JveFz8yϨ�jo �T(��o�!`�y���\P=-O3�z]�]Jz�Y���ب8�p�=����b�q�"&�,��}�菀q-áwv�B�GL�%��SfJh�ɴh ���ڏ��c ���>�)���*J���2@f�f��~��ѣN���<I��N�zGɤ`�xP�ZT�{5�Ȅ���0�y���9�yRy��!W1�Y�{ow��~z�O�iv������a����S�s��͵��� L�xx \	ʇ�7�ǣ�4JL� �� ��9�RW��~�S~�|��0(�激��0�g�d3�3��a#Ȋ|��P�P(GVE!�s1}u���ٳgry���`$�Ʉ�B�5���5��Z�cv3�gQ�D+i��S����P黗�|+݋sy��\\H�B�|A`� Lŵ'�=�Z�bD
Pm�VPx�.62���F��d6�;�P��m?W��N���unY=�9��Aɮ��9�"H �8:�Y��/��E;t��(b�e"%f{��n��&�4����Z���H�Ǯ.��q5�ojv�OrTFO�+�5�qƓ/s�[���� �YO�L7�z|z�t칲��*&�����٘2k^�gQM+��
U��v08 9�C��Lv�%pd��w�-!6i�",17�dm��c1��{��¡Vzg���lH�PK��&���o�f ��܏�	�ߩ)����B.k5���E��8. ���j!�-���;2�L���l*w�w�<�Z�=��k6�8F�`p�3]'�O�ua$=����f�Ձ�4�����[�ڣaE���t��؊�a v  G��gx�7�LO�nR��?Bɜm���4Au���%�/Y��nl�R���ߧ`E�Xϋe�nG"���z}�� ĩ7x �����܁� �DX$@���=�Aml<'Hj֑gx�jxafǹ6Ӯ)x�5ʛ��mΞja^�"nj?coSi��!�z�1����r,����V>�����Ӈ3�J`&�#9%}�[Ê�����)�ly{Nv�i+J+sD�h=9�Pw��$K��� ^<X@���o<�A:�b�쾓�Zc%"�s��5�s �P�����C�q �.p)X�L�6g�D�e]��*F6�CQ9���Z���/@��q	��x}��`%޹������&�+�4���p�6��@Y�7�����PF�޺��cs�<�`��~6N��[)7�(�,��U�u��.����)�u��\����>#��`f�Yp���#�԰��~�Y�G�����}��$o����*���
|����ƒ?�"hg4~���T{�w����\a�'���8��XDJ�И�����Rv��֘+GT��L�Eԡ�1I��	&���O({u0o�cԑ񂗘�.d�\�Z�̵:r�\_����Q� �>ʹ�/ɑ�Qg�z8���ϒ+y b̉��h��`���6I�RZGO�^Cdm�"��d�.���a�(�`��B��^Ɠ	��.>�j?!D?��R:��,��dYX	�������X~�3�4�Ef����]�L >B���[��PHO*���Guިp�)5K�cX�6:���@ ;��Qu��s�Z.��$�O�sA0����V���nFP�NL�Ρ�ҥ�/����;���A�(W�� p���M�H�AC�2pj�Ud�_Kp���L�O�g��gO9��r������յ��.�^q7ΌJ���hz��w����(7�=���?�mmޙSk��H�d2��6�﯒G���ޗ���ҙXcu�1u���5gK�2e/�A�؀o����w<ΣE�[����g$3�d
�^y,>
ĐC��)�}Q��.�㍙'�	s�p ���I�S���/|	��y�I��3�X���f�d�����N��?�'Ǯ��WP*bX���#��.:�s�A����"'@X����$�����03�����<�=�jj��&"��hP_��̧��p�6hi+�`�x��D�L��b-iᨈY�W�/��ѡ��a���`HL)}��參�������@�&Oԡ�lN��s$��s�2)��ǉ|�ye����&!w~�}�db�X�H2�@m�`�3)a��{��D���{�o~E�I��a�a	��pT2�	��n�<����~7���3�S���������d+ ��M[}�gp�9D���Gc�1}}}Ͳ�k�Y_ Bd��:��SE�{�NJ�{���R����Acz� ���:fE�qW,�#��x@��=G8�Ҡq��䛮���L�~�
��Z��S9E� +æs&��	�X�O;�,���r|g6څ����kH-<�U^(��������z�9�:��}��>��l��fŌ�s\k4,�6?���`D�<�g|��ݬ�W���f���b��صF��Jk@�B���X���t� z��!(Y�Qֶ�{�fڄ�AU�2����̱��6��<��`�"�/��˙y]<�G�V'^C�jz�a*�?�&�y�����?�,r��]��R�f�VdM���$�6��GT[l3�u;JՔ�O��9㱦^�3d�A�&̌T���.��ڜ��O��g����z�`r��;��"�	��l2��V&%�fl8��y�#���g���l=z���C&u ���w���ޙ�S.Q�&{���V�6��Ү�l�{p�Ԗ��9~z��ԁ3��@V�L�5q�{�2�,4[7Z���W�zR��<9~���"�9����(�Ll]�l߲r=d�3��c������I�C��r
�B��;�y�? ��:�v{y_T�+���W���<p��۸S��tϢ�"�?�jo�r��`�����6�9,fc�X��z�I!ŷ$�e�^q����	���L�IF��Z�=�TLR0k�$��L�C|8�3�__�CGGLox�T&N�Yד�'�bsy{+��Wr�������ӫKr������t-}M����Ǐ��q��5�B(�T[c�W0�20:���_}#�Ȍtq�5
}vv�~��~����˺	�����ͮ�{ׅ5��2�@���x�ؗ�aRR���C(��J�1dp2h�\p3�:��I `��X�3��4Vbg�ٍ'�a��&	��t�jfKLd g$�f�EMp���奫���ً8�{�t�{�-:�1���d��p�w岗��p �4[�Py��9�`�B����,�k�-��/'H�������ځ@��Ѕ��N�Ec�����9����d���[�4;_�\7�a��}CK����k��s=�X3;����*ȝB1l��gz`����n�b����e����k"$�L7��k�:�~�Fzz/�ӅL�]�R/ײ�L������o_3��7_1[���=�"�tԉMond�F-��Ե� )�Tlb�ٜˮ���lV�Y.$5��+s>�xbx�{$�t$y�A6��<�l��	2��Ͻ�٘�M�	�ډfw����j����I�Bˊ%�8Ψ�@j�n$[�)p�k �윣cq�:0�'�2�˪�\ ~#��NӸޅe����~j�c_	��5P?��������? �O��B�ݪ^Ǳ����ARd��m����@���4d��J�gX�C(ٲ9�[x� ���v�!�4����?��|�cRD�`i�M|�a���P���o���VM�m|������4A&���#��G����Gv�H����І��|,o�������|�N����L4@�+(l��mm�)�N�~|NX��`$���_˫�/���X���A�=�)Y�5�Y:�3@8�0<��+��ş�"���@����Й�WV
��:���̀���^f�?H�<��ǻ��~���Aܑ�(�G#jHts��M�-��F39����J>ܾ�ɿ���-4���A�ޢ����-�uM�����z)�nN����al����r�����7��Pa|�O���h��L��$��H�fr��^��ƿ�0�JX��Xň��uΦ��@�tZ\K��\�njmp�[�^�rPd$M���bl[����&KsY;0���f��FJ��e�k�����:����;:�J���z=����zz=̍o7��we�қ��L7`,�{Kb�#<���W�#[Ƽ��������1������s�֏�,���y	pИ�=�V�Õ��n~�O��kqW�Rh�шx���>�aڕ��R�{� �3���A35�z#,jGFl��f�������N���T��J��D��V��]��^�F�ȾG�>8�e����t�kU�E]���D���
����L`��_����� ��������S�����=��~�w�9gذP�����)�uמ�X|o����E{�U���)�Ms�Q[�>�-��Zee�^�H��3��X�W���s�?�pl�~O8:�u@�cm���߇`��.�k�HY�<����ޱ�as)FO~��O3�������֦Q�%r�t �Ӂ�h���{��Y|�O	���c:��Xu�Z*�9&c���}D�S8s2qF�
��f��|��!~�����%1�اp���6!S'��5*�L�0��L�p�5�		�5��(c���7���N���L4i�X �q�ĮU���p�H�=��sm;A x���I}�q7�� ��� �B0����_m���G��/��E;tW�*Ա��MC87,��!�L��xK��F���5�:w���2��W�3���yWb��8�\���.����.�o%;ԆyȞ�G���$K�X��;9'�N�+�|
�n�iF����Z���$��=3��b��mL���no$��_����F�nw���9�D��2�f���>x�._��Ci+�������eKg��ړo�R*�c��%���oi#M�T��g �����3=_����g=��N� �5k��H�׺9.(�i@�F����x<>����4_�Yl^o2��;I���R@���q� 1�������A;b��{�����\����ܥ�#N����h�u��8a���J{/^��b$[}&3��@E�L#���@F�0z���93�@�g�q-��u�sT1��y?~�Y�5Qe�<��+T8'v�w������C��� ?����N��=�Z�ާzO�NG�M44&�۵V���ھ!�L�a�L���FIcxO^j%�B��'_U��T���wLD�'���z�� �Y͑+��22��78� ȋBi؅����(�+5�g�;�^eFylf8n�R�d�a�^�lghO�|���fZޕ������G伵3�Aȩ�>���}8	^�S�k��x,�����\q�YW�Y��m&�棵V5���&?۴�r'�鬍�QJ�w<�ez=�#��5J気�b��g�8�3�8UH$��v���z�TK϶���f�$����tod��
���gp�}��z�vI�ap���݈��>�����l�[���Bբ��|�@�l��xJ��hdՑ�PI�L�V����~�p��@ۡ�\�&�Rz�&�3r'���_N3�r��1�J`N"���7~���'�J�ݖ�5��桗]+�dþ�_���3Y��2^�:�?~P�?���Q=�F��	�L�:��s��������}�����wG2�z��]�h0$�D�\����P��f�::
�s�18�>zE�e�z�q�F:�$��G�Q����Y�S����P��Q���m��8�2Do��Mj���($c6�K���M��+�A�V�o�$i���c�T޽�`�x�3����ɹ3<���5�?���� W�鞝˳�s����h�ܿ���L�ܲr��sF�A�蘁@�g�dp�ϟ?w1�D����72���H��K�W������;.�&�]�0���A":���7i!_�#Y���{��9� �މ5hC6���A���ч)�@-��\��3f�)˞��h#���a���P�ҍl�z����~�ZzÑܾ�kr�`-��PZUqK��z��HL��*1�1#�k8&Tx�T/$�H�8�1Vrc��V�>f7�\�������#����-�������/�q3HX|����Ҏ�g�������5
�em:p��4����|��4���9�q�1	�3 ��c�ӏ���Y���<��5����B�FdKȪ�x�e����E`���U�a.����[��GH|����	�hc����	�<Xy��N''�����k1�;C��%���DA.�ܐ6�rШ�a�@w0��_��J����J�zM�YOm�f�h����t�N��w��V�/��l)�=&>rc�8���{������dQ�-���	?�I�+�-�G.��d�� >�����(ۘ��`�$4ݎ#@ׯ��(�|��/ڡ�N�0�6�}��fb)�q��FՉ2���$@o��L��JY"��md��B.^�K�YO�n�~��|$�.�%�0�P���d���1�]�B ��Fȫ74��ټi	F:�|�L25�yޗD��#5�e��6�GA������e�f�-�IU�$]�L�ﳫkq4���Ys&>�*�x��ob�%}b�eP!O0G���iY"�8�K��uM(�h%�c|����'�6�t���ip�\.x_.�� x/;���$C��,���N7&Ю=��{#YO3�~O�Þ���^n���	u�%L-�3jZo�(�S�	�G2��N�|�Z��od�?�T��]j�9�4D۪�[`d̥2ן�WGRhp4V��� ����ʺ��5��F H<8nh`�N/�$���0�C��]��	��}��A���[��t�4�� 0��:� ����D#�{���zm�TB���-��`i�&���+.��M��y��Mq���6@V6m؀�J�TE��Гw��;�Vr���{��&��y:�֢��#?7mY��U��8�����	}d��W�B��J��l��@u�����a����d���OK��"�?��O�io�t.����pf�.��e�'b���>�Z�q)�
��r�!ڍ#��5�-��i% ��Wζ#co|e���2���_�	���@�k#�����t�T��W��\\=���~CY���Z~���ɰw)��3��kҠ{yn��/6���F��A~\,��v��n�Gɀ8q^J�a�j��ȯ���O�2�jЏ ��c�Ӊ[S�� �&٘����ܓC�������
Uw�|}���G��y���O��u.e��P$�?D�І�7V�F�Pr�p��RV�R�����}��o��OA��5�Nֳ��u��=e_��~)a��X{4+�|G�>f��.�S��ru��:=G�_ҍ���"ug��"���4*�k�s=��ك,���8?��F2�b��,�2#��x��� g S6�&��(�i/#�`��g �VȀ���Ԝ�Шz�Q��v�񏡞{�z��v#�~�q�,*�������^�����l"7%�3� �+�>ʀ���@����̘�!*�_�me)�n����^>,r��8��q���\��k#�I�������;�q>���H�N*ϯ�2�L�F��f�y�B�z� �8�:` ���a�ރᐨ��z��27�<�!VMG#b��F�����������j�fd33ӂ�.��2&�����F�b�!�#�+�[U�R=�g�2�u2�w6!ad*�����{�D����y��O�ٜ:ۧ��j$Vj���kx�M����	b��a�ÜN���$ek�u|sԔ����{��w�H�G�t|����a�e�]O����>1������/m��Ϸ�Z"s��
�UA@��2�o�:m��>�%(�5�,�2�=L��aygN�>� Og���SD��~���p���Xk o�^V{g�����n2������2��+Yk�4|��y��N���ג��+��S��Ӆ��5�� >%����#�{6�ʫ痒hP���y�@҄c�)t�A�م,>�仂�ɼ*��%�Q
�pK�e��h���V���7�\�J�ثp�[o��tC7�UsP��M�^,J��<<N���� �P���9����d+�Łz���h�"`H�&f�O��A��7�8�$�诀ҏ�Hq�����7S �.���%G$L���"Uk��q";=�{�'��k��+�%y�Ԡ�z���9K�.�1��+"��������9���y���A[�|}��y�hS2%g�c��~�^H��ffF# i��h��X���8���ד; ��x�.@0�f�B]�4C�w��7y������J0�>��dnI��ۛ��g�΍� �H�r������aW��Ų�t�V3r�JLN%q���{��s;0~�@����;5�$h�X���۸Y��hP���n���&��B�k�H��;i3ؘڳ1��J��ʱ�D��ɶ9��gD*�n�Z�BC5;Β�:��Bj,!n����1��	|�C)�̆k��dLӺ��9����RtFZ��>��5s0\���G~|��k�8W������f.�0jf�ՀTu}���e��|O��OqG���N�^N Z���I���@fw{xߏ�8�"� @!p����m��/�L���Ǻ��<�)].*N(�׾ZG�9������i���W�J�փ��������(�E�Ǘ�/?�f2[��7S�<�$>�e�A��jɶ��^h���W��ՠ/��'Ii~kW6�z��V��y���z��i���f 'q+Rꦤ��t�˽�������e���P�VC�%h&NJ�__�C�Ă0z �a��5�Y���P B�A`R��9�s	��cJ8�_������$�4j�8���L&w3Y-��BM��T�،mBD�x�G+��4�@+~䰧X�J3�Nґ�f��@+ �D|&���W��.��L5d�@�2��=�&ƌ�X~��F:gT�B
h��u�i�	�Q�Sg�W���	* ��K<	��T�>CVM����@�u؄�(^����,����i/����7չ`����
kt#)�Yl%�g�7y���z�;��w���!:�R٨�� ��p����e�\I����V��X_���љM �č�O�6 �l�A��D6��@�y��F�4�ݽ�{���w�p#�mI��Z�HzCY[��f��yc���`*�l��>��������\�PCW[�ÀEȸ�h�T�Mܾ}��5�����=N+˄y�8�}ݚξ��c�Io���eN�W+�����V�5�R�Γq�*��m>�r�~�1I;^����>��E��}vo��ȫ}����_}g?�ئD!{���Io�O�NK�ra}D�ȟBN�f��g���'h����i`p��&���JԼ6�+?�UDkN�$�@A�	V��"�l*�N�#��-��V�#�^���=T�a��~t���y ۧ9��1O��2D�?|F���w&1�-@n���jϞ��ݫ�܂x��l�����ݍw�%� =�K2}Fᜭ:r��YS��L�x�
^81篃k8��`���� 7��ε�A��E1x��>ȦKP��* �D$���Lҿh��W����NHq�5�ڠ��YA0w�����g�\�6Q?��1��l����Fa�������6J�M��o'�#��f��mB��Q'�ȼ��Dr��:a�ڍ��0�8��Y����b���9!:�X�T3��:pn0���Z��4&���aO��-����@$施���$v)�:�~��:���v���x S@���g��1��j�v�u㙐�J��������iZ���"�د��w���/V&���q��g�7�\v !�Z#�jR?���N�fI�WG��`��!����y��AD7:_�l68��U84�⢙�9���;�%��H�d�IRz1�����ߑ����T�-�,�����ٙ\�h���xuq������e�p'�r%��+���������d�,���)L��*�>XR#S�������	�`?,�r�CA�Z�9cNX�4ɈL�W�^�exǱ�&8���.M�T��[�<&O���)-�BI�Pꎼ�%3y"�w<�Iy�v�j�#r�|X~tx>3�ѧe�'���Ϧ}�e��ש=u�͟�����OG�Nz럖���&��l��z�`��KT
��V{���l��o"r�@����W<���43�l����vN/#��#�Q�Nﴭ��\J �1�
������z�;��V���'lI���Ku�H<4 0�
;�P���L�&������5|�8�MQ�5q�ߤ�k���J�~��/\�r6'�g���<��9l)x/���Nj������L� �5c�r(�&Ҁ��=���L\�ι�Jrz�0 L��U�z��ŎP�Gqq�gr+�z}.�3�CF�7��Ǜ������(�YID~^� f����H�#� �H�9ew{�B3Ĭ��\��-��:b�����~-+ݨ�������+Jo���$:����B&�����w��7�v�O/��A�F���P2V�%��ȶC�9Ъn��5�XSG��K��5>��J�4(���'���7k�������k�]�*[�����HOJ����u��3��2����}+�5�uY���y�r.&{ȇ�XЄ
W��߼QЍ�D- A�9��t-�w�����{z_5`��v��Yn��=�<F3�D7��潞��^^?�A/��/_�����H����`����ad}��t昸HIL�C�� �T�ǩ�A=��KP��[v�a�1���D3����e-BU��h�"#WiX}�
L���mHRD�{ρo(&�BF�x��x2_�`W�6"��8F�eb����[`����L�3��Q�:_�ʒ'\B@|�����D��΂���v�����~�[��{{��X�q|�� 0�?<9��'�PZ*��ec�D��T��#�e0�e�X,o�<Ɓ`P1}�$267:�Ґ��� �S��4�n|�'o�~�T��~t���P	5z��W���:Ϩ�^p�j@��e��S8��$	G`�>� �gٸ?��Z��ԏ��Bo�������5���6��R7�����X����.��hvUL^k)���}gb� ظ�dGRMO��������8���j�{����8Ki�]Tj{k��;6F=���S� u��8���րpi0�ҘF��6Y�����መE�2����N�w0���������	S�(���3�[]`@����%��K܉�0

�e���F�wL'�4��������z>P2����mB,^FB���<](�{p�m�X�O��L:R��y�l܏�jo3��_f\
!��t9�J���A;�VK�6]4f%Ns�4�v���E?4�� �Z0��r���5���B���.�x���_n��ƵB�I��U��t96�6zmt�5ؘiЕԙ���g�7���1ы�X�4,�9cI�zޠ��TV���\ݸ��G,�[Η�1d�T�"���:d����i�ڂ��~���<�>����S|�O�s�V7t���7����>;b�̽���i�
��eE�����F*W??ʡR�T����	��[�7�R7�W�lK0�h�ЗwBtsR�>͢����t�M��_c�<#1y
�:�Qo꧟wZ��pY�����W�Uפa�0�c��g4�`a�\>+�U.�ɛ~{���*���n�j�ʠk��c���|��^	��=��p��믮�[����IG���MCVp���-�F��t�EXz���z���/)�^�P��~M��#�N�A�#`*ڪnc�(Ώ�oA?[��;�߭c?�o�&��W؛^Ů�=�k��#ûڴ#=�*�l'�?��E;���8��S�;S��s�b��F�$���q��Xٮe���*2m7s��n*��Ր�������Gu(@Q��8�6�����XJz���0>�R��f)�ل�񢫋mRqვ,�E:�{�F2��'^aʺY��m(X2�vdM�f��%q��s��t�:/0im7��/�s�˃��l�������(�l2��G]����� ��ld�f/���p�>�!�q�7���[@��\V�����  
��ݜ�0�2�0Jd�`�����zm��S��[�I'3�fi칀s{0�X��V2�<ʸ�h�S�X�-'S��9
�Kf�9 �N����� J�c��wn%z�k`��%dkw3ʱ"��ݏ �i���Z�i-��cv��1_.W��r�7=�H������%��ă�� ��tZ[�W@���YM�3{I�ЯC���MNח:�]e��@�@8B�^b^��1�z��޵s�,}�y^|�PVmd�Wf�m6=f����@5l~ea\�� �PEИ��*8�9r9J��D��Қ[����9�+:����(R��+�SS�<ƀ���6��y�8f�IL!�6`��[���[q�1����Bd��Xc�`.��Dz��8{�`�q����"ε�88G�#|�5�"��6���;�#���TL!ý0�@P
����P��hF��L�Md�k���0�˺7rP�)�W�
����,b��8@ 8QYR���g|�b�ଝlt��i%r����X��o�=��_,���#�	����PDmWV����}���>od�;���?�������/�]���Nvn�RzÞ��,;&.F�c����,��j�]7˅�� ���*�>F����=�ڙ�L���C7����/��E;t��5g(WC䒯�
�uobO�`�JF6�w�:U�)��P���Vzx�fk����J�b_*D�bY�Z� ���:��.�l��*�l�����md��LVSpu�?�N�N��K�� ��^�����$f��C���+�^�T�}O���<��Vd:Ӡ���<L�Z�\7��]�'��"I�7�����ܪ\����:�?��Xy�"��G�DY{A
��tG0T[�sǑ)�G�X��d}��g�>{)�o1	�R��ز���P�n���*6n��A-6G�"}�c��t��#;(٣/ �8��p1S'Qɚ�F�48T�[� ؠFT"�$#��cv�g�r6f�p|]79��>��L_O� E�F��� Jm����d�6�f2�@��r��v� �b���JZ�R�ZاYb�HI�.ձ��ǿ�!�E�a?����l��J����*ԝ�%Џ�ǝj�6๤'�EG5@;O8L�J����+Ip����Q�&>h1\�>��`���oٹe��g:��TI��j���L����1���L� ��pB�����׼Ep��6�风:��7PY`�����VF�񃱖5��	�MG�4�Z�e�&�{��`��WE�X��@Ѫ���^�1��j�-Afk�V=C��q�B�c3��,GYl�- '�qĺ5'��"<E��՜��������̒�%�.���ʙ>�l|�ד������B�q��D��Js�/b�RvS:�P���چ�;F�	���L=�$>���0���W-�ƃ9��:qӂ��[A�`\�����:�YZ���q��1`M�&�`i*�C��Q�^6�t�1"- Z%2:;����Q���%�>��1X���V�$����Ѽ&���c,  �(+i�P�֧j4����\��8�Dʍ�4#��Qr4ˀ"FZ9_K�����+�����nEn۫Qc����2�,dF��Nz��������=�>��6��'��P����'������|�]?A�����F~>Dj�����#�PoȬuVL�o�v�(�/1�ȲG�P��88��z�f���}Pg"���Q�
9�N��~��Z��j�F}}`�����b���(\3�N��W�2��>�L�c��Xc'd���A�|6Z"+ 9��c5R�+����m��ո�S���9X�dN�y�궀���s����9Ijb�f������.?)�z\�+{�|c�`&�t�<c><��9N(��	�Mb0�=eL"p��@`hp�x�pfi\�����&#�1�GL��ʚ�$�n���Z���9�01�S��Q��ңSN�J�^ۗm��B�*2n�VH}���닃i,2v���`��i�K�%�^��Y �f���|D�a�z~;�k=��ǱJ�v��AyX"P��ߛa���(����F���G���A�:��#i��U��*n�х
ϧ#n s!U��]!�Fy˩��pt��t���DF����{�1d(�M�e�^�o��a��V}�Ì�eX+y�;J����N�T��j�w?�~4Ǟ➰�#�"ҥ{\�x�##�a0X�h�}Ig�wP����hQ�JX"��q:bf�Hol��fM"��WP��;�=����X*Ps�L�������+�_�����2�0�9�bǲ���c�!��E�3T��睗�l�����8�¹_o�n���d�3B��'o�z͞F�~���@Z�p�N� �uT!������n��N�I� T�NiҜ�"�5�l f"�{��HP�,�##�AvP{2��+k��Y�(�w�FH�Jx&(,]�	� ��Qß��c;l{5�f3�|DZA��Mt�cy��O�}%�10���!�rX�$�������f�Z�C4K����{eϸ� A��)4�5��/�&�&��ڪic��=:���пD?{��t���Y-]!F�`��T�N㎌�y���+��������d���=W�5O���f���k녧 ��ׯ��lf�͑���߰�j���_��P����ɐuL8���'�����@z�f��E�G��l`�n6���A۹������&ө�ypn��X�J�����Q���"{�3P�1CZ�ԫ��X���o��I*�חl-��fG�hv�\�A�:��Jq��G�ѽ^N�v���5��UP�Db#z"˚�K�^��Y*�E���t��dD�q��7?���]]�=bd���@:h�Pj��r�M�����y���	Y+#�9��Y.MB4�k�Β��@�֐�ě�Q�?�Jv�2��g3[ȏz��o>2P��R�<���w��,ãJ
M�r�a�z	V��x�_�5�������>Ϟ��5��W�7�n�ƆW���N�ͽn�E�&�(qvn%�W���x��x�).��������C��_Q�,��[9(40�-@v� ��^�"_o��K�P<{�R._�����䃾F̹���!A����{���t!��:�f�{���$d���6t2J��	u��9�w4��	�Ų�(���oD�e��)I��#'�A)͙��^���6�t(�Òi�%�"w �9z7�BG��,�X�Q_���2���;�0���i'.�cBVJ�)7_C��l\aD*�H�ID�����_�3�:�i���|y8�II)rm0����^�|�����e}5b���J5�����p8C�_�kz���2Ӭa�!�>�-��i^�q�h��&|� ��2�i[<qcm
�\\��yT���k�H2W�ڷ0�r��́��Y��8�����U-��d����-sI��AԩNwp�T_#�\�β���1�_���ɥ�y��!����k�a:TΊ�_>-Y�x�2?�Eq�]0��,*o�d<����9��=(u���q0E�;�{!<[-5�L�� F�W +9�b@?J$=��-�\�5Ph��|~v"C�=�/����V�D���E�Xf�g����?h���~fDS<��k��F��o�B ��@�^Z��!I1<���p$��'蟯.���ŕ�?��
�Ѻ�/ $�+B?{d����������k���a*�q�<h��k����]G鞁	���}�=d'z\W�#ia�3���݋ж������������8�����,B�JNM�'�xh�t��w� ������������_Qu��k�>��0t�� � ���5^DȘ	m��ľ9�[���C��V.��J�o���_���v�2t�̩�Ƴ��3���&�#D�14m�>f_���Z�/�9�����ԇ|�8&���E..�Z��\���=1��Ԗ����Qu������Hɳ��^>������ܢ �ݤ]s�I�{�ȄtS�Z�}d{ܕF��F����SY�e)%B��O:���І�����X|ٓ�%���8Ud�V�M:�X��,26��
%�ꓸ;�͜d�'��s����>�?���^�s����>��h(}:E�s �9�q#}�j��y�χ�u	f�c��N�Ԛ�jKÞg}�&ѿ�p~�5������&٤/�L�18C{v=�1�0Q��Ud%\���rH(�R�o����x {�@զ��B@V[5�+j�;g\�_�%8s���b!>�?-�������� k5�����z�6p~�<�����]�Hf�O�D�u\�'���37
W�r�bds���֣DY�N|�.���܎��02`2K I�MG�cg@���
u�T�={�3�Ʒ�Z���d���3�	d�=b�2��{�E��
@d�����4X���,�3aM���
���i�u/#��v�q���0�{{Pd���u.��kذ.+��4��&
÷��pG�#@�o��(�?H_?�r��( ��H� ~��u�w��5�eu�)*�a]q�<�M(7[�&d��m>�(��g�;Оܓ�n��
0���}�QG�����
C0pf,��L?��9H�ALA5È�r�4q��8S{����J�w��!�q�F��z"⠺W��{=ή�k%
��>V�����^_�C/]�����:��_yb�����k{��\k�6�Pưg�_�����AA�ד�Fs(�?Ne�^���Q�
#�W?2 ���p��|u�+��_�D.���eGD�k�<�X��[�OD�'�(�R������`��j�w�Xp���~f�j�M=��ܺR�k���d�:�B2u����Ǐ���p�Yчl���[���Ӱ; ��1��cR��ű��/�\N�r��'�ɳ��G޾�s}�P�oB[ ����C{ŗ�GfnB�\ج���1���B����[��Q=���<�{��B�����x(ы�d����{�甑E�PQ��������Tԑ'G:4����V��_�����0�VV��k�y-[50���K]g����:�QN��]����w#��"��G~�$5�[�]���9��B�],
H��s�\+H�$�a�z�$�/I����;yn���N���p�Ȏ+�ie>x�k�����������"[��>�=k������v���rsilY�X��2����'��-K�Ya�`e�u�̮�������Zx�F3<�1K�M�ׁ3�6+Tl�`(2�P|(2��j��<��V�
Bh/��mc�Xڗ�&7����D�ӟ={&�R���`$��Pv�U�G�v��0��m���d.��d��3���|ns�j�G���0�_��=�L�l L����h0��XW,SoBUH<Kf�Y'��
�툛���S׾JĿ�]��lo���W�Փ�8>P����~���2��ݐyi8���2���3��O�!��-��i�J��A��bϗ=��ϊ&�&����ǔ����Њ�"������ҹ�S�:~cw߀$�P�A5;]CXCعf�o��Z^��'��hz�c��a�K8��W�2��xo?���w蠟Q�HD��nQ{P�I�Vy���-n�nG�/ա�TƯ_�D���F��f�S}���d���E�A���QbjUqBzԕf�˽)zE���x����ܮΆ���"ݾ�[u��G��]��H��o�8{������Z܁�]8ƅ��qcN���JL`\� p�ɘJe :��3��/l�W@Q����\x�WU�w8?h������sd(���٢>��a"?|����"�_-�x@q8h �>��j�^�O��H�l,S?�cH�ߡ��������c|����~�ܥm�ڗ�C�N3ڰ2�~G�����7���^�l!��� z��_]���Y�����߿e�d<�*�fi�DÒ>9�=���,�sX�P�:��'ǭPU�K�Sr�hYpGC:��"=�i�w+qlI�2�w��#�C�j<�}�MC�j�:Na>ې��� �i�S��쫕C�-d�y�����K���Ծ��x���ޠ
����S<�*<;�hrk�����;|G�(�Boߪ/�s7P�#��}�ٳ,l���5񔯼7q�*G��u� ��V�6z����>'�� ��T�B�4rG���;�E��m�S�׫{`����7�����兔?���bO���YE)*?��>l|�dc�G2��O2u�B<��%62������}M�4p�h�p�i`��WkV��|8R���A�HqA�"/�_y��J~����|����;M���*�M��z�����_�A�%b���G�dS&��[��8p���W�{���}�?w�Q\`�j�C	s����G��ei�Wz�������^pv������=�w�N��?�9��۳�Tj�:��a���,�Ƀ� �l(gbl���Dd�\r$�:hV���N7�Bw@�b͑��jx��;��Q㸅p�f$��J3�5{�$�#���
��J�E��J7w�n��Ȝ�c$K���ȶ^�X�w�N5���^nN�S˥i�8��.5h(���7 ���Tyj%��0Ɨ���yZ�:��������'�zcc�)^B�)&9ʱ"����� ��z~�:HdS۾�tr'�F@I�7S�N@�3�E%�t���'
�\6��?���������c�@3���AvS�L��y��8�7�r���>�DmA���f��>Anu����ۓ2S'�a<�K+�jp��ҽ���#ˢ���S�Z ^��-VNX�l�G<Gb �ϱ��W���	�`��c�2'gp"(�r�_���+��g�+н�ԟ-�D���m�+�:/��?�0�8���B�>!3�d���rB&kA [~F�=錣_�� �<��DG��a8�}aA��N�A�Wt�A� �	��D�������B�����x}P�a����|�'*{�|h�(y��w{�$q@u��O(d�qR��o�����wr���p�j������6%ɏj����.�j�6�_����s�@���\�V����M��I�c���f-+��9D� ��R�
BN��p��1��BW,��B�g�k'�+�U�e@��'�%ڗ"��8��
��S��;
��ګ�����g2��$��@%c�?�ՠ�_u�>��a��i����q��s���cl�N0W�'�	�R<gyjӸ���g�Oz}��Ew��Du��m���������=IG3[�e�ۍ�@1���ܾ��c86�}����6[���Im$��I4J^0��Ϟ�tS�|�H3�H4 D�M>�������7`lS��Qz��hx���Y&#dB ��>0J��1F����Ɔ���)�ڊ��U�a	�ml\��[�1{�0u�gaq�81�ِ7�����Pl��v�E~������}�:EQ�%g~t<6b�ڷ�����Yp����G#_P�folS��t�)���^�'5�=�i��j�&n��������k��5�,Ӫ��w�@Ї[��=P��P���`�X���ni�A��AH�$Ʋ1�����\��B���fG	�`\�� ��|Y�`�
$ƈm��E��AeH[OE I͓�|��n��,�'�ekq)�7�;�9Ƣ�[�ư��ap~F���X��h���upO���D�o0��x�D9D�Gt�)���,�z`�����ǵ�����y�6�c���⍑��]�9!�xq� ��Վ����ω�z�6�*��0~���1D��C�A~<�Ad�x�(�5;+�C`�nZg���S\cD1B^�7���(�̧T��7�l�dVC=��6΍�rX������\�k,��F+2~�����k���F��T�nN�w�Aۈl
'ԡo5�Y��t�Q�����>�yp"����O��]�J�?�]���)6���� �LPgb� z��߽�����aB���tگ=�ePs����[}S�V��d���_m8�0��y3���N�=�؞l��E�'���m�^��ח��kt�C�K �XY��2�°��H(���<�K���Y���h�}6꫱�5+WÄ�f�˃E�(���3�t%a4d�lI��U(U01���S1�Mu��}��YK	1��7P�C�If�H������G��2<��Ló�H.�� N�!�!��V�N��+�&%���Ȳ��J7�H���-I�C�s����@,pxOԙ��=@����Y�E�H}( t��:Z<���eH�?�)��ד�*V>��BI��\��� j��1��ifxyM����?�d�&-c�����\��v�R��ymVl=@lgqx��Ɏ���P��1��r嶤�ԢI�������ک�@p���r&_J�2dTz~Yc*Wx�V�����b���F�x/5�I#�,\Ae1����T�Ԁ�ʃ��kSp#�ȉC�C��?���u�_��Y �f��	ӞG1�C����:�!�ԗ��6s�և,����
i���d���~�j|�!�ht����y*a��@`,
2DwQ���)��=ÛȨJ��@ ��i{��8�E�Pz�aL!����P-�l�S�s?�@�ƪ�ld{���������86�#y]T`b�4���A� n�2ƚ�7P`c��5 �	 ;��8]���R�?e��}q./��<;���^����D�DP2K�z��6��O�]ڤG�#=&8�/޼���|��Ǟ��p��AW��	���C[@��f!h��j�EV`��|�d���R��N�܂U9��vc�b��@�a1�J�
���^b� �M|R8�>Ӎ�TE��yym���<Z!���6�9�mQ�sB�Y��-.^�VG$$2�r�+{���__�Cw�4nx3���-J�g�#$�B�%\a�U����}��z�q��6R��Ǚ�����=d� �G]�?�dno�^��aFr���<{񜟿Ԡ���~�n6� �Z�F'AFmjm�х����<�a亠��L��[��?�su>ٮ�(Mg�e&@�
LY���xT��id��w�dpv.}m�qJ�[�Xd_��ٯ�W��| � z�S�'Pk�?���{�Ɔ�{�Ě��5p�c�����0�����{��LM�}����t�ʱZ�Q g��aO���t.H������3]\ʳ�H�[�6�Y.e������1@�eÆ�]�'豜sc2 �P��A�
B��(��3�;A�4Ե7����f��j.���sG� +S����~%o�ƲҬo���5$u5[��+[�������q��d&�r[j�cF�4C��gN�F����K��O=�����Y��F� ;�����l�H�)*;^�@ƴU��h���F�կ�w�������D�q;ge��
�}�g�y%ݟ�:@֫���Ĩl4%T�P��k3�ɱ:L|T�{:L�(L�#Z�$3c¿m6�
q^���s>��q�>���[m4�r���z���k��ΐ�e��*�y-��8�k"KD����5X��:��A�`������)]o1�pa+=i���,d�O�n�{� T��C� =��])����t�=<N���ھ�ԕ��J��B6��+=�?���[�����=W���O���b ���O���HNX�;XK��:��U��~K�%ޏ�R��6ńtn����d��	�r �)�8ں�@��ī����L��G-��V�Y�|,� �8��	�!����OU��g��^@��D�K��A��З���HXd��id� 4��PF��D�~.���2W]}]D�bKf��n�T�tS�ԁ���(0��C��5㱜_?c	n�yw��������B�`5��<�{��30XⲮf�J��\�tQvw��u�v ������=�%4C�Q���Đ֏z~`$s��Pbè���d��*��w�RCvU��pY���d���,t8�1�z�X�"1>��@�J���}��O˧D'��F�'e��9u��0F[5r ϰ��5�$�1@�d�F'Wǚ�Aːil׌�I�6F]��c��b�Z	�S^
u݅[K5$P�K�g�)����5ru��S"˩��#���gI�Me�����R��KY��@����[��2�lVU�j1��A���;�4��5�4�Xu��A9�<a�9�{�<�۹c&�W�N�Ó���q��s\�? >�#��<� ���7Nc�A
�0nI�3��u�'@֧_�<9�X��W���3�mv��Wn�ɓ���hbs��3���V�	��η�t^U�U#��p���}Y��K��j8p�G�;s�F�H!+�����{B��?�)�$��f�C5(b��q���(�1��u����tMu�ƂN���:�ݝ8r�o�^�k�j|� :Q.+u�@�Cԩ(�	W2W[pxx�����W�w�L���S���o�sb|0)usf�`\D�@��0ujOμ��U�m̳���k5g��G�&z�hv�Hǆ=�B�O�?�ԯQ��p|��t������=�g��'����8��{�gh9��F<��rm��� ��%�ubo�4 K�����е[��V/��F��n��/}��^�}Ťk��8�m��kQ@�z4�E��H�D�������a�/�CGv��nP�ܫ3XϤ��ɍΘ��q`�\�Y�Q(�\]���Pz�XL)K52��J7M�2j`\�+]�~E6n�~WG���,�׫�[��b-g�ݨ�s@�\�'R2Yf��q�{�Sq����#7�%J��K�tm��uc/�z\J������e֥S j7�L��DH�9�Ԩ�=��Q̲��X�Դ��&�6}>4�S=�?W�oNJ��;��&y��,�H�^~>�l`�ʠ{~��q=[2�g�W�w�ר���m��I���FP�!�sE�5�pa��I9���a�hp8��,��5x@6
`�(Q��p/i�"�;�Q�ѵ���R#�������?�(����x�``9V��9�빌5��`��k��wFW��+S$|��C)����'��s��t?�ύ�����S���`�X[b�-5�<"��z�0�d@��/T�nC�.2�Il�%L3��0��Z�T�I�؋���(��`�T]����p�:ed͍��=�4�?���b���/GY�f�#Ϋ�>Ig=s��a�j�t##��vg�qG%�m���� �+�-P�m�^�~f�*�B��B�;�@�`���*T���'%�Vg�TD�� B���p�QB_�S�hж[k ��h*i>e�s��[��,+�C�4��	{�{M�����גB��f�,�2u�r6�[Ƕ���+�_�'���s/թΧV�jg/�#*�mVH��jș��u���si��o߾�;@�`⣨���R������>;�@}�ɘ:�gW�L��ۍ�ݏ��GY>��pL0D����o��m��{l�fb#�X(/�f���B�z�P��X�����ʭe�>�R��cZ���hp]  �M,�V��!Tu�Z�i&���M:U2؅:_�i�#�R�f�����澗�ѵs���}��t5;���l!g0��h�IX��x����j ��3��SYL��1�t;��7�1W�(�`�z-�Ӆ{���sr(C3.gv+b�`�3��;T����@`�~&��1)���D��!�{Z*���p��f�Ա���~5�e�hs�u�U��7�2e�-4��*x�;����T�@8q5J����g.�@�>�d*�@��7�- 3 \�i�~q1VG>��c�6_�=�������+�;5�����n�^ʃ>�9Dy�(�S�X�	�d�9BI���s���z�0��Z��ʘ������V��5z���J����i���߱GH�;C�s��k@��~#�ਏS�m��ƐǾ�ǲ��hDR�ϒ��x�9�qmU���%��Tk߻.=۞]R䝦W��#�	/X�(ra�Ͼ\����G@��#"gϷ$0��
���������Q�@<H��L���IÜp�#>j*P��>���B � �$ә�8И_��Gb��k����zK�{����Q�oN�Ӑ��
~���؍�`�{� 'xX��f��-�(���$����
�`O�kn��u�\~�Q��"*�� �^[�6����+ZQǂB �X�]W�/_ȫ����o/�Ŗ���gW2|v)��,4���~!�r#ww���}[��]6�I�בR�X4���_��U��-�����ׯ��{j�3β�<`�yv/@�5͡�Sd�l��r��_���ʃb*j47,�`C�6{Yk$�HwGƳ2j�c�d"�]�Cۡ��߳g��o�û�\��#}� ��4�������Q�������28u*�ɂ�7W#?DO�?f�����L��5�D����C�F�3�%���纫_�r��&�~��Ѯ�"=W@�2��K��ݰ��^����+��*ʀ�zuS��$�oO���~�b��V�|)�m%(%i�z�������\���F�"	CY[	�r�@�/�y�~.���bil|�Bu���+"�&jw����� !M���r�x#l���qB A �b�:�^8O'3*��]�3I5h�K��1b$,��%��.�9�˂���l��f���l��jKz'����^�8���PVOfҨaD)e_������ݍl՘��w$��O5���L����\�Nz������\Y��k6q��!g�W R��?r�F[��m�?5�Noe��{�f���n{�6��8��x�A�࿫8(��J��3����lz<&K���[+��&'^ �U�� h3�\��p�nł�Dl�-T&���}�k
����(SM}�f�v�b��$�| ���hӭ_�#d喉�1n<�L�%�/ #Ʊ6��W�l�0LG�y�G��!����HZ�t��={M.���{bA
*m�>F���L��#b���k�� I��]�8�X�m�!�M�\�ZEk��@nS�{n7k��ݱ%��0�E�����n�*�s��he�����ޡ4�M����_���d��(>|`�~E�H�m����������L��_�Uf��{�z~-W�^��3yT��i�l��si�=7�.��%�`�S�CAGFBM�
F_��ꝟ�'��@�w����J	�e60�� 	�������/
�7F����8Ӭh/�݂Q6&7��nt�?| �[�6��g����#�BJ�_K�1 2�ёqZ�VҠ`и+��+���|f��S��=??���u�s1�j0�1:�M��4�"�&_%�p�W��y�A��u�K���?�~�*�lb�+�paC��܃��t�����5�F�����!��w# ��0�u�^������{���c�Q�,_�o�V�鍞}�Ih�#2e�L{�C��@n�>Q�j	��|��B&�ѢE�]�D8���ޛ-9�%ס~F�@�9�ح�Q�݇�v_�Lq���"�4RF5�]]U���1c�t}-� "��l=�)�FYVdD��}��q�Z̲�yC��"����`YR���g��8z���^>�s��5�E�4���v�4B�,�]
�9�]j�2׏�N�h�uD.���*����D��3)�j�r���9�to��~����I��:���Hh��0(��5F9׿S��h���2��aq.vg�I ���ue�"�hbd@(�Z��g��)�-d�����	eÐ5��� 3M|����{�>#�x�:9D��2�i�L����):�+��8�o��*��A؂b� w�x��x}�U,�b4Nm#܏�| ���:�;��x.F2z"}ll�3l�DV�����bD� oգ�;ĝ�B<��� ���uҸڮ��~�s�AP%��Jm�8 /"aSY��&Dԃ'�f�N� ���}s�+�.����ggF�]��Dz�!���9W�	���,~k ڂ
��o�u�����&{pr��4@�-�گ���m���)��F�c�p�$n���Z1��:+��߮	4V�~�$ր�����bvj� �� ��r�l^n�d	je@��������`�dv{-��Bb̶S��읁Zʑ���P_�4⮫
�9!�_�X��w(o�M���������5�>W��-�G��sQ��$�۱ޗ:Ud��x4�,o4�[�(F�q�ژ��� tRL��%4g� j�CB
�_�[CIW��O���g�mW7�|"óK�n`X���LD���Jh�Q�k8���i��Kz+7��&=�0ބ��'����nv[�:af�˶��v�d����I�j�w"MeN��������p\s��n�h�"�
2�Wtš�	C+8��q��V�G����xy�GO����"����c+�"7D�]F^���'��}�[Y�uB�z����-X�^�y#'��ނ4B����i8�zOZ,_�˪����|ƾ[gpJp���b%�V����,E�IT>0�{�Y���N�NKu���o�4H4��&�S���_������~�3=o�J�[���D&�-��G�HvR��RR�92����=���9�\�����nN�����͋[�0�\���p�����㠙g�<��]�@R�Tx�-�;��+��g@���O��Y{, ׭�}@�#ˆs��Y����6|q�<౟N�鵳����FQ�����?�|T�qe�0���wT�P�ºB[�?�	��q.N%׽�P�-H�� ��2�t�5EP��Ŏ@W<0�J�@�3& �U���:��]��WWzV��A�t�d�~|==X<v�	�DT�UM��U�eP�����{�į�;�H�li*q�,�{������Ē {�N����������]����u�����掕$��b�r?�a68a�S�k6�b����>�l��8��H��ډ�AP�H��e@8>�ra�Q��݃f�cF����91�~�ͯx�P�_��BQ�.��7��"�Qz�d{�dP���rNCC5*2���1���=f�5�*{���wWrzq.���wr����Vsyx���ȄO:�t�P��9�����  ��IDAT'�:-�.�c��c���9�}K��V�Ǿ�|	�Ȓcxp��gN��z����3W��`����ޘ��M�=��lE��%S]�:����F{�P2u��=�f���ci��hPԘ ��W*'Xil�'	�"r0�!D�3�� {���:����J�l!˼���^�����V�Q���j2��]*��kub[���ou���0������ک|��F�o��e�L���|���/�>�D#�_����B}�:��s˩Fz%F�`d5��Z?AWx]5,�e�n��-�J�U%����5�L���׋����uQib2U=*Y��z�8v.�g*���>%Ħ�#/���3�e��Xϛh2�a�<��,�'��!��}V2t8�����1��E��k��ǔ�9)U�����{�N2(�vk��R�)`��㏁i����>����g�~o&`���_��}��̘�J� �8��y�h�/�;ݓww2S{������#V��h5��ۡg���>Le���D�i%]��g��L��G/���s������S��}�Z���t�iT��v(�G����;Ͽ�>�+E�w�\��b����H��a0|��B�v9������\>���խDU�IK_��2�l4Q�SHi6Y�-0�j��=19�'j7��<���g��cJ#f�"OI2��F�q$���J����	�X.�#����힇�x�D*��wz|�K��ة�Wf�zh�ݵ#C�"��]�*Q]����-af���Eo ��s)��r���c�k'���;��IS��Z�F�]d���9����Y��jI4)f��h�P�{R��7�y{�����ͷ_�T�����ꚑ�bZ�=�'�N8�W'�*M)B��`�pXD�m�����r���`�pȣ4rA3�|v�	�~B��1G�r�f���U$�H�
��*��J���\Y.�m]!�I���g�rd����a��ʍ�-��s�/3�ƌ;����a����X�o��ʘi�> ��~7�F�6��6��7��iv��v.�j �ɽ��WT`�M%� �G���+p����R�x&K �T�i6��ý��� �}�]/�8���8�Y� �3����u1O������~�%��bN�)kHsf|�t6,n��:𮣯������7 nC����k������Hi*c<k�����]{#������{��>u�7TCF��|?=�w�O��^�չ�ukp��5F��$�������}�5�����?�����qvn��OC����p�K���`5�=>8"P"�|�d.��,t�AL����:��/�4�\�t�@t���6�{JHO~� �	�/����1��w�v'��{h%b�sT��C�)v�-��2,���}R���l�tɁo �1l��j��^���%���U�8�/t��|���}�Y[:���}��f�������Y�+��Ǥ�E�Ӎ#�*u4�^k�VIT`W�Z�bDF$�!em��6տ����E;t��Y��|r8 ��@�Aؔ�v�Պ�m`�z}Y��E	 2�s���~�����H�b�?u�Z�҂���1[;�F1�D� 20�ci'�h�?����I�x����"k��7�~'�:���@5�h��`�tv.$C��肞X�6�	@���}���#�0�}f\��T7�P���%�*c���2�
�=pi��l:��

�D���ȑ����ѾT�H?Y�����=��m� ���:r8H��A����8�����%�8ҝ��� |�`j��m0jf�m��1�����r����LW�Sg>�}4��h:����53�}�J��=��{�4��?]}�߽{/�ٌ�N��g��c5���9��!+C=}�n��A�/ʥ%���4�|����R��C	{���(]�&���(h��Q�)EE�#�MW�k��O=������D��N��v��W��P	�5D�qC���I[���{=�G��m�.5���'ZB_�s����@���5��zT�hu:f�<3���'OH��j�z�co]�HP�6yt��Y1ҙ��c��@�/�"�w鯯@�@,"F�b̭�}fj C�jd�x�P��� &�8p��VH�N~��{�����)k��pI��P����Ag���
hm�QM�6�V�Tx�DAD3���8�AemF �<���S���@�??�L:�����f�$nK>���Xħk���g�sŘ�Vm���AJ}�o�cF��.���Ann�H�j�ח�%;��� ׅA�b���4-�k��n��,�E;t�����0cjQ�Z�4�^����VF�]���%EŹ��2+���FQ�|�� P���D]a}N��sR�q
����ƈ0j�{K�h�ǋ��
��ܭ�O���9����k�P�jl�u�I`�G&�ϐxِV??��`��j_ݠ�.U戨5K��=�ԣa�~�v����ຖ��}0���� zE�6���X�6�G��v��0AfI�>5��?9 �bg�2�8����z?�zp����D�F��%�c�����'��i|jJ�xAJZR�v�cfj�:�1'���,�u����D~�����o��~&��n6�3�ek �����>x֗�W�{�L�!�����y?�ɵI���� ��5ԬN��L�z���dA�!J,�7�d*���z%�NW��Vno��4-�D�!V�c�5B�a��x��up=�O�t�����?�U�"9̣C���N���pJɏJεV�������pn�nk�)�Lػ��k���>��f��=M�G�{�qg�4��������k=r�������_���#����&EX���a|_ ��_��`�ά�N}S��/��bx�ޗ�a�R�W�T�MqC@��R�[up�[u�& �/���+ �&��p��.&r����k�x�E?�0\�ۤf߆P�؇#oI�k�`�(����5�.��?}�=�R �"`)7P�,hвĨ_��}J��L&8����<�N�4�����~*�{�F=��R�zń��&F���ڜ�s��{�o���{<�h����)��Jb���̉����0�F��P#\��r���@'W֓�����f��^��o4���xRr		A���0rXl�eD��c�9]*����X7&�����f��lf+y��;����G���2�χ��,*U�".;�.2+E�3a�L�c�l+�h����j�Xa�I�R��k.jG?o���1��*�Z��tOO�;ԬR�ۡ~����/�*�D�O��$�Ou�o� �����̡��C�N؀rv�a0@�:׵�׀l�׼%B<���'���4��d�
�Y�C�-���O�b6��%��ə~�vK�.Ne0�x�xW3��/d�k��J���������շ�I���l�OhK�ablY.�� ��tz�W�Zn*�V�� ���j�&��9�4oK��tY4r].��|)?^_�V��g��j}��5kv8���j�E/m�Q�Ħ�ſЪ��>�e����K��5>uΕ�z��x���]S�����t/?Z;KPY�ϕ��:�qb\6�uh��Q�ՠ���3�-P��}��'(�^��<�����#��gK�ʙ���9|��Q�j�y���l��B�y� I�-��A���ص����ŋ�r����o~�Y�>|��jt/a�����f��Ӂ|�W�J+�����+�:�50%�� �y� �p�/�B��K �qm�4���$�%�:۝VH�E3�1hkG�?;�DF�aO�q�E�^��[�����Rm�G=+��'2E���c>0����&���ܰMЭ7Uq�������&Zm�=����o�x��̐ݶ�V2P8��*�=�s��l�������!
�4;���"�e=��#u j�C�l�F�}5�g'�-�m>������Pƚ��kX[�YC�Y�Q���T|�k+�i��R���p,j�)�]�5-�'CP�d*��w��cN��ћR[�/���Q* $�:���j�N}�����������F��m�H�qZ�*��5nqL�R
8K��$����1�oK�F��I�%wM_�NC4�7�Q�O��T�sr�w
�H#�J���	T���F4���256͠i����zvN"���`�e�P�����W8��g�c�������c�H>�o6�W3��,��U�R��ɬ�����˭��:����?�X���tC&t��]m�ǉf@�G����f9E'H�b }&ӑ:愽�{�����2��oW;IgKR�~��7_I�Ӗsp�#(�L�W����ZZY�G�џ��#��Q&��@�3�5G%l,+�2�9��qd�2����=9�e���G��G��0����~x��Ge���m&��������*���C	ߞ`�;8U�;�_���Y�ѷǠ�����V�G���CdH��n��@���j`� =�`�CfKe��Jp�vf��s�Պ��#�Ƙ�����o����d�^�L��D9��ȑ2��F��jƫ�(@���rKpf�w��I9-�|�Ϋ���.��_;�Dm3���I������` ��Q�e
"'0;�� �݆D>��k������z���o� ����&?���-��~��n��ST�Ff(,����� �ŕ&C��[�B��|q��/ڡIX�Ω��Y9/%�Q�.�cـTd�1�
��jmB����j(S ���#��#�"@����7����x�+kU>?���t�R�&��Fm�p3�4�E��;}��{0�D��W�l��V��| �V@��弞O��A\wd��K�6x�/����mK�{��b(z��@���&�ې�:���,�H�̝AGzg�4�xw�^;ХW��]���D_����t~@�ԇ� J�=�@wp��/����Nf*�O`� �׈�l��]*�r�jYj���L+Ø����y� "�p?�|�9� 0٦Vt��v�\�p����[[�Ԟ%U�tf���Q�r7$LWj��#2�]K��Q°'wz-л�p�5 ��{%zO��is��=_l��n#m��~G:�b�?\�(�c_w(ﯯe	�� 9 ����
��<OO�e<<��.���n$�������:��|�6N�y~?�g�v�*�Wfݑ�^'��u|��bT�!W�&�&)p:�L0vG#hOyx�wt���Rz@��~p��G�w���� ��{�E3�h����Q���f��U����=����-h��Г�*�1�����~'�9R�?k�X���wbqU��>r�$%��$��ϭ�����B9���4�+�b*�场�-�s�a���7GGƏ��2S�k��s�&�P�T	��# c��(SJA���B+�����LFL�@�g��iꄡ����9����u=l�?OR�R��e)in��1z
@�I����C�%Z�E)[���ke���~@�L�cH^;8�>r�_&����Q�G����j�%)��'������R<���#�����$���"-}��]}�/�N"&;��A��V�T�1�2JR���#R:��)+�"o�5�֋����T�5�<���˗�_���+w�i��nN�9�I�L�-F�� ��j!#N�Td."�}#m)˛ � ���]
]h��Y��d9]HK3U�쿭�ux2�����W/�Q����ʽf��w�������.����6����K�YmW����Rd�'���$t�4���c�]�Aǃ��/5�;�n��oIQ�ĵ�ȵ��r�"Tق�����#:(H�2(��w�#�..���0���F/.����f��B���ܱK�QC~����(a�կ��o��f)?_����y���L&��:vڧj,��7`ہ�YC�Й�:�ӊ�!3�GC�z�Cƭ��d��~�~?FF��J~^�I�1TC���R �5�j��D(v��2���w��q�|z�����0gh�ʦ:�D�gN���{���q�80<Vգ�AE�WU�#��h�����c?_��e=ή�{���s�#$}�y��������;\s�E�Ǩ}V9>�n ����#��U�% ���ƒ�*�����ivt���[�u���.$!9�z����,~���5pĨ���R�T^�h��pn?�����Zv�;������������b��%�%l(D�p��$4	�kn���,�թ>hsus-�~�j�������m0�i𚓊ّ<����[�?������Lk��A�͙}�ظ0*
�(TI�t�">z�$�o��F��o~|�],K?�P�� �3Mj)��*ؕ42��u��&_�����D�bN��N��Q�f(=��-JD�[�#7t�'��<%u�G����n��Y>"�a�U߱���Mm��x`C$��Ě�}���ԡ�=Ld3y�rz��^q��y��v��55�n�����(vU�T�!�:j1s.���]���N��� ������v[ryv";�΢0i
�I�-k=���D��������b�ia���г� �H�jl�$;�ܼ���˦I������)5:Y�G� �;3j8p@�����IK�]��=������+5HZ��J�2`�+6��tQR�$���w����F{������r�r�k{�"��E���Ʊ:Ӭ�{mܰ̍�y�)̐ӏ���{I�VO����9}d
z�f�
�J�r�h0��S Է]@�jA�}�Z0m�7��5H�b��E�Z� p��ˢ�=t��f�h<������2��`�����F�,��i.��1p���A;����@	Zy�g�Z�y�q���}��P��,X��e�j�����w=e��	V��A���}���`�v8��̅F?{`��6%��/d�\Y��e���5���z����l�T���-��	N(c ���Z3Е��p�����q���A� ��M�v�^�*I-�$;�ELeH��7�7��qc�Y1*}�(�d�Dk&U[�#�b ̇�t�:u��@�
�u�5�q��*ri�3� f�� �-+I�Z���TG���פ42�Q�Ĝ27��d�ɀkƨj�B"`µC�����ꋱ<���2�-�i����b���}a�/ۡǇ��?���J
f�C%�r/�T� ɲ��Ι���u�O�L'�0�YD +5뤪[�Mr� ��BĆL�s�KO]=�n�&6���g�b<�)�e��0j�Q���A�6�L�Қ���Ԣ8�힔e�Lf��Z��b�	A��6�������\H?2e88�����@����}}6�)�ɋҘ� r�C:�����Ȁ~�P��<2�V.�@d4���j�S���5��jc4���+�B�(��'��Q"i�}�c�s����#?�x�.��}�ƳBq��}�{v)/]g^�����0�-͈��L��Lr9�^�%��%����`��j����ȵ�Ku�UF�����--���JM���Q���M�k��7뵢��}Iiw�R��F6#q��%���{:������������9���Y�n����TDX���O��>��
�nNuVsL
�׬h�n�k:���0�U߬�lH�ĝ�!���U�����s^�����[����Sg�L�?�j�\[�5���U̒����x��\{˃Ah��F�w�r��;jcB����s�M[�;��H�r
 ��#k$��"�O��O��2�V��s]�u��yFÍ�Y�]�g���dc��pSט�~#��C��.�=It��//���ԕ����i 0���<]=���k9A�|b��Q���.�g.�y0¹o���IL�Pu0�9�k����������v��hLB0G^��Od��lgDl��z�&o}b�8��f�~��
��k��C�se�z�Ҏ#v�f� ����R�evd�GF��s�C�_�a ���B0�VZ��Kv��k'Ihh�ч�A�ҫ�����>ș:*h��43�uz&���?�-9��^-�:G�������*n,d���E
a��#C��Vg�w��8S�ܦ(HI�^Ia��A��o�u�r��:�t��9ˬ@@0�L��~����>w�1Q�_�|.ɺ%�Ȳ �I����_]x�� �3�e/]L#�L�U�&]͆ ��ڒ����S�	���񶩑��H�* q�[�t �0��h	2|�~?�_-�R�qic�XK\��EA��e�?��j*��P����9��DƩ?�@��fj�0*s���/%����a/�u�c����`KC��jU�&nIO�a�e��"X\���[ir���}���?|^�5u�A���|���� @Ρ������9�f�gK�z������>ϏX��Ĭ/F�J�DXZ^3�!��M���%��e�����������Q���>�g�����@!�ң9�����G'��;�_�k����CU�^��Ʌ�;u�K��Hr�R����v-���ϵj9�K<(���Y ��"o�My���QJ�ĸ��?[v�+�
�Yc/��7^r�i���:T��WR�Zk%m��P����N������(��4!�ggRi0͑7Hu樊���37��e>Y�%�ԇ=ka��j�!���T2�&3�?a�v����������ۤ�M�D�w7a/bx��A�d���*��*"�c����U�>��ӌ��_^�����<4ڥx�����lj�jq޿m,�Ȣ��(Q���5#G��W������JRuXy��*5�մí�xVn�.dF���@�i�B�)_��~ꨆC������R>^�Hk0�D�e��[�������;y��joSJ�,�C��}�����ҟ�0��� }�1T������4�޶�vQ�^�Φ1pK�Ӗo^��ϓ��DE�9�(������i�קgr2<U�ޕb���dl�5zȖ��$������6���T@��v�����jQC�d����=;�>�-ԙg�/��� ����^6�B9��=����_���!���=jft��(�o�(Zǁ��s� Ԅ��2��N������y����p'��L�o�3i�����<F&z_����ږ�����Bf�,[5BK]��:���O_���j ߵ{,W6�Gɩ~��*s�iq��??���T�`:���� �2�l�'�c���td�:7�v�s��E(�2%2֚E%���QX�
��>2�VdG�ެȃh �K���_�ӳ������ ��v|������Gp �=��Lhj�r�K�����Z�6$3IO�G��9�럁M�@�qpa�����^G��� ��W�~�(O����W��$0:��:�2 �Yi|xe���66Mj! ���*���9F��V�����4�$U��(��B��?��~\>{!��	�yŪ��h$-���dT9a%���sR��N��Q���~.�^���.�%�{w�ҙ�Lt2��{P�D�	0ᘱi��W�>���9���+]R� ��9
謅����f?�3o�(c�#q�B���&��o�4l��8�?�Q���ѱ!��vXGs�V���J-%�]��Qil���F�l��׍�5�l�����)�ׂ8Inh_��nԹ�4���Ʈ�Yo�vA�x��1j���*gY`�S:8���V��Br�4�oߒ��B3�S��)o6��Z2<5�˻�L�3����#�J�ۅf�;fi�+�*a�����X�3fds��X���v������C������C�O�|/�:����:t�~�+͠[2�C		�(y�a�k�36��ۍ��l��*1u%P�fBÂU[3�L�W�����O���l�x�.D�L��!9~�m���j��f��1ā"W�:�}��������um_.5#/r*SLԪ#��d�	���'���7������,֥�����V� *ti�EF�x����^}�h�����
����[����"�LN�^轎d����@ b��.��\�rq>ԏ�%G��L�f�3p@����;�_��~��s����3s���b�#��-���p�k_p�x�2��4al��~OqO�xO�/v������S=�{�\�i��E�m�}�nۇ�chN�jz{l��ļqK-H
cu������?�8d���b�T~M$6M�2}B�ob2���U{̏���O�s� ���1z��!�G�D��
.�_��^���>�.B��D�&k|L���!{��/1��\�b�V5FP�@
iVMa���Z��jG��8��UW���w[]᠇�U��A!�Rm�Z���9�%��U޷G���˅ڽ��33o�-�܂L�]��w��@U"H���&O���C�,j����ҡox}�b_�C�"��Qi"������"����վ��^O�k���Ʉ6�y]�c;��.5�a	�����@ɐ+�2���ȞZg�����ci%8#�He����9�؂�58ث�T���5;��h�ݺ���ֈv�rI;�r�����p�[h�]o��,MD�3��"�Q	��u�5t���X`�����Q.s���N�5+٥F�ŻJ�].���eV�����g�&���ts���-=�(3ɩ����������6�wb���,��]���zO��Q͡���-��%{u� � �A���,�G�콹��K�qT��F ����S��gi�����O���߿���7[��b�c��U��͌:�`�//���_���}'�Mɵ���(70�UCd������̯�� �T0z���Z���LRuί��5{_ˏ�5�I�A�3f`�0��L���~�6�>/�N�|0�K�8����-�	���� ���`&��'�L���&pt�V��p[pȃ����L֓���Y�8[�Ш�]����T���@�����+���,M�cl0�T�����<�臑�c��n����cǲo��1�Y�g��w'2� ��O��l��C�@6�^[���v���:޻�g���<��Ǒ<��1����7��#N�J����!t��v�U�rd��հr��&�4GJ<��(�\R������R	��`��W��ȮǊ�]5�)*1;=��?�(?o_��X�o�����G��ӳ3eӳ�	���G�@�z��J�M��G��-WcQ�L��9/�P�� L��/�AU�cz��>�9x8t��� ���
�{/a��a�,	��'�g�6�3i�������X��&�Ц2�R7�VO�늨�*��jdQ���C��B,RF��f�u�43��Q�42��6>�� -i4Q�#ӡ�Ju3"ӄ �=6gA��{$ `�:�,4��H5ڛ�\�@ֶ �~D,s���Hvr&W�Q������R�z�s5Lg���#�sm�ۜn4Nd:�%�
F� ��9�2�xt[��N:�[���H�-�z#��k���Q��ښ�C�x�)��Mֽ��;��,�M�H�q��5E֯���"��e��ԍ�������L��a�Z�8�� �$�)k���Z�fr?��� hͦ�c�#�()�obԒ<�0�@�j��cB�H���B�*/��8ˍ!;�A���jx4��Ձv4���a=KY��2���lK�h����N��ΗLU�Ufà�Ɍ�,���'.w�(�FTt��2�"��V��d%��L���s���g���������/�d�?8}�L��=�!��G�At��$���j��P����B�| kp1�R����X������c�Yp���c0vB�����!�t�3�5hE�[dҋ��>��z��?\Lb�N���F�k��r&�A�y��ψ���x��Y������K�#r�̉�&�P���
D3��SN��*�f� ��C&tkJy���f��x����~�ۣ�GE�cJs���^�
�҅%%�L�W��@���`L�ĴMfSzz�C�<��T��F�48f�Qv��Y�h�Mm� P�湞��>�֪YYd��s�\�C�'��"�!��A��x�D�~�,޾�>~�����b����[�ݮ[9��ྂ& ��R�~M;����Qv�~'���D�����Ϣ{	ﵞC�_��f��-���߁d�����^��)|�I�T�mC�&���7���-=w8�Q����HZ������Rr����ʲ��� r���rxJ�6�cKF,��V�s�9A	)"�(M1-!R��LW3+�*����{��iHbf�p8Ȕ��lZ�L[�8HH�bY֣���
8�(6��vd� ��Q��|�N�b�'�u�����{r��.N�{6"g=���z(��ݘȾ6%K�k�2^y��+1^^%�d�Juw4>у�w�֭�� �Zj|v0e�Hq��:2�/x��G���^`���yz���t���A�m�f��	Ev��h�a�a�T�kP��J=�-5���H�O��Yh���rW�G�pPah@�������s��G�{�%�� .ii ��hN�����ڮ'3�{��$�2��:[m%U��|0��,u�eE2��ud���{�6�m=��C��$�����L�1gx�@9J٢�Ƽ��/����)z�z���7zϓ�&�9s�{�:��Gi���4pm5���.J�N��8U��8u1���4���uD�]ܘ����R�i��eɤ6�7OLe��$pA$��޸ږ9r�DA=��s2H���w��O�؏K�{As�s��x!y��G��� ,�7r��|� ҧV���-�2�E�,�_���,�'G%#��"^}���뜣T�ح�d�5�。��	�����1aO����S�m`�"'jۀ�5y�m|�W�I0&��(f�&�TǏ�������|���'�u�=�Yǟzi\��P�V@s0-�mYb$X�k�s�=o'w8�g��)H���F��G����_پ#�iߊ3Wa�E�9�ുHM'�F!�.� �����p��޺
X9t�#n�:�K���DD�C��0�����!��P��B������֨
V'�S�rm��ؐ-�W����&$�!�N�"��*W�[�.���A�O��l=�r�;'�����ސ+`�m|�(Q&BT5���B��I;C��cd�݁�KIO.�����a!?�Ld}��C�w��ǡ�"�~NpJ�g������j$\ ������,A?�ޚ�ƿ�G@$bx}~ڵ��k����mTp,�!����]oG"GML��ύ{8��Nt����*wt
'�o��T���I�KP�Y2�$*3����M�`( ^Lk˾��?L"5/�c48���ܵ*^��x[rޚ�~�7��[�0��*G�j�u98���3�u�g��}��	�\3pT@�]�F?1�~��=������쇟d��;�_0�������EY4�c�xC��z1�������#[ @=�Ѷ�3�ō�1v���Έ������4jTQ(b��É����omDAId����¸V�TF������Lm���9�p��sԒ*3.葘���cd =N�Ǟ�=��e�S�+�������ݳ��	u.�0x6�k�sL�>Kئ��P�/lo�~D�yv��d%��}���=�sM]ު�6F�5�I��8��u�rd&��l!K���������*
�v���P���=ȱ��v����_�d��#��0��v�g��6����Kc��+kc���;&��z	�C8�NY)��h8q`�������N�)&L�X�Ԓ&/�v8�^�W6��`#��8��c4@� 1[�8<��� !���!q
�#Ϥ�&������z��<�C���Bh^G�I�_���r�l|����|�0�c+�"c�Ə ��Gg���Ma�(߾�Q  X�=X�o0�8I��ʄ��	�I��)z�Ȗ�z ��W�G��
8�����gj$��d��jP2x�FF�����+��r%o5Û�Ŏ�K�.mK�Z������f��������j(}N5ӛDw"�o�s�5��r��g��z�5�'��G��<��G�Q,Xޒ��U�6��!Z9U/��K#
i齪�}�s�;��P5sVg���2sb��>���LW���%��V�f�n����\�~�N�.1�8`�=4<�f�}C��&��$���6��n/���*K�Å�@��sᤨ�`�F����#�z+����~N�~��3����K���a����=���䇑�zE�<�
��&�Q[��ڃ��;*	=kR��h&(���C��G�B�b�^E Q��.�2���=�D���v$<(#�/<;�v�s�_�<^�Q��#s��u(�S�V�EB��y`R��Y��������6�P9��>#��
T?v 3;.)��3�:o��(�����f����c�~��ݕ��MZ�2@�0?*K���%�:1���q�����s��X.�*�@f&
�U�5Bt)r���bB>�>9�GK��m�}ӧ�����hB��|�`����"��F��3�6����ϘI�@l|\/�!���'����n����������H�e%��w�<�C��{�F��
j��F ���.;�T�l��m�ҍ���\]}q��/ڡW��Q�P��A��d5K���o%�J����{��k�]�Q����P��� 7��������3�ȼ��x�[l�����4��y�K�{d�����N�Yy�����~0��a�Q��"-^Ƥ����]�ƕ��\��b`�,$x�m���1���K��HGd� �m�3�u/o�z����{ B����,F����)���+f'��RuH8\��Щ;��]��p<�EB�@y]ݠՕr8�F��D����A�m��K9�Q~��Hz2��م��"��g/,ݙ��uMs����5˹p�H!�Z/����IZƕ��듬M�o�� Vr�P���Ĕ�p�j;"��� ƗV�Fy2gf�q�y|^����򄸁�:�s��Q��aY1���WD�4W'?��be��w��uo�,��%�Op��S0�\�ew�]V��L�2�C��v�-�,��1CM�=q�v�3'��l+�*��ڣ3��{�Ec$-].ip��W�\Xy��/PQ��Ĕ��66�?�ُa���
|�l����J�V�ӿ���ä^$�����@S���u x�x6[{ ��H%:pꁌ�|�\�XRK�=�ȋ�<�O8�߇8
�a�k��FP��v0@��(�͆��D�5AU�2�5e�)
�'o�E��8Oc��F����W�p�+�R|�U��Ċ��=��8�ȧ�u6��6�g�`jK��i��ڜ	+uB�u\3kP[����L����~5��:��E�@����8EkľA���r�
�c&�kP�w����8��ʀ�]U95o} Q�u���Q��w�q��#�((j-�S���v ҈Nc>��s:��fu�,�w���S�#R�I����j�. PE����ice�(D�q�9��M��eŚ��Ic�HRYR�"��%��@4��B�s�����(�"�Q���d,s���F�{���J|}#�rs#?]}$:Br�?�§�N���f!;5ժ��~�L��S�|?�� ��J�]����3,��M�X,4�,�Y�eP�s�c_��_3j �L��D�ņ �x�Y�~�vl� ;DҬ�6t�`�C�}���f��;��h�w$ۑ(cLs3�ʙ:��:�w��}��RU,�8МZ���8��i,A/YnI�3S#�y�v[�sZ�@�h4#�xK\�hl����M����'�`������D7���0��YI�4��?�0�/�A?Y�d3���g�T�wHDbr�"�)f?�~ 6��*-c#�+���c\+�Rib�p���رc$.�B!�2��?J��n:S ��N������<���d��n�ҌG�n[���0�<&c�υd%��qy��O�r_6��sw�m�!���D��1��~7޷�̗P��?�9l�J�!�A����m��yP��*+Ղ����D ���;	�6��a��j���`@�R���Qdb��)�N8kd��v��(���֠���f�?/)�j���3���,	@�ۘ"*�yڭ�@�ZR>珞N�|��<'.�S��?�F�r`�&��� �Y�p������ �zRk����]Gvͥ#��w��}; Y��(������F"�R��zWJ�A�"�/,���|I�9��5[q��Jk�~ˣMoX��=��x�H�V�LS�m��� ޕB@���}l}-ȏ"�ق��,@�T��G�rS�$�G�A�!v�!X��˲�ë}_/э�y~.���c+���jf�=�K�=��rJ��	h���Zx��w7wr?}��1+XԤ�V�V��\���@.�������\͒y��5Ǖ�ˇzZ_~[����?@��]5�6,C�k��=D�W?3�XV n%zH�j�K�T��+��b���Qg� +��70w0�K �q?��@�[9ɝf��}��ב��n���e}������p�S@K��;:�5l��o�I���@�P{����5��76,3
�<�<���8 ��>� z�0Pn�뻜���R*m1E)�齅�� ������L��l��{2��4�H�M��a� ���J;�l���dw���v�t:d�+M��*Y)��?��t5�v�ŊֹO ������V,Ň;�
m����[ތ�3�	�k�?Db�7�(q���TF�Z[�Ô��ө�5���;#s8f+�HLc��t0��1i�TK�*�����N�R�u
�a��x01Ƹ�Z���x�|���Q-[`����;R8���g��2ϐ1Ke�����y�+m�17�}<;'}�t��U����3������o���m�.������T��o|�Ň`&<�?^;�����s��FE�Ѡdh<���8%qX���#�|�1A���3�������o'j�n����� *�e��`�;�]QZ��v`r5�.q�
�yK�֋ׯ��p�J_��`|w� ���'&j����_�CGj{�0��b?�>�4C�ۤ���DI�	�C�cp��dD��ɫ��{�����i��0瘘�� �^{$i�>!��o�Ș�֜q�ȅM���Ky������F4�[�8v4'�n��Z�������_Uc���}��W�z�B�;Y�_#��z0��
���t����N��e�Fb52��\v��#5Я�z#�_���F �ł�V�%f:3]/0�U}��f�5�I�����n(�v4:���><p��}�B��N�׷2]ϥU[��~�YU5,3j���1��-���P�ػ|&��Ki��OdYM%��d��5�ɳX�Cy��+9{�N�|���=�Ia�Z�m����íf�%!�pd�
 dDN|�6��u����
E�oBY0������-��R|@�a&SrmeN���+QJ�	!hC�_0)�o�[V�G@͹�ت(iY[�'Z��T��ĸ#ʻ�Ϥ�E����u��ts��WzF�H�>���@����'��un����f��r�=w]ǹ:���ri -F��eTz-�ӡ.-��Y�n���<��7�d�@;��	��j��2��p��}�ǿ{���=�ȡug��23Y���I�7#!(w��t���u4���MH�,�>�L��c�gDy4N6�4ܛ��\�_ȷ/���q���z����H^��'X<�J��������q�+���v" ~"�s�^�l���:������] �Q��q!xD`���#����ԦK@�E��y�~-��sY�>z���ؔDY5Ã��v�h�_'�Y���l���1�W/�ȷ�.$�kz��^��n��:��=�O~Nfm�þ�Ǘ��q+�0^��E�쵩�9;;��\_��kY��(����~�����@��_7�}ͥPx�\��.6J�'�NG&�a�вW�k���Kh��ﺙ�'�����Cv�����d�����k����Q)ǝ��K����R'��F⫭m�@i�f��)A���:܁:�����R��!�J�b s�g��F�z��(�?����k=����R����D�k���t�i+���NG�y�Z3���{#�R�ԧ��sP^k�~#��{Y��ɯ���9{uk  �zu�A�jF�tQ!���/5HAf�%��C\e�C�5xY� ����|)ST-��gy��wV�OD�6y�Ã���qb�*Uip���R82k�i&�Ĝ�:��a�vjr�'΄�=H��H��Ĳ���6G֌�98]�۷��{���t���0w�&;��@��;S;#����˰`�DY�p�H�����N���T6̠�+�{(�S�Fe�U�]eH߽޸�?��ڲ1����v�9g�3��z'��	�Mx\_ݓ,iz'����Lq.2�Vi7��}i�n�g�५�Aߦj8�Glr��~�.=&�	F|�AJ�wΑ��,�T� E
"-�T�2�|�{��W͹�WΞ�ص�x�L��]#8���	�A.���cx����+_�^Z~�|M:�ڪm��L&��5'`�THD�v�pY�"�����#�I��r���=e	�ݟ���by?[n���
`e�D662ׄ�J�a�#|���@��j���k�A"-�k���vW�(u����t
Y�7{Py &ׄ�
��Q��"+�(���b�����m<y����f�Eh��/rfM�x�^G�X��ӄ��󋡼�慜���֙\��d�0�!y�n�\U�l��g�Md�Gz�P�={O�'�I��+.H ��fb:�ؚ�#O���jS����"���Z�Vُ��O?�,W����/��V�[�QL�ahR��h
@K��ث"v�Cy��R�^ �!�P��8:	TAE7�fF�h�D��%�:���tt5㽼x&ϟ?�ϔ�l:�wj�ON�r:h�ӕ��L���No����ɦ�#r1�4����K�&�ywrYc<	�d.���u� H�v1�+У�SP���Y?��d�d)su"SuEm�˽"�Nf�ov2�@��fr��Jڎ)W[�a.b�7������p��VT�ʑ0���>���Mз�Y6�����n�G	%�F�̆t�� ��q� ��F��O�JB���q��:H䖬��:�㒱�0v�ȍ2� 0���~XBa�5�Wp�XoRgz�B2�Ap�d�J�DC��E��c��'� V@�,�e�Nk��� 4���8�4r �m5`E��^��=���La�L�	R���Uz�l�'-
�7� ��'�!u����8Xl��u���ckE�� $�ⱍ��}�WV��pU;ŭs�E�#�'/8G�ϔaO&����}BlI39D!�L}�e��=��4`��`�c�0h��֠��~��̮'3��:���a���HX�?��W�u� ��:Jy�ݴ�:a�鷃��+��=	�Eb�$����w 2k�>�N�M�j2�eTurkp������>lon#H�t0 �� �%dKrE��h�ͧ�9���#JkV`ck���~��2���m|� ��x��(%��٩��<�|�ɿ��{���4�]���9������-��~8B�e�M胢����/ O ���Æ��G�Qe��(A6��8�6�����hKV��g ��lj�㹼�,�O�u��\�5�s	x�s���ӹ��?�N�X�p{/��Tx��� s��y�Ӈ�6 <��F�U��� �ݩ3k�gUFV�QڨcE�� �1�ǭY�t5W����&�S�!Cr}�<D�]TT��Z�J��՚����T�#�����:]�^_z=Wj����f���2�UbfB���Qc���em=H߀W�F7K8���(ذ7b�:Y-�"���ֵ��dWBF��`���ǈ��^HL]���~�,�5}�E��~.71ǃ,h�Q(��KSy0ngԒ ��,qƽ$pIC�j���LS���x�=�,� q�C�S 8'��@���N����}��v��CE޲����,���2V�Va@4CMz�5�L6[2w�&!�e5�u���x������H��,"�N*�5�+4{X-���[��iL�f�ks�bm%�[m�W��QI�]��(qp4��|�$ʱ�7��P����5IH��|�1d�ھ����/�/���'��>6���rK�A�[,��@�X���S�%(��w�S��[���M.8#�Ҁ���(�gڏg�?}�Y�ck�hL˃�GD>Q���9fX�O1$�+bc�P瀤�9Ƭ6L@,뻉\m+� �W��:�����i`���&����U�ʂ|�7$7lpa}{8k��}т3�\7�j2��kh�Ɔ����@�s��K���Q�Q�<���Y�Յ�W'�<Pb��A���"��s�r�?��hH�T|oXl(�(�hL�{�=% �c'�'�6�d_^��-�J�UcDfK��*�^�S4��d#�(���(�0M暙�J�ۖJ��	�o/Ԅp��Y���,i��r�D/�9��Kv�#_7@��	;�˾Ȥ�V!�Q_@^!�U����!h<��9�9�]��(�x�iC���A6@��������&����k΁���=�FO�v�����������d��}b�88���(�#iIN���XJ�P{C4?Oe2�#p��ꕴ �״�lI���k��I1#��SDF�㞃���p����@e�/E�(�g"�<Rw O��=J����e�sѐ��o8G�ڢB�;�pMZτt�QJ*�B��m2_5���j�)��\�:����C�0�5�y8K��pl��z�8[s�a�.j2N���d}C������R��Fpb���6�ND{�#��9}�BJH�"�l���O�]�˽�i"���PJ��F/V�B��*Y:�����ꙍ���U�})?hF��_?Grƹ�XM��[����z�H2�Ń�Kj0@�@َ��H��:��^ �Xف:7�7v���������1��p���|�N�Dn}wT��&��F�Ɵ��?���ڊ$bu����m��:F�����a���n�u�,���M�P��YnX]cґY ���J�#K��� ��Z؏)�@/���8l%����,'c��| ���K�+o��#$p�<h�;q��_�C?z<�o١�A���zO�+�v��1��XZK��H��E�n�����	�u�.�V�xb��@n�%R�]Ҥf�}�Wn��2��T��7\��t6z874A�$2(��-i��4�`Ij��٩���S�� ��?�n}+�U}�X�9�\$�f]5
�NKN;�:�:��L7���R�\�)R�BX��=�[��}�q3�2⮚���r���G�b������SΦ�:ܻw���P��q�}�^���r�0���7�/��F�h��Є\*RP���*�KAT�jL��~��^�����}�y�\�)��5�@��p�Spg�S�F|�4zg�&�'���1��+�{�ki�3���8p�F\"3��{X��2"�>$���ȹ|N;�Ձ�L����0Dֻ�kl?E\r(_X�ƆC��;#� &=r����q�H�ʣ1*NX �[��e��	Q�UL���e��4��R��勗���3i#i]^�X��|�A'��D+����z_<��4{�Q%���CY06�*Ǽ2[�"��ˀ''�<�����zq���6�bU|MJVĹg�0G�G���5(��)����&rہɇ�h^�j�	�� cC,
�6"��4��{�D��ڪav�k�޾���>iÿ;HЌ+ ЪثӅ�2�'���3�C�޻ʻ�^�����K^��]?�'�F$!��)���T9�z�u&��&$�Z�����dpvB����5'k��Q�4|������]��iwc'Ǳ�N��J4O�n7:�=�o�kп��v��֠�ut�-J��������	���~��`���W��r��ZVz��Zg�(lT����hӲn (B?�ѯ;19I˒��$��j�"u|(9q��g"qn�F���y��NBz�#�U'�!���ɺYW�:�Đ�g����.$U��P����~R'��S��oU�$��F3�#y>șf�m�è��d�������f2��m�W4�TS�������[md���������� ��L0G�;}�|2�!z�� jhw�|��!B�GyX�T�iӀ;��(A��"���cYg�ʄ�qw�e�m��¹����h(�C��F��r:�1�	XKD��tY������	?�5�E�~oB�7�}V%fǨ������]�qz/���϶�b�p�g�޵�%Jga�2�c�S�����6�^{X|�~_�N�T%��Z��O��u'�Ib������9H��Sh:{]Q6����T��o��t.Ac|&�����[f^Qb��$jr��Uwއ��X�2���8��b��Q#��V{A��ħ����A�n�k�c|����cT	xqXR���Kٖ��V��P�EH�l��	,#d���{�ef�&L��)���p8��1����'��8
�٧@�Yup�́�f�rǛ�6W+���+;��߫PJ?rXO����C�m|'4�"����j8;�g�v��]d8  >o�qN:>R�J)�  ���2z�\��ͯ�L�������?����1ېi;���W�T{,��Dj���r�C,m�K�T2������k���=�h��U;.	���]̖r��+���&���\n���G���zx2�,:3��qL�'�N��CM�78l��$#��#F�lu"��myJ�%dl� H�zZ`0K�v0�"F�T��=TG<���N�l,W?���˩��r%�jFR�A��ɬ��'7� �ߠ�&+����@�(-u����Z6�E/�c5,��AŪ�]�����ִm�9ܳ�b��#Ya��,�sGƙv��!%5 ?LX�����l:�@Y���H�uٔN�RY�Z��9a�72/z�u� �I��G� �AUcV-��2� 6�ﺯא��ְ;����j6�,���I1$pgG.Г�i�����W��0�E|�d/rA���F;&���`�s�F�D!bN0�j��v�T���PUڟ��M�l?P��0v3C̗��}4���|>�O�EG6�eev��j����'�d%,J|`RD� �M�&��4��yݣ-l)���x�Q����� L�O�*@o��^8�N�@�U	�=!Y �zl���S�$��>�Hx����~`���;��-�8�~��}����1��[���B�3�9 �ז!8I}�2��q~=2>���G�<���!�\(�G������v�K�!Jy�{�ט=�^?rc|�o0{���0��<z-%j��ta�..��lyÖ��=IkK�I-#��g'���3y��}��nd�AP'��#D�u�昝����[�(c��Ap�'>�h���E�
��:�J0,$%Vvܭy��G����KA�1�4�m3 �����w1�Q��ć�ܸ�b9��ğ��0lcV>��$�WG|"�t[r��g2]H������m�����m�~̑��С䵘��CD'T=��5$I�z-3�7�p��i�e���@��Ym����W�-�r�8Z+0v]^H|v)c��"����c�2.�T���Lc]õ��T��KW�h�,�	��Y����"�M���s�P�k��Ո�+�FI�+��'����ǫB���p�ʈ}���Y��M0�:�Y�KI�j�T��B��)U� ̀�t��s���q4G��`�@#���(줻�c�7�1Nc�2�~�"��d$2n��	�HO�xY�GܙRU�U �O�{͸Sy
���F�(~#����)��(�V�QE�D�5"c��v��at�@Vs����|-�`Ҫ��"r>� 	�`wW�&O����m�K"����ι�t�Ge��M1�8jGBp�:`%XUs�g�E5���\���r�Z�ۿ�DS����h�K^�rwNt�O	�]Yp����H`��@�ۦ��CY����莲\���Z���L��I�rG�G� �	@_�����h?��q�����w�qG<�qI�료?��{�?՟'ism����>�2%�8����#���'\9���O�DB�v/�hh��WӔG�O�>���1�O8��0�^Ǐ�)��5_h���v�D�7�R:{U�ax�1��~L�������V{�+t�j�vj��h�S�3W��~kC�"/�j5�UD�@\:�sT�hiD��<�1�Գ������,˒��S�e��UY�Ոb��%~៘_��@� @�.gg8�;�ե�R���)�ٹ�#"��&A2?�7��"����}�i�,��ȖKP�;�ٮ���S��]Y���{�_��2�IN �Gd^4�wK�Ȫ��^��v2��oo����Zs"I��^��[�J�����ܦ��#���ȕh�]�g�/>�Ϋ_�E���Ύ�n\�����=�Y�6R9���Ԏ��z�lH�}Sqv;w�jfJ�]�}�̭P�{�o��	�[��G�in�[=�!�Q��X�L��fg� �`��S	L� ����`Y�s�t줡 ؅#-����U�5�?��i'������導C|��k���Q�6y��qc��ю�C�ɬ]�/��K�AOTr�^l������E{���c�*U�
@ۆ�6���|n�ն����X
묵�;��.ǞgF��6�3����WW�e0���\�l]����s�
Y�$0�y�Dg@xMV;�7������D�y��TU��
�#a��G�g��V�3���%��	z#1�y��l�ƻjʱv�����=l1k�r���` k�X��O�8w,??%SacZ[8D��=�h���*�-`� /w.���"3{3F�yw�sJ	3���mj�G6�"��r�Eն��rx�Gs��cۊ@����x��Uġ,;�s������.>
e�g�^!j�_��	!lhJ�``�Kj7T�����������Nj�w�G�ˉV����R�Y ��9����� ��e�tY=�]X�l��\�ڦb���CK]J|�h���{��y���XW-,Tl9?�*�朵
<�谧YQJ�5���v�&�X�&D�9�GH��ȦO_
|��L&{$��KS���7�V�޽�-���Z� �QP�tu�>�#s�#5��)!U�>%�ɋ��<�i�Qfitv� QF�۱�����
f"w�^��d�b��1®��t�<M\fp!�٘��N�F�^n�V ��	���iì����3�K�~.r
�ގ�?i7���V+����lr4�1-�n���'Gb]O�����&��mnf�$P�x��ژ���L�)/����;����g�EU5���g�1�����$��u�ΨS�JDNUz .&z�!{d6�53Ŏi(alh�(smk�������2\s�����K�����E�O��U� 2��b�̀Ơ�[p��&�=�-מ�e1��ܸ_Բ%��/��I1�e��J=w�p	���/ܪʡ�Ͱc�-��b��,LQ���8�^����u����f�?���� 	M�*�<�w�R�����M�UQ?�l:a�+
V@�8�&��X��]N
�Ԟ K�������*+����q�ʄ)MJ���
'��:�JBD�)��B�
��-��/f ;h��v�xN}5W�kSS�	{$�8���4����oDye"�;�Rv��b�)u��Lf��@�>K���	pÞ\����ޝ�>���ڂ��O��hZ;�1aE��DE2� ͫ3��!�6�rčh�*�Շ>����_����C�i��,�]@�šQ����������y�eBU�Ю����HɖD������T�9�VB����å�s	��k��������Q�����9���g8<����D<�6�ޒ������:�_���&�[�ȹ�l�(�m+Q��Odv�>��y�a,�6Kz��砟4�ޘG�H�c>�8����2��2�Tߍ=����y�}d�������RdL-F���S��L��b���u�6�O�x����2�Me2����rF�?�֔�Y��3��st/��t�Y��Wk�Xda|�*��� *���%�m�9	.Ⱦ�?�k�l�''�����\�����]l��!x����+�ƀ�N�l`��P���ar��!Cp����
s���;���a�7��z��;����bɒ���IO�v,�rLmI����b�m9�.��AǱ���SG73����C��FU5���g�w_k\��U�cY;sǳ݇��;�h��c�ad����7F#���)e
W"�!�5��q�*���~n%);����ӮM�Y��^c��C�b��rYY��F�R���#H~�k�5qqd�c�D�y?���{����S�����|\�r�C�n��MW����2sb�|4��p�)�J�x�\�_�lE��2�4��R����w3�S�1%��>nY��녳�!@H4ۜ	;�J������%��cO��]H��<����LH��:6�L���mőC�\~�9����v"Au������@aeSY1o>�d��n���@�淮!K	�y�x������3$1��^y�H�h{4 ��5o����ߦ�0F��S�R wG�� �rzn�3���ݭ-�Eu����]�U�~VDU�Oo�x�|�*>ۃ�h���_��s�@�O��(��ۥDNr��!���)d?��R�z{ݡu�=D���bC��9�V�t{y����e��P�D>"��-��&��O�4�,&�q"n$� Zx�q��k�l���vm�a��ɰo������F؀=dϽli�����s���쪩	�V�����szɈ��.v�i������)䢹��e���bG6���b���]۫��m:�Z����ڊԑ�E��y��9GK�4f����uW����x�어�[8�-2�X�~�6��P1��B�*��Y���H U!`���(�t$b��G}�4Q���,��_�7��Zδۣ�W[���{�p��%��|���r0r�����,g9��f���ӶkkW�HcHvS���"r��:��q<jԷV��m�[o�^����[f�^�������(7K��eÁu���]c���_~��6���\\Zuu�(@Yd�ُB�0�u0�a8j���w��P=�
���Pn���a��=EŲ�b;Df��r2��)OP��Q+�t�xeG��3�ý(�BB��Z��=C�����]N���v]��4HI�d��6ć�|�ѯ�F�!N\t4�N���8�"1�v��;"=�DqR�uH Ĭ>��}
1E���z�Y�c$!a�`�y!P-�*�8�<׈_�<�pRs�m�jL�7�8����M��a��|=��ͯ��ZӨX�����>������B�� �=�_���uHt�t�X	�l�A��nZ������@���v4,y�=k����@{�ٰ�5̏e�Pg�j�55��b�& ��������C�ˬ��[��DqX���"zR��u��B �"�c��񪃃p�����kԞ<�}H� �X󖡌}F�кP��Ɨ����x�!��8���ʲ�Ljkg|��Ў�ω5z� P鐀�"@�ѹ�:5��|�d���O�͆YK��r���]퐩�;6<;�e�E��W}��5���X��p,���bk#c�͓������h�+=��Q������@Kr����@6�#���7�vsu)��i9苆�O4>iO���cc\c�6yĈj���<�j?@���U��~�x�S����ғ��������}��֙�m�o�$:����B��Eb�<3�� ,�X��v�$	�0}S�t�%~��H`�P2�َ`�(�]SK�{��V�m�꾔j���V�F�H:��m��Ń�m"�;>{iYf9������-A���Vu���z�u����q���g:8>�{p�dM���[�ʸګz5���i���m���rU9�4�Y���)~��tU2�8D��ω�%S]8sY���Q�j�3U#�T< ��E�s6w
�ݑ+��)���{8�ޫ
��`]���Sѐ<�vqځ���A'EXYҘf� �*����y�6>���!�j©�gU�8�m���Tm�����G��������C�\�|�=p���c`\s�E�M�u�#�����N����X�b$��0OZ�.�C{,���	������N���=���n�p0�7>z�-�F�6��q�����'��?m�^�v�7���Q�Dm��zM��f�H�s��eN�s7���r�^�am6e��,�<Q��|���|6�u�	<bO|�rGM*�h��՛�6[.,z�����b��y�%{�{kùtk'�Q��0��_�;!<�}0+�=�%���',�a�8ӹƵ^�V��綽����܆��=3�����m�|�s|���ikd�F����nve۽nǾ�6;:a�/"ko��s8�)����|�u���#N�p�J�,�S�%f���*�j��%e'b��u�=�� ��H��4:�ys4������Pv�=���&�&����N^���~��m(���]���nE4Q��u`��,���vRͫ�n�#�-�ؗ���K��|��٣�lr��r˱@�`�Α��/6#
�U��WM�S	��9���Nײ�D}�=�7�u;iY��Ot�7A-o�@�����������M�i����>;ԋ�{l�hl[�˩�s�o�H���b!�YQ�F.O*`$y&'�b3����\8Y-���>T4x���oO�t8���Zε� �/����}�Ԭ>"Ǌm�X�B�ZS"��ry�P��d�<r�g������jrrd�x`�����M4Y	۴!�!������kIX����}�}���}���%�	77�`���
	J��	���ep���t�c��;~�O>-��w�C�2�Nu�Wl�6�NDjEF��l!\��#�]WC��n*Nq����U}�%H|R�j*�ͨ��4S�(X�d��A�4!�����������g�nT�c"�4ϯ5�F;�}�������)��n?_��������k/K?��>���:���aG7�;5��9�v��2��_k_ظݓ���Hh��x2Q�U��bc��o�Q�Q���'��d�_`j�����]�P\��ùeD��gv���9�Y\.�������|��������fx]ʺ��u��۶��a4z;+�<��X�,퐉Swkz=�Ѫ�[�PZ����~'�����"Ѿ'���ڋ���zo0�Πk+�a>���9�B��ŰW;0&9�{=q�a,�u�N�^r\�#`]J��5��L�!|��d$�nVc��#{:=�?��ޖ�W�_o���
�r�ǚ�^v�ʠ3ז(suST#���1���Qe��yt����߭�^��Em� ֑?0��*�|�B�"v::��Ｐ�#����w�,[�@.7����8Q�Q��5"���m�tS����Ѭsx�Ǐ� '�<�c�<����A�;�J�J��L���a�Z�>�i�[�`����@-K|�!�co��[K� �{Q�2�-��ms�@X�Y!ƀ|	��X�Bs�+¹������ػ?���;M8���TE�����`+����E���@Ӕ]{I[�����Ԟ~��գ������|k��)c[��o�����Gs����Q� @����h�r~�>�f.�Ӱh6�F���zX�2���
^}������A�ʡ<�����WMp�{Ԕ�,[t<����wv6=�w�����|'u�,�x�&q��"�d�ă�X��^5�x/��e���̢�B��Z؋H������F�ո&�i������I��)e����zY��r	��d"�m͙���<7�NR��4^Tl	��.#L�>î���a����CP�@PD�S��KP6��5�9c�ⶀS��%Y�"d�g���a�W;�X���c}���g�sG8��!7�\	 !��9�kd�9Sg<���=��P�D�_���U9��3,:8Dp��L�u�}�=K�k�am�������d����Rj<jG6G�Ktu�d*��>2�N�G����$��ߎ4��CK}�N*�$���p��jx�G�&��
Z�qZ�)���J��әk��y	����F�M{#r�ѹ�9ڔ�����͕!� K&�OXC�I��}$��`<�r��$��uҶ�L]�>�Ofĸ��!@�)h��a/8ּ�g�Iz�.��*�p��[3s�P�����7 �|a��prkd�\�5}�{�a���mx�m�*w	������W�N���M{�_�ewa��ݶ��Ng%*�ثM,5 F|��n�kz����V�j���J��w�V�^s��$"]�_մ�CMY�vh1a̬���͞�e���\�m�ϿȳO�f���ja�8#��E�y���c�$��#�I�sdh�\��mM��=�(��9u3���[gb{䒵Ҁ'�qvX��C�u��\*J덓v��jZ(��KhV�ͳ�*�=2���~>Υ�d����o��A���&���<99�W_~eg�'v�u!Mt��2���
۲�m��T����̅��p:�@)&C~�Ђ�6i�㑵s���VH��k��*o�?��Z�J����k�~vU�~����Oڡ�E�F�S�R�b��x(v�2*��R�����\x$#`�t����(�YƁ�ß��HQ�8Ӛq�q씯���0J[�^�^%�DYܞ��4`�}�J�3Zo2�6�v�d}+��R��3?��&C���X^�ʝX��3΋\�Y难��c��xl/_��_�m��z�<[���p��ٵ?bF�����7Q9�[���'d��&u��V�E�'d�k�����0�"����uI胯lW��+� �z~bѳKY���'���'Dmu��*���a#E+��ݝM` G���o�msw����>$9(�Pg6E�OG�Q8fۢ@�!���SF�P9��-���K{�����&,�Z[U���Ȏ^~���Ӊ�e���l8Q��o�����3�؋���.�5^�v�P�Х=I\�Lc���涺�v�KfF��[F��ٌ�6<:��2�O*����cG��o��`�6����+	=wkS��^^kfy'��N���Q�'�;B���Ԣ�swq��jc�ݠ���:�������y���/��ɅU�9aR:AG4	M�z�X�ff�t��& p�l��xT�$��y�x�9�8{�e�b�4���f��V��S}��~��{ރehH���D���_9�R�E�J�#�A�����4�\���T|+��w?��Q[:(f�i������I��|��1ٟD��*�I��sx4R5�3��w��V��&���o���ь��؋_��W<�n��bZ�������m��J��C�-^�*)�[ym-�Vcӣ	��?���E˶��s��vv�ą�ƓV�}D=
f۬���K�i�t}�vK����W�:�Xnl [+�%�U�|,��w�%q��u������G蕹�X�{���T-��&�c�>|���/:�)4�EM4��(�Q4k?g��h$5�7�VkcS��� �1:�́6t�4�{8g��)iDd�L,-=�pm���[-`f�ޖ����K� ���*M��@g����Fi��k8�������
���P܂X�w��Kӳn� ��_��K���d8��^�b����Q�<w0�`ص���ru�ޓA�bX���V-��6{�!H@����y侦&2	pp��iX�J��YWu��x��)�	�6+D��{� �],WV^��q\��ӆ��!�%}l��郓�e��s�$��Z�h��"�'j�o��9/�Y��Fyk�/m�_�(�"xI�YF�����|��:��WU��ᷰRm��:s�X�x�*O��b��,`��@G`\�mL3-�Q��>C;B^�|�+�S#d�]�@�� ;{���a}���yq�+?����<�L���ښ��q,`�n�"��D�u����&N��Z.�zVfp��#Xg:<d�h��3P�1�p����@ �'/�?�˩��3��d�f+K����AF�ｏM1���[���ap�N��}�PғʃT.����pⳲę����⫮�s֦4�V ��h�c��4�}�ĕ���T�#�R�fadO`���� ,�\�g҃�OwZXwR�[<�����FA�S�����m�ąn$�R�S�:���w�q
�`�4�2M�6]��������E��� 18{��zjs��-ߥ땒�����Q���}��y���~�\Y�J��=��|m��ǁ'LBh����Ke���PEIu��M����g�̟��v�vb]ߛ��${ӧ#J29􏚬�#J^�~� �b�"N{��|��N�>�
�;wNg>y���-�rr�=�ᰤ��n(�V�Sv��P�>���tP��V�cԉf���I6����{di�9���!�4�H�X���tN�&HC6�QO�ȴ�v��F�韈ЅF�$��H��I#����f���DI���2�ա��U)�5q�%8t[�X)]K���~���X����7G��lh�8j�J\�L=�̍AT8�Ǜ��=�k�x�d��x�tnߟ{鞳�	IWJIb�"/if�T�~�Y)3�`�ɡ�f�
�U��̉@4��/f��5;n�P�YZw�Q��rnn��Y:�s�'����$���8>/Y�@U�X-DD�s�N�%ub fp2���<�n�bcՁ�'y�٧U��[��:�kLN �L�<\��,�mV�b��M�� 3��F�EuLU��:{�cݟ���Lao(�J�De\G�˩ą��X&�ׅ}����v�&M��M�h��Ye,���w�uK۪:Lʠ��7R��b��)`!st^t�7J�^^I�~���������K1��$�����q���p���V({�팣���Bv����Vh�ծc�c�'�rq��^iO�] ;�q&��HH��s�J�����&�TK�eU��X�I��aT��S��J����Q�י����9��瑓���on��n�cD��6&pFĎʯP�c�ׇ��m%Ǫ���g���������ݥ] x�&{�_���[�{[vz,B&1e����P��Y+�x ? ���p¡\��jG�@�ث�ֶ<ِ�Ϻ�)l�� ����	�����Y���N��ğ��@�<t�>��M|Q��Y�&�z�e�? *i�7�!M���H�G�C6��G/��(���I�P�ٴ������#�s8H��q�%q4+%O	��2T���(Fa&2	"xK�ΐ.r��0�����	���_�l��1�L6HUֺ%J��@�B
�t�X�����@��0�|~�
[����xE����i�c�q����{c�"|F:�ک?xm�ɉ��Sd�II
�1��^=Q5�6L؏gƟK޵_{���~6�w����r�{r9g���3��0菱�b�C��o�T�B`�>-���ֳ��i�>BF�;�*gW7N�S��c]�|g?��v��0̄7����9�(� +�o8��Ϟ�wL��������Ж��Kd��Hn�ZU�c$�mѲn�A$5��
�ܡ�`��F 0ku�Իp|u�,��G)�q����U�-=��`0+�������_<xν(Gm�V�s�="V�G���&x��Õ�!��-Y<wW�s��!+��t���S
�KG�U���d��f۱�_��ɶ�oW�Ua��F�}xJ
3����/#Ke��/𺬞i�L�,��>.^s����~6��X�Z"���v�8��U��C��3x�U�u����6��������G����v��m^i=X���@��u`[#O�ą�_��R��M�� 'eRC1�(jHpM��s���|������/���x�[͏�֚��`D?��2���k+��GC{��x��-قY! ���h2>��b��#^�z��X���"; ֑�M故T_���|�p��,i�'.�����V�3T:��s���x���$Op�j���'��?i�^�%��q��*A?(	6�Hb�_�%Keb	��B��68�F�1z\^o����9y�x�}V�&e_���p�pd����%ϱɪ6��ʁqM:޻,�M�<8���НH��GO���7K9lV&���*���HY��ptkC��� �m���+I��o/�OcԏZp����Еr�i��68'���� Jm���C�q��A�a^˙����I��*;~��� -޼�a;��o����~sz&��p:��|nW�Z��=�}z�k{��=9���o�i�lc�K|ö"g�R���&Uk�#we�-��&N���9�L8�M�T+�+��t,�+IӒX&�/��w�ۮ崷Xëׯ�`rwX���0>���R�#� 2�YA�����3����l����cs��j|��������6G��z�a0ȲrȌ�ȝx��N����8�n�8C�����z��
�t�I ��օH��y��>=^�g�
������gQ�ڲ~�w O��LcG��G;�g\���ƳV�l��dBWh�%��,Hfr����1�	��\j��E�5�@Ms~[����YV�{C�I�Z�v8��H���snX]��Rr����P���@ZV|�T��{_#ΰgY(k*����r��\n壇t��{e����r	��M�C`�+�m�"
T��o���qV^NOԤpܮk��{s�Q�FR�W����&�$��N�׎Y-�|���78h��]š���{US
�ho8�����f�`7	�7+�Ifp�/<&BQ?.C�T��S|��r�[���û�k�>����߼��~��?S��÷���_����6o`^_���&�J��XO�'�M���ř�n��W�(�&|���͘q|�b5ͫS���/��	��G��>��'���rb��a��{2�#[�8�����>ph���CSB	7�=�C����e�z��fѳu�0��F 6���A��w�D4͊�#/�$���G\�K2fɨ(c�� �S��f��Le\���V��&T:x�Q7�!2a���fpL݀��oɰ��:�Ӻ-��#�}���iQ`���C��Q,|�����3�#��}t��:��8�(���!�[�����g6�6eFB'��I3�˟!��p��/�	���>�����Vñ���z���ՄOH��� 8�B?�$.�|>]��ke[�C;�i	F�Pe�q�`4c��[��+R>d�Cf���\���]-e@�����Q���!k3t2��"WC��cd�my�����=©��x�
�q����)�:�
�X�nZJI(q�r|��5+(1�9���@CI@P����U��9;e�ބc� 8��=>�G`'>d��6;�yaґ'�����`������_�
������4)0�>��˯lttl����Hc`:ۓ'Ot��76�8���~%�!VVNP��䩏��oUrow���u������w[��\�=����xM�#�ZnooPά� {r|��#��{]!��z"X8���+<b]�O����N�2�[��3���1���n��m��2{�y�:r�+�X H�Y_yI>u��Z-�ʖ �?�#{���֙��{�Sy����d����7}a�OG�p/�5��i�J����p���&��l�u]̖r���	�x��F52p<���K�����8�%����f«X�Q�N=����2!��v<qp��JҾ���������'{s7�D�w��Oֆ����_ۓӧ6����q"�|ly���
d3��b܎���gώm��2?��b�DB�$`�QW����D<U���Z��.@�P��x�X��O�����t�F_d��(�בz��.b���Kh�vf��� ��ތ�y�������K*�/$�
C�쨍���ᖴb�{�*��V9�KR]b�[W0�d�0'VO���/�k�C�J�h`�>���O�P�s�mʢR��I,N�C��-BVV¡G0�G�o��9B%b6+7�lj'3����$�L�@	 a�`/��ڔH%&3���8ʖ�ؿ�Une��|���#��`d�X�.��J�(o���g=90�@&pn�|#�Ӱ(�U��m&|��U�b<�F	��
�XG���y���ZAO$u!��@�Lw��E솇륌��� `���˞=�P'�8��UA�['Dβ�{�l����Y
'�c�2���g�m��v���p�F X��}��ƶ��/
@kuT~�S�
U��J�dW��[�l�8���i���V�Jש*0�:������=�9s7�Ш�>��VLi�z��:-8&8�/_ڳ?��������F��Ȓ�B��N�퇫3d�O���!~�@s|�����7D�r iM���:=:�U��j����p<�erk7���[��T���������X���z`�m|dǟ��!^''x���6p�l���_`�綸�P�����A�1x~f�ڏ߿��|�Ԟ~�ji[�A]o>H�����?��)�	��g���6�{�p��nV3K�m��'�Lݳ'��
9�Y/��{+%�Ao2o�Ɛ_�iA���N'6D����U9i��m+�ww8�q�x�t�q4��}�������=`�l�<��A_g���\A[�0	j�jӡ�⟁��C��D�č�5^-���X���9�;�9`���^=yibM���g����ʩJ�3e�؈	�^���+�l��.������O;�III��$V	�K$��
܌�5Μ2�l�`�V���w��r�̃���C���D8="W$z�3╠�N6�DV��
ԏ�7jz?z�;G|3�MR�r4�g�I�{���L"Os'�h������$�IL�K�������F�
��<׌k��;?C\cYʚ�mJ쳅]�9,�m �=������Q�tA����P6?d`����2{YTԛ\gf�x�.1�r�<��[-�>�)1��x��8ݾ��4>ƹ�5M�ϱ��!*G�}E0�B��vNU��X��F�����C���&�nt���LץW=X�&]QpR@�=�a��5ƿ���0~�rn���,��_�Ǹvz�r�hb{>Ն(�	�#f<P��%p�Ds&�,v�0�"�+N��_���v0�D3+``���^�em�a������V�۝��U�2��b`C��e��6W�5��w^S폂;Q`R����v(8���m�~nTݷb��%ּ����
Ed6b��u9��0���n���]]��wt~�gi����?��=�9���E�Vx�o���H�cj�����֝��2�'���j+FK�sd���bϢ}4�dԷ+8]�S�ݮ���Z(�۪ȑ�}8R�4�^L�=�?=��x~�5�����Y>�����Փ����ɉ�����Z������PP�ɋ�v�}���u�{jy��FcY�77�B�M���&�k����2w��(�q.q�arj��j������ro-��?��Q�!5����Y"�>�7!�ܳg/,z�).�o�ⱷ���m|4���c]��n,޻@N��q0G��N���h��K�3J *m)	��l�a8s�G"�I"�=�Y�2��n�e�21�dq&Yl"������������^o5�>�gb�2q;K<B+q�]���WF����
Kֺ�����C���1�ƙ�&�;�/�IǢ��>8^/�;�v2щV���j��o�Xݫh|[p�C�K���bn)����N�K��f^*r�9F>�����&���J/
=��SD�,�I<F�f%�X{���,k�מev�����w��W6#b���ʖ;���(3��Y����xP����XH[6����p�v��t��������x'PJ�4��TH?�Û�X�H�g��Ø�P�!���z�m�����V0jk�[)"f]d���<�E����&����j2�U �`��~��h��%'S˩p�]���Of9)o%����(V�� tM%8d!KN �G�N|����E
�'�_�t�'�`��F��Q����M ���7�\��7��3�5^o�v�Xa�ֶ7@z<rpN�x�$�S6h#�m�7YQ�1��7(Ac��Y�r�{^�+�sXƨ�G&?VX~�u�/�o�9ml��X�P����)|9�@�NL�e��� �Ќ��j�T����X�AuK���;9'�����8{��5)?9���hS��νM_�%�V2칓��i�S�J���㛴� ��s�ݿ�+˖38�;���4g_sа����k� ���
�[����mA� ֲb)���g���A�'�o��ى�^�ޒ�i�u��G�CF�����
���'�0@��9����3K?�Uv_�Yr6�K�'c�&֍ҷ1���^�ї�%J�bM:y�J��m��X���E��b��Q-��\���֦�l`�lr;���5�&t#�ݝf�Gþ~2����.�Zu�ϋ{����t��A.����Z�� ��A�*Ϗ#��@�$��0u5��%��Cm�Q�2��ԣ�@	�3��n��� �������6GR��um�`G,���P�w�EP`�i ���SVX%.OV�B'�
���b�v�
d+�&���[ǚ��Xڏ������v��,�>*s�W󟕵߬��Ry�h3�&o�::���{�u<�f|����~B�R)�+$ez�Q�f�O{fW�n=�|�|W૝�F}q�=���_ps��za���G.,�Z8�){�$Uaٖ�31����W;0�r$&0^i}�2/���)��(9����
u�9��(���e���m|���>�}ƹҹ�֥m����@x��Ħ�Q�X���] CnS�ͼR��I���>Ti�T�Ԗ�H熷UF.gE��)?�)B�F����!?����S1�Ͷ+��{��n`��>y���>a�'g���Z�V�.ȝ>�+eba�լ��O���g��!���w�5ݣ�ހ���Abb��"J��r�=
�TV.��Q��e�H\_[�F���YSԇ��-��U�}���;v��+�'#8(1�k]��@@���	�ߔ���ެ��)�J}���X�%�L86�鐓�2/�.����ұ�u"C˷�@�g�1���#d�#�&�
������ ��,v��:��ݠg�8���n޼��f����x<����׺�.�#����jL�]�D�W�V��w8����~�y����)�}����m��������O��tt�ho�~�[d½�Ⱥ'9��c'C�`8��������X;�s��A-�/�(T���$1"d4df�o�������{��S"p��]��M�Z���u㚑�r������6X��q�E�Uk[�,Ւ�~w�=�3`y"T~E�g`j�'��r��a��a�l/�]yo�$�z�~A͙�p�sN� *hOO,A0E6?&G�^�>��C ݲW�>Þ���wo���\{*bR*gU���I�#���ё&G�I����x�#�nWn[�Pr^d����p�|B�c�)K�����S��zχC_��)�w�R�6.��Ot��7ܼ�L�a���ytﵴ���<B�&;��@�$�����ѝț�pN�z��o�O��%E-7H���"��ҥ�gW�7���0ݧE�HT�S�f��Şuf8���h�D�6o,B�$w#O`��T�������T����V�ō�\����y���"3�X�Tf���|p�dS�\���k�X�u#��D�餒��ahJQ�F��Q·cb
���Y�L�kg:�5�[B�� ��*��s��$���u�Ū{�L�!S럞�ї_X6X
�0�A?O-�����^+{M�'v���m��]v3[�ᵝ�nm�L�(%�>��vT�Պxr4�/��uN�6��拑Z����������!���LA_�vX��8��C�@�*O�qN�Ֆ�2��m���9�	�b�?㜺J�����W�[׃�>����K�~گU�L�g�n[�>���hS��Ճ���x���^�"��U���8��ȏ0`�p�WN���"a����<���)��8��9F���ٙz��]�.�\��A�!`��z~cw�����u�X�r�Dk��equ��r[�`�{:i�"���V�,�[�Y$u�p�w0�H����?nGO���k�a�Z����:��#�dj�Q�E���9�-�{
G��R�o#�@���9���c�D1J�Tg�m�T�A^�&r{�����j��>+Xt<�m���D�uZ��z��|k��/m4Y4��8N��Q`�UA���'v�쩂ׂZ|]f�̲%A��H��(�1a]������hD���E�em��x =_��x�կ�g�`����v��9�Ǎ��c�[��Lkc��	��cy���'��(�8��O� ��.����~mؚ���h4��njڡۅ��	�8~H�2�񋭪Vh��XP'���C'�q�Gt�yss���'RB�ff��K���?����Ǐ�hM��.��<��5�k�I��:q�T�Y]k�@F""�j��s8	$�f\s�Ry�Z*��d��Wt�-�ڲo����@ȕaM�����m����\u$"�2̑VZ	N����B����[���B���p�,qdj�=���'g_�s�![c�s�L5��)"�铧p�	2��"i+�?oƒ(�Q V(����N}@���5��N�ǚc�x��nߝ����?�.�����!���\�Y�Fܘaѐ�󽂱�� �HN��?"d�p$K���.�����6�5
6e�<�,������d�E�Ӈ��i&}8"��ڛ��~��[�pq)�:^GU;PI$C�Tš%$f4����i��C&>�TvH�m��Io:]򖳲$�e����ɑ�����.w{s��v˵uH����O�iL�D��D�Ӄs��C�?G�8�>z�D����;����S`����ϟ�~4����A��$|�菑)ท.����|�̌}cfuww7ʼh��,k�Z���
k ����JDBY��|�?��Z�T޾��'���;+7�����k��+��u_�X]�j���
I�Lr�k��!�)h9
���S�_��.�涼�Q&���ϑ�[�����Ҷ��I�"'@��8�z;/E����>�)Pa
p��c��Y� %��vD
T�9:T�½��k�}N���N����W��Y"؎��w�k��[{{ip�'��zO#�g]ح\:����)��Ȫ���=kW���K��Q�ؖ��;ti��Μ�܇D�gu� )C q��=����]�>b?�կl���]!�#>yq������U�î�_��t`_��ͱ�$w"�[�h%�k>;��)+c�������&��5���K�=�-3����D�R(�m�
-=<�O��?�Aij�S{IX��ȝt��֘�%U>��p��QU7Z���EҺ���4$�;xå]����T��>:���
3�p�Vcdx��ςfo32�2}@� �Yn���ޙ�:$XI���k�=��>gV���m	���%�aY���j���1����a��������!ˠ�X&��,D�-M��\���91��������,����ŇKd�9���FϞ�ӯ���/����3{��G�o
��Lk�ӺÈ��������� P�Bw���Q.f��=����
"���I��>�r]�bͲ�^B*IC][Շ^[�b����3��&��^F�AX���Wp�7Υ�ͱ�G�.�q��z)��~�kў�]�0���o�z�ڐ�
�MgØ��]�.����G�:>b��5��H`�������\���>�� e����I�K�&O?�yrG�rOP��ct��n{α�8��'!+��%C:�G�yb����f�5�T*�R�:
�i�S5��ʱ�5�x>��������~�	`�pH9SN�$����$����d����Ӽ♯��5���K�� {ne�s�{A�!J��s���W�{8��o���7��,٭m���n�w�vY�����V���ى2c�f���w��p0����F��W7��;e�������r��ƪ40P��?���~��p"G�}����Z��̾�`"r�3���Ap<���=����.����A��M���C���̴O&+�F�d+ǁ�i� ���*����a������LV5�Sf��V pOGZ��幟+������ɫ����3@�:�<̦��"�!>����Z&87K�	�޽���J��^�xR�>`��	���P#}�9[9p}ʜԇ:�=���wx98j������)����(��N�MGЊk��S��㷙� �CY]�'���:�H�Ձ�2D�4pI���J3�G���0���hL�>k��m�
�ؚ������$�ϫ�W];�%�����7�2n�&p�� ��$�.Q�Q6��F�*���6�'g��0q�pHl��d���o���Z�ȴ����7p�����h��)�c!�XU����Ҽ�ė��a�WS�L�C=Om����3�-�8��WB�2<��w,���WPY��<y�+8>RÎ�	Na�DL3��|���6��i�\�H�o??�wm���w��V0�Db�pbd)[ӈ���$#����삊t�a�ĜM`�v+��"G�
�A�f0\ǟ޾�7d�c@���0�@�:9�Md�vW���Y�Lf��J]^�D�� ̙M6�څ�4�C���@�7��+Ϋw	J8HT<>�ݼ{o"���L�����9	h_?�mJd��}`�[`��s9[��T$����wU��Cn�+�2h�����PU"�Yu��"j����z>�)�%�5V$N�/%�lt8 D��x���D����gpb��_@���1#��]��V���� �}�Imy�F HV;6t��HbC��W���0���s�#s��o�:�\�۷�z�@��;���  =�T,�8�x���ji��K�n���ֶ�\����|9?w^�ĠǊ���#5�S��VVH�B�"2R�R8)�M�R�.q�x��L�@	{e/��R�l2���X��}��{�D�����9m郧v�V[���$�;��E��gE� I�W�e++s�V��{_��J��u�]����^±�~��>�\JM1/6���se���l���$?�Q�NO��%�=�%e�M&���K,�o�����N�4_��k�i� O�q'�(�*3Otmd,�@������S��G=�:G[5|�Q��lJ;�"'ri�&��'���,���ׁp�.�1��-�gܣ@2Ԥ�R�a^��O|{�MS�2�C��j��e�sX����K �rp�b1��q"��
�Ԯ��jƹA�GN� ��_��.����H��E�o`��Ir�R+���q���^�x8��eB�T[|к�^�@��pM�(`T�}�:޹�i:��e�|n�߂�b�y��B
-����A'Jz�Lk��5�e�M�HRT��v`$�\��LW=�T��|~�w�K�{�7
�1�5W��g����/X���8_㠳�\�x=d$0��ז��;ݗn�qT��?�V��O��4�"� M'ic��]�y����۵0F�& 6Zg~f�MT�Fhh4=C/���`�G��C;H��瑝���ad��39H�i,���{8�7�����yT��RHi���G�������S�.���w���{X��;dA�F�jQ�&�Р^߈rU#��k�孮���nmo�D@D�X�b�]�m�w�C�� ������:Y��z1�X*�^�c�x�S����\�����]�v���'�$&¥o񙉾���ť�f��5*�O���o_[kŌ��*�TW��j�[��?P��p���r����s����!���Y"\á�:x���J�yYx��;\�b��-���b9�g;��f��3:��F>*X��b�G��qϳ�s7Ezztjk��ij)�Սs2ԁF���7��'g�t|�s�Ɉ	1H�=��e!'1v��/.�`S"��=� y���R���gn��R��'�Y~��������_u��p����������$�gl�zZϝ�W��6�VG�GV����A0u{~��94SK�e͈�WOc	�$���w�o}�i��}�=�'�O�J���QR�����s>R��ƛ�὚��2�z������R��9u��$q(�"\`�\y_���� #'�'9	��As�;�Ci��X��}�M;QN!�S�J:��ၸ��#ߊ����ػ$8���D8�2�AH;�~���:�)-`��6�q�(:̑�b7إ�n�_T.�N�@*�w���B}�Lj�Cx	���1�^�X��|{�S�7�/�N7Y�d=��$���奌�Mwd78�KO>�J�|��9R�#	N�)�~f��^WF[x8��f�+�d/�%f�eR\�N��a���W�"4)3��s���6KJ^��y�k��������L��tV�G�S����l��������E>~ػ
l����B��oH[9�|���0�m��?$<�L�m�iZ2I�wz p4Q�����H��(ej��ᰴ/q�	�J������Hu"U�XE`u��cK��F��k�]�����S|��mʈ�jcdB����c::s�F-ᘢ���O:l�BY�k�
Ҧ$�Q�E3�"� Y	3���x8�^!U P'�s�K�*���R�D��c\{�����ou~iYw-n�6�>��[�����#x�{H�u�W;UA�R�#𗎉�ى3A!sKD��l�����8�+��Є�h�P��]¡"e����u��C&��l6��:�L�#�I�߾�����YbG�� [kK�q�ly�G<�����`�	ǌt���c�|?_��^��j��� ��)��`�jM�V�r�3Nq_i1iw� #���� �F��l��d�U���
װKJY��7��t�Jy.K�^y�ʐJc!%?�=X�z|����sg��3�Y�X���)G��������s��� �z�	�֠��P��%��4��U��5�o�;�c��Vm7"��C����vG"r���ؕ�i�ǰI�KCS(�����2�z�p`��Tb��)�{V-v1�=ߝ��*5�hH��
��r��шF�� ��V�#����-�� "����[ö�Jp*e�4�z����}(�q1{1|�O��������؊$&��֦�!%h��,�-�f��]�܂���f��'N��o��T�!���I���5��h$�Ɩ֐��������K�fa�`�#n�}%�N����@#u�>`o.��tB	;� ��c`�?)SE���T�����>��?�Y�.άs#u	�2�S����l3�y�Fj�8���%�6�@���2�v��r����N�c;b����e:,���� �8X�ќإ�s�����2@Ǘz���A�R�x\���8{�����L���pΩR�r��+i�x�:���\��R��NJ���Z�B�#�%8�cv��Ip���g���Ng���A�n�5�"��2k�B�)
}����k��x��es_�NN4�����<[B��I���;ʖ���w�m��p'NrI�"`e�Z��x���#���2"��Tj�HL΢ä�����q)+��ןN5�Z�l>����Y��-?��F�b���X��T��Y���k�/�c@�	��U.�K��up���v�-?ܩdN�8.w�K��Ǜʭ�J�.�J��֥�Ěk��Q�K�k=TKL3���s�a忥��?���hd1+4�Դ]��=^�����p͹�gw3��7���z("�����@��Ftmog�eau{-��(fUT�Ǫ�F"���>
��&0i�"����Ock�#�d8?��
����Z䗩6Ԩ<>�7��QU?�|�X�M���������h7%I>Ƣ�M�jZx"��yI3����^(IFA�P�ER��,�m����;<h-)-Վ!�<c��f)�(�b�-�r#W�P�5]w�
�ϒ(�a0}�U?^On�=}"�c��Z}�6��>���He��!b@���
�BԽ��u@�2ި� ��>�%�@YI��<���ɌE�)_�z��c$љ�pw�K���9%�7�)(�qtr&�����ý����w6�eֆA�7�V�b��+���	��3������Ի�:�R���>���'��3d�3E���A��s{���n9��d�U@�Q̇���"P ����=�`��q��å���o�N.\M,
A��sێzw�T�/�-��о������=R�G�싅*Mt�)_ +'
h�S��oj>,��>?*���ߖ^��Vi������E���-�%3�9����Ff���@�g�{mq�sTT�k��8���sc CU��HU�8��?%�y��H��C�Di[�������2�'+����lR��
x{MȨ�d���P"���9w���˝� &N�l�!�%�Jd}Y��OZ�c�D��Eq�5*ɪX��Hg;ҿ�N�:J$���(�� T��}r���c`̚�VO�U�z��!�n��_�~x����7���I��wP�}e+��$� T<19����B֊|Z#^����*cl}�â� �5m�G��*��zșs��Uɜ[����.�5:t^?�l��%�ٖ�(��ds:o�E���X-a2d������u������͟z�̃|�{�+#w�4��YB;��}?l�73�Q����t����#�߇�:`䛿<d��3�uo�?�%+��Z�h�7k!+��-��F�"
��-vel�� �����K�v���[]j�j�t_y��AM�'eZ5��D%�m�l{	6.�%+YY(����{���F��Y*Z&���s{����R�*�yr��G;���M�|e�-_�nm��Z[�/�R[6����x�W)�j���ZF�x8����[����^����sT���G�[��7���cS���d#�'��_����W0�sd,`��,7_�`�����=��WOG����޿��%���\���1� �R�Z���n���+��g�D���"!gO5���yhop?6Jp�\��2��Y�r{�>�;f�8ų�;�=˻��R�[
���+U/K�D�a�|�9h�ڌ]6�%\9B�t�,_ܫ.E+�m�9>�Av�u��Js���Y(�-��/��/��w_[����	:d��ead��?�dw߿�w��{e[�uh��~֕S8y���O�l���Î���|4��B}�^��DME��z�R��h�:���k�`pUo4���W_�`2U��I([1*g<_��������9;��g|�X��w�O�*�����;˷�Z���r��@�"�k��,�i�[8����A82Ƞ�j=����b�e�xf��/4��	�`�\��q?�fҖ�8i��������V�f~���UO�G*�ṫ�&؅0�Cy�j;ј�$N�`���&P�����z��Ǎ�e��pAi*�;�ӝX17�!x���Ԟ}��%�ʿ�VLq����:�*�c�Pd�����߿���PG��$��8�WI݇��(E�a��J��̔ʀ%��� �d��CGK3TבsysqˈQ���s�Q��P�C��lu��{p��L_����e{�������t�����o���Sg�jG����0�K.���Q0<ܾ�>xN�u��jҌUU�-��Md�*d�hu�m�*�%����#��վT9@6�C����S;WI������4@ӧ�$�5k%c��,�
,
Q���}?�3-V��\��鱽�.���o尩m�e�A�4<[�D)ds��j'{���Jh���r]Iq���f	���p7�);`p��#�.ol�	,f뱗d9�G�܌U 8lC�2�b����#�����E�Α����?�����T�/�����H�
�I_8I ����Ǳ�ɑ���$�,�&��i��y�0��]�43�(��1d�7��ʝQK�{f0��v�.�s�*g}c�2r=xeP�3gβɝO@�f4	����0����V槏�Ut_I`p���Ǌ���bn���MHP�L�1Dq����wrlm܇��t���LƘ�l�`�߳��'�}����=�B�Y��~+o�lK��d�{�A����  ��\�"�����	�s�+ $����W_[�Oh~���{��#�坭�.�-�7jX���x}��! x��_������vv�_��?�4��P>.`f�����{�����-�+�f��0�y�����6^�6�#(f�� ��o*�q�����ģ"�Ĵ�,e���d ~F:����;��q���X�*m��J1���YǺ�݄;����dO���38��I����͉U�>�$�鐃�&���w��N�VۆXs|m�D�RU2�kVe�
�ڦ�^$I
��!���B�z�*���$��3��v�02��iĲ1{9	[�0Ճ�|��������Е��Gr{��?r�|4N�o��� �s�9���rt84���ci�q��;�nGI�,B���B�u���1�.�5�EAP�v��|i-#J�'-!6t�2ܴ/�F�By�'�2�Hlí�M��h�`t�;�tn�wMNԔ*���o����dg���I�ڱE�evW���M	7P��J��Y�뜆�
�.f�T�Z �`Fߩ;΂�Q�2��{�%	"�]c��SL[�x�)Q-�:hf@4�IT ?���N��bfQP��^�T�|!ęͲ�L��BT��F�����������r	���1���H)����|&}��S�ޭ�G�O,B���o�ʲ��X·	�}�_Ni@IC++]��t�S�jB6���4	��2��ER#��B�28�g`ՈF��kq�r+g���:�9��fɀf��zE�5^�x���}!�B�t��kq�6t��p宆���d="�9���`8f��ܵ�A�zp2)��b:���s�,G7@H�Q�`��"Y� Sns�?Vo��N�����y���=E`q��}�������E�õ�^"��nh)��M�u��~`o�����_���/U����G*/-ΪQ^����j�̕�-�>o9k�\���bA����pM$��g"W��S'����%��yj�- A��SX����i��� ��xX.������d8���3;>>����k5��A�3�.mD�~څ�Kq��4l7�_��l�A8�m���J&��t$�su����6�k���J��!��|.�zfd�����r`��1!Z�
� �56�\�T8�(�4�r{o��PJ:�JH����h�'���z�#��
ENt��R���%�Ψ:8��=���{�������V������K���{�.�ʲ��
��.ܢ���E!�T+�}���ks+bo���Z�#�P`���C�0��D��Ʈl�6��KI&�c�~P+�B�f'ǽ��\E�w|���C�Z6S�CSG���d<�ʻ��·��X�|���:)"T����'rv�����/lw�;�y%e��Tb�"؇���2���=��}��Kf�R��Y ѫ;RS⠳oH�+Ad�t��>i O>���M���n��Y��6�]X�%^���P�$�+u��6��O����ֻ���Y�g�0���y$X"�ONΔA-`�jd:4�ŉ���"/�V>5=�N��~�_9K�׫wG�{\�g
\t�>�c>�W���#�ʅ8Z-}F��Y�e���\�?[��(�D��b��C$m(2�d�G�z��������������X�l����U��C�Χ�Шjtu�hl+8�~�ɏ�YOi4�Y]B<��ԡõ���Z{��	� ��L�?�|����{Ζk�%�Wo�{�H���D��e�jI�K4��ѓgr���~�-�P��d"�Ϟ��I����D�L@Vé�#�hv��O�0H��ƞ]
�jA^|渒����+9�D~����۷o���{�$Ok�%�˳�8�	��B�ӳ'��ٷ��_���!�L�|!�:�w��9��Fc�y[)�(`����\�|���g+�F�pO�N�ɣ��G�v�?_����ێ����
�Q�t�hA�5�O�5��������UαQ:/ �;z?�����	���՜{�X������#3_���k��MhϠ��}�aq01d{QS�wWn�YM�u^��m� ���� ٹ!U2F�z� �K:F��
jpҘ�<�s�-nJ�UdZ	�����h0�,T�s���^��FW�Vqo���4�H�����g��﷫�MYe4��4
F:��bf;� ��W�v,Q�͇�������}����\���4F5۾�!�����dM&-+�O��jL�������A3(���5�a-"/� �٢fs=*M�;�@��ƺ�����������c]��;�q��c<d���q)��>�iz�I��*��؍@��o����2��~�6aF��1��&����t�E��p�|#ws� _ڡ,�4�i��Žf�TU�����G���0+�y�?��l����ļ�����,#c�wm�i�ug��h,!I�:�|#��~��V�i52�����F?���j�@�s��	-D�3��hu��jS�B���f���,���wҌ����\�a��Oͩ��j��2@�$m�� ����>��s C���Q�^?�w�\u��"���r�AP����`���f]��_���Y�.��ǟ^s�kvV3����8�RP^�^}�N����ՠ�a�7���K�]ެ_[�!��'D0�\j�yu'�w��N�7�P	�Ÿ>��G_}!�|-WK�L�K9���x,�:vȫ�:8M�6bL��� ��0o�[�ƅ`�@@����?C��c!*:<���B�\��_���-	��x��6A�����F���Q�7����0*��|�AF)���kI?�����4#%��1ދQ��b�U����SH��K}G��q�/�c`n�ӗl��X�EZg�ZP�� 
:f屯Wj;��{Yk�\h���ӧ2�9Y���!�"�W;7�L��� PN2���,�<L��X�D��n�{{+�3���>*L�F�,�o�-E�}�kt���L�]9���	� $�0@�����2�T��q��U��bp��k�������Y�0H{P)�=�M�mwec��c���%�+��#V�4i���|vw��?u�MC���b���~�^�/g����^�t�����uw����W�������������9�N#��� չs�jlV��=�64+66�?Y��#�[��	Y�c؇����?kﱳG��Ɔx ��C$������4�H�����X���2+�q���6ךEoY�����Ӭ�,X�(�
 ��"�������?z,w��Q��#b@h��l@ߘ���Ò�>U��RD%&�Y8?�7D���祧)My7>�ioX�V��8��xlPUy)ru�jV�b���eN؁]�0�*�#�K��������a�d5(�Ao�D�u�A�Y�}��K�O�Wb�|<��	8e2�1�%���P��:s��c�/`4����N�J��r�qE68��[�Cttv*�5���𧋗��M�_N�ӻKy�%*�s�|�M`L�ݷb{�A	�}0�d�#"��M5#��`�����X�#����K���a�0�}:9?����e���jz'��|C��O���8!�^Oﱫ�=�L�����tt�L�K��_���3�����L�p�@�� �;���W29{!�:@맦�Q������/dy� �����-$������@�#���q��˩�v(0�����2l���Ӿ�Q&�*�E�f0� �[�ca'O���}���?����D��~���7.�������N�dD�c����#>�߿� �~����_�����Gr��먪�5"���!k�z���	p%jxNOO� O�=*�M&�Xl.�,�&��l�	����\1�Q�u������=��=9��Q$7�I����-��2���F㳑L֧x�i���4
#W�p��Cy�6��$T�J����I5;V�����-���+�puͶ�h2��	x�S&M	��ck�`�,�$E�J�cQi�S���� ��&��'D�l��ك�����m�?����r�p�j�[�GP'GIE�S6�e����2�X�O�ӑ�G����j�{��~�j:��F��z�{��l�n׻ɮ_TհX/W׽~z�����>�xXn�����:=b�	}�n��F���Ԑ�S���H������[��ݽ�i]�IT8>��0��������s���J�Il�N8�� ��i�\�~ಔn�YŦ��n�#P����t���MTF2C�O�h0f�(��e�p��ĤX4h4�h6�%Q�=��=�� ��0�� j������˅f�z@j�p��t�j� �A%;�Z�E�ݜ�Q�N�
Wĳ�Ј?h����GH��J�uhi��	�������P �Ӭ�G[/f@�V���Hc-"�#޲.{���06��Ac}}"�9��1K������]Q:c��,��<�Ȉ>�i�aּY"3/ �4����A"�1IX�n�(���G��"�d5�WjXzF��r�؜6��[C��z���*o�1�y�5P"Æ�F�a�p#(��+8Z�!�z�4�z1��N��2 /�h�D~l��i���{\�_:ŎMS���_����g�.���W��C%A�H�]��2�Y�����e
}������M4��?���쭔p>�������JyP��3�'���WW"(�@�2����j�uEC��01kΕ��Jm�|�Gc=�X�b��`\dԇf�:T$=���[_m6[5UD����D���=ܓ�g��-��5�]ۋSZ�#r��b]���"̷[�9�,{���۲ӟڢ��w+y�v X�!�
�+w����ż��s���A�Y�3�:ɻ9ch>gH߲؏5���Y�M��u� >�:V�N�jo
��SY��>��Ŷ���qĥ�xQ1�J9*��}Mv�#�Z���Po4�5�K��Bz�@������Űgi��2���b��"�1@gi�����AD�)��.}�-�[���]��KbX�/��=B�B���a��0HyV�����|����x�>h�N��޼y�T�UU���������|�o6y_Mr��\λ��E�--j�_� {���f6���=U�f`;���e��Ǿ:m�H���^��s�Y;���-e��R�\ڭD!��fI�����h�G��	�08ͱ:�a�ё�̌t���2a��Pd�,��`d�XKeN��y�[ |a��I}u)ѯ-�٭:�~5΀��k��u(�Fa{���z!�I�������U;�g���d��룙}�����%��χ�b�*�U�ʸ������j��wӘ�t�� Y�<8(:t��
�RQɰ�5<�����O¾�{9�hd1��J�I�ZZ�&���G���>�h��L`j����u�{+�^��;R��'C)�L�Q�2�S����^���ͭYKR�����v�֐��	cjc*�������S�v���L3�'�gr��q~w'��Jjw��Ϲ�4h���
�������^�#u���F3�QґS͜�yCƿb� ��|��ݹfK@9cr�K���m$�j��9Nl��:��PEUl=��7����i6y�ו��lQ&����g�����+
��C"���!�?2�{l��`��zOw��Is}�*��~�o�����p����Cg�JE�_�����cRO�= ���dؓ�ѦvX�?a5�� ��j����$`��YG������_�^�w��u��7�����Dz�1$�82��0(�,���ͯ#�
�Oa�k�A���#u1����F��E�&E�.D�Mq�5&)���գ�s]OM��G�YS�G�i�L�2Y����Hwڐ��u����h�Qy���(9�vd�O�(�����e���[�М��?��~NG^�@6u.�4������@jɒ�	���1Ld�[�	`.=,��K ��A�!�uA�Ʈ��O�%�cha-�;�|Q	��oWD�M���;���ȡÉ�f��j�����0����\3���j�������cˌh�J/8P����Q��hgd)���!l����1����4AU����,j�����ʣ[m!X40�5Җ�C	8�I����} �m�*s��g�FG�b�A����@b�9�L��i�R9�@�:b��`�H]m��jx��[���*M�oG�����=-o>���?�F�/2��<+)(K�as�@h-����)��ҌsF���3���0��wΡ�+��D��"�����8
3~���{�޼!�����#��3J���!�ͩWN l����@�e���R�w���>BP�(;uU�0�]7�`IԞ@:���s��W��{l��(g�R��
��6����V?J��:��xYu���p>�rs:��m�-"{�$詌�.K-�,ʝ�J�g`}s�)�]y��T��ꥼ|�L��9>܌��~���F�;�hV�#�pU-%Y�����$���/ʏ�s'�[nHM���x���f�ku�k=wǍ>K�N�Y y�����e�Y)Q��5`��:X�q��1W�����{�&#���x"k�֦|��MO��_��#]G�iGHOZR�/�2l�5 کs]�T�93��ܱ*r�c
.ypϫD5'�e,���u�������g$)�C��������Ͼ���Hר�����?��~�{_���Y�y��3����m^����>�����m9cm4�RT��d�������*�z8��!KE�a׷��WǉYm�90�K�20ރ�Alb�#`v�#�00��P���P���g���l���kkJ��Ȝr���$k�{ôG��z@g�)T�j	�g�Y);�*�?Hٙ��Q���.���%3�" ����Z~���;y��N& z�tG\L�W��h���}$�Q1��Y�g�Ӡ���tr�=��p�^�z�����{�O��O,�K�"��c�B�:%ׂ��*L%C��?�������:���կ�'�D���l��x��Ku���Oҟ"6��2W����|��={� r�ՙ=�=�3�x���z�m�*�)�P���Q`V�dE�5�`��L�P������w�Fa��4aDl�s��U���I�����F`�s�#fp�}��;��hc�()�j�jK4�PA+��|�`t�;��Ԃp�����L�z0�:Hмr�dۅq!/W;]�)��Ś}�xhU�gQ3+�1+N�I8�&�Q��O|4�wڭ+;H�?�(4N������&f��1#�a����`T�����*�ICr]�?����ţ��P�>�Uze%2�2+��=�k���\�Kk�46W��0��k��&2�����iW��.=*	+ X��Y��qm��x�u=:�.��9v�I�0y���)8��}͌!%	�p�O��!X,�|dA�l�����ؖ���Z3��[������4ۉ�˕Y����I3Q��i���t4@���n�Fw}{'s��q S_Q�����J��L;��0�1����~mO�8�����;�-�iFK^����pNS6���E�\�����4�7�
Nc���������m��t2��tx�b=��� !
����n�{�A�?�j��yQ�}w%KMN�����&�-m<�vu?c@�����J��c/W��!ƵL��\�t�U��ύ�
������J�:��C�5Ko76&����ؔ Do���0�����b��)]?��m(U{0��GL��#p�B�67�������m���Ĩ��}�:��C^4l;5z�Ͼ�R�'�tXA�k�섴��Áڲ��ǎ7����vh]��8�^���|]0�A��κ�QA�+�g�i���{��P5��W���`�62�>�gd����&;I��!������O�>����?�/�_���wo;W���Mh�A8��8�pnx��Ñ�Ѩ5�<���;�#Ȕ�^G���X<���C9z�ic�BDyP���lq+�y&��xٸB(��m6^��!�J ��}�����Pd�(�s:5BUt-���'{�5�m���Q��]GkY�����n�>>��z�=��^ܱ~3 �0��i�hDB�]C�yUX9��z+��b�x�5B�ˊB"�E��k��R����!�q"˼#c��r�Gc���Q��2B��a����YZ'J�E��/���z�6���sb �Y������?�&c�+V������UF�̅���,$ge���%R�jM�!f�����>����G�K�brl�G����{�CP��3$w��;�9��}��_��MǢ�$#f����ou?L5��'�2U�H����! �f�	�*!s�PF�5��>�#���h�eC���q��ݠ�Ux
��]o�g����_=�c%~��E{�˳�Z�q0ƹ��#�� ���4k<��hL�T�c�;v12�I�D=XuN���J��5��@b��R6�F�eZK�H[ ,W�N�%Y���@pmT;����G��Q�g���D>������y��\|��<�4l�b4 x�N	���� ��ؠ��>���2����_Au��b&9�e��NX��g lC�����x�5���F�bSC���W&YB��qy]V��:�x���1��]jJ~���HA�p"t�K]�u���R��9�g� 4^�<�Գ�u��U�xq���3�)帪�sV�A����`PC���'Pe�$-T���u�_|�\C�Q���~Ǳ�^��*o�̈������#uL�}h̡#�\՚�k��\�s�r�ȪH=�Z�u�֮G�#ɔ�����o'����v�������O��ͫW�:`B&6�Z+��Ea��Ua�����FF����r?O[c�`Gp���T.?��0�ÌB��w.�P�L����(�13��L	,S8k\�#�=S/���\�" Z �\[9�:x��#d��H�����4��Vf;"��ݞ�~����&gTj����j�٧:d&\ Iyi��Jhj��� &��c�_ץ;$xe2�ȝ�ww�|�Q�D�4�Q ���}�F�ZJ{���{�F$Z�ےP[8�7�3�/�j=g�����h��d_��+�L�0�8�]۞�gU6c|�]sp����ฃ,jQ�m��b.���Ga(dYVb�cy�c�떳�\���ct�o�1H��m����C�ld��)�\p��f� $��Fdz�M4 t	d<x���5�q�@njY�V�Xf�n��������[G��A�������EQzD~�.�����bιlhB�q&^E9@t�KD�r������4�a=l�` � ���eUƱ�o5��g������M>:��[��߿���u�X��!�,w ��J;�:�t��X@�k1�jAQ��tJT;Rb�pv�G�#�h�P6Kf�A� `�~l�y�O0^����c�o���ɛ?�(��;��Q	[m�̨OV��4N��_� y�ⅼ��o�ݏ�����F!#��.gSy� ����B�7���w���Ɔ��$��tg7@�$g~B��ژ���}`�׸r^�>h3�n9z�j��J����Nc"7Xt�aC�~.@m���x��K���h�c�3��ߢʈ�`)s}}�چA�����LL���TXy��pN�,	��n��r��J��������\/�Lj�>:�s߱ЙU����toDww?����d����?�=����p,c�I�/�ZpT8�5��>�)"��Eb�aݒr�p�>�L!����v�������.�cF�݅~2��8X��"��m�
@��w�NLH�Ê�ϳ����`�,�L�|���Z/ū ���
j#M�H�|q���X4�l	��v66|���!��p�f�(���>�ܸH[��
d��B�l�`�K��
� ���t�/����2�����(�C��K8�ѯ�[D�C�Ʈ�� KXɘ�V��枥��3I��ב��j�۠h{_q|i��������c(��;�&��,-k&X�G��IG�����Ɏ�B;��yq��Z/�#B�ZY؊Ĉ-0{�����;�	��=���
L�N��/1�^N\��3�0�>�-I�3!�oM �5؋����TEF���| ��w�������f����1"+���Ѳ����e�;����Էy~d��`����U>J���,)h���r$ 1�[ZK8{Ȅ�8#!�[=[�4�s��o J����G�Iy ��uz+=od��2����9�1f	�5��� �9�S�ޒ� Ë�{+`�`G3�هK�@�������r>�	@@�<PlԢ����
�5��3�i0"
q�Y�V& �'���ͭ��Nz�`%����m�}��f�o������g_�.t�J1]J�-e¨�D&��:���G������I�����M�Z��I�dd��,>9���cQB����*���*�<��
A�6i���%F��3'x7���g�;�Tu 7�x	B�웹4 %�� {�i�#T4;>������)n'��"1*m�� ��1�E��_�p��)�d}w`�k�����W���X�����Y�fԗm��k�3�}�7r{{/?������$��A���
r����oy���|��� Pq����[���3=
VRk��I���ſLEв��sp��v�U���E�PP��z㌆�Q��|��~6�B�;l*�;�W5T�x���D�#���p��>+5�ԇ��Ai�I�U��9��:���~�	1Uo�zt,�9�Z`��j>�[mu�"�D���5]�O����s���!���[{_��8@�@������"SSĬ	�w�d"C��ܘ��5����&�3�YR�E�=�+��t`a�0+��W������m%*�]�����s�����L�����C����C! H��5�3GE�)�g&��}�?����'-�'��+f9udϚ�k�<
���'�'�꘨�3�V����"~��3K�Y�bHR0�p��I62�0�$8�s|
Z�Y�zL<EmҌ��3VR&�0��&N���Ğ�~ 4�+R�6�A���/F���QMXYS`���t���5�i���L�.)BR����y����a���(���5��'ǈr��(��W{P�������$�z������E	g�1ִZ,M-�!2c�	4��?LɐȬ���WþX�e�$��Yf_�!������{v5ji4_c���N>��k�u���9�x��z"���T+��M�^]�=�-|� �ɑ��ܐ� ˁ#ci�c{�6	OT�f˩Lg�ܳ��]C�#��5E��H�m#<	eiSg[��1FE)2:f���>��O����>\�R2�i5vP�uނ�5���x9_���z	�߻[���d+� �sr7�7�!|v��!d�sv:���+F��b5(�%j������h��;�j��M�d^����p�+�ب�vS�:���v&���G�r'&�-��A`G�=0(;���}�ҋc�Gp�!l�P��Q8۶� ���������Sj�D��9�tU��Ũ�88}hu{��,Fd,�?����d<�����U�G��~&��y(6q�Ԉxp���m��QU��VK��Z��CCe!N�����0N���N�hy����т �w�<�B�����m����5�̔��jČIZ.zHH�P�it����zࢼ��C��S����r��c]�uD D5�}�={._�x����ܾͭ/3��;�ϴ�7/��X��a��(\͋dj�և�p|�(���K=����$<�)hBv}�0#�������}���c4.���V��32�ӓc�UØ`�=\]��ԟ�� T�h�J�z�G���rFG �������  *HD�� �囿�%��w @]��bǔ8�t�Wյ~�H&�ϩ6����7����{���2S�b�H�7����K�W�d ����~�,O|�� �����׿�l8$�y����J
�;A��ƪ�1c��kvrqαɓ�Sf�ؿ+ۨ�ޖ��� �p��Ĥ]"0s][�X0�
�Ӭ� �H9��a��5xf"k�@	�^?W��5;~���������<z$70����@(�=��V8V�~��+���-3�_s� Z�q�>,d���>���É �@e'�wZ��"A5@�͑��@�Y!߿z#�����3���蓋�t5��h��Pgry{+K�$ UE����,?\��h"���q���C0m��������D�4��� ������|� y����)�j�<�i�i�jg�) �r=Dw��}��)!.}��5[=�xĳ| ֱ\���,t3h���{�� ������-�J*�YkV�C�d/�f��6�K��bk�w1f=�,8�8N�K9=�V���$�cY%�`c�Q�tU.$B�7�P�m��(q�AC�![��@�v5�b����2���~�1n8_�Y����xUɡ4v��b�'f	�%aA���JzM���#ǈW�}� ^}�9EQ�o�/��k�����Cb���6	�0_��t�
��$��%^���U^����ޡ��ʁ��?�y�6b����JRg�S�6 �ɣz��~g�
$�,IzǺf���017c�Q5�L��Q�PkYn�6/���� �ɸ��ӆa�`
삘�����x�L���gS�l�l��@k�ib�7��J��۽�hX�j=���-I��ʂ#8{�~�\?J��Y5~X[|?����0b@�v50�x�Lz�' ����_?�T۰"�POkf�G����������bÑ?Vj"�ŷ�Þ�>z,/~�3I06��3��n�!�7�G(��yVԉ_<./���5�R�j��_}s�AZ��}�22���f�r��1����L�׷2Ӡa-�+�^�m����_}���/�����2[&���o��v����]dbj ���s٨�{P�W��e�#�@W�� �K'4~X�-Z;(庐�)!F2$�]"�J�jd3�DY���]�̎���+f�5�s,nۘ�5J��1s�J�  �a��$*�nrl�	��K�V�o,�K8���(��c��@�g�&��#xj�����~�K�;<��������X�.!ȭ�5�E��0��i$��\۹,v���́Ve��볘�CY���� �pB#{��^�ǃ����-(�j�v��� H~H��j�������P*�@!����饰J'�%:�韈��#}1�4]5��O����)�D��l��(��bP<���C�k���2���љ�q��v����@a�Z2h���X��4����>	�ab��=��/=H�6�gXRJA�<P|�U°�g��zMF�OIZ�xo���at����!qK����&z���G&1��Q�� ڒ����r3q�őo�)��0�	��}�x�+8�8<Ў�"U6�x�L`�"�l�B����x�5Bfe�L�w�~P�h,Ǽg���[?��ݱ��|L��6(�I�A�m�Ca�35< �ầ �h��ЉM��R���@!�y�d����
[��g�|f�~>��Ww �C��G��37��Ѷ���Q�8�����ϭay�f�B�
� ����^2	��'{ǳ*f�xn��c�"6�-K�Ec�o�ϕ##��ob:ʨ~L��/��jf���쎑�������j�|`h���%�؎��1�#��j�����d?h��k`��َ�ţ� ���6J�����^�k<씂�̶σc�2k�3Ќ���I-]�2ve5Q�3wlA�!��9z1>~�����!� ���Ӹ_�6Bj����\0�6u���������M&���Z�d�Y����Q[0��Lo�� �'G���X]k�����'m�ΤgC�ٹ�U<����:��%{/� ����	�#���� ��4��:vI�s����׬�aOāW��`O������b�@`���6�= ��U���	��$��``��ed��(6ɜy���q�X#��4P<b����&Ԁ�f�k��LS��1Ѡ���wl�+�+2�j%ɔZ��˵7l����a+�������zP�Gr7]H�A�ӟ}+o�w'����#�,�2�OY�L�	{�Y�Pؠe�!��}wd�gv%�-T$0D�~��XQ~ol��ϫ9P��W�o��_�8 ��S<Np[�M`zeuf+����{jg���ơ���f�(A����A�)��^]���0�=	��Ցe��'n�3���Q�fPO4����ê�����Ǐ�]�H��; f��'�^b��x�^G!09p}(K�����$3ؑ�J���2�V��y�\�z�kn�߷��X|���k�F/on5�|`�V�4�����U����|���?9�vp((o��_�j�GHD����\���1rd7�g�����p����em�c� ��W�� '͠�[��}]X�I,�x�t��ԯԨ��[�h�"h�q!��D_N��˛k:����,��	��sJ@�=�v��|�e��&�YI��c@�2�U���t���1����(���N�l[��NAu[[�b%��d��*
"�)`D2��[P�-5��u*�ŋM��S2�7{i����{�^Ik|����9��5=(v�kq�_�1`H����"u>ż��'fO�mO�=V��4 >����kӀ��~��m9{%�a���(���� ��te����s}��j��T)��P���˜8�S��h���A1O���Ńbx|��~U������a���6FNu���!�z���u1i"Q�F�� 5r$?��wx��FS����?���0�V*����.�cN���쌚���R� F���i�?sw}%W77�X.
�-�(�!Ȅ��P�F%>%��kEMl�C�1�gEm� �YM@��5 05�z����4o�d����/e�yq=WÓ3u�Oɳ�$��O�:�f�$ߙ/�	l'���U�;�i�je���C��Z���ى��Ipl��dc������l?�ן��=2i�^����!em�#��#L�37sx�m��t��8�oа��ġu�]U,-��s�fµ���}��+ ��~0����{�I I�b�@gqh+4F��L�:�{�F�a��0`0�8��가m�}�4�g:��������Ҁ�Yz����zԕŸ �	�}�_b��m��3ݓA_�j��h�4kV%\�������]9�)���^�2�����c�܀�5q�@85;.h�#�
`K��c4-1Q��ϙ�V�w�s�e��MV��"K-#�A�M˞�ҽ�'D�3�WÀFĆ"��\�WhAQ�\������U&Gj�{����F��ԛ����Ȣ�h�	@0���td��@6	���1�+k���Aģ�Nd03#]4��&zÒ#H5�R�pv�h0������V��<�1��+/�+�`FV�`A5�슪�°����\Ѫi�����.7�*��e��@:
<��c#�M���\���ￗ\����H��@�3 ƅh�]!��wD��j���w��� x�ږ����0�I��Ѿb���?`uh�]�u���*f��b���Qb*d�����A���nC ��s�[���*̑�x�a|"�-�<;��%�}ldX�8��QI(�Q�> =Sc���*m�MJ`$5=8{xO6�`SA���}!���D)�6���&�x ���F�e���Ta$a���T�ț���22���]�{�V�э*Q�!HXM������pШkg���A�����'���T�?еm-dtQ��6[NX=�T��G���{�=���~�`��bA!+�9;=�Lmb��*R�@�yh�œU1�a��O`��/a���D�8�A���G��<�?n��C��c�/Y�0���%e�;i��S����C��a���4K�b$�%&����3�ӄ�h�P�G�7�x��d�9��@��0W�R����wb_��ź���*�Y��LY���`��)��	��@ک q�z��fgrt<$ك3���V6�7�������Q��T�R���i��n����p]u��-�'�xK�[�����>|�ƋLa���|�Dt����'�����S�� =^i&U��-3�(���</~�W^Y���AA������~����j�hd�N]��z'����*+�0���v܉	����:����*�_���>9>�L�x�����m[thW ���}b�+&$y_"�׷�-M.?�P�
�}���,1�.�DFCyV�<֢���ןw�V8�B����u��>=����``fX���OK�[B;��r2"��| D�q/d{2�3�`#�@���{�ә,0K���trD�u[c��_�<# *'�����ep�8c�c�d;�an�]�\E �� ��Q��{n:  ՞IDAT�M� �^��� �Em\�%@��L�٘�*�D8���N�S[����A���,z&�t��b�{�*���%X,�d_[�3!K����p:bs� k�Ӝ.�l +���z���G ��@8�,Lo5N樠(���@d�HP�@���\�^�Yԡ�ry������t)������L�S��Wz�G���?��5m&�QF�����'#��!xWy���O�as��3���-�����r!)q�$�>׾OqL��W��������p�W7�Dc�;0c�7�-�D�R�V�E��,��/�͇�.yʝ���6No9��z�yE���~yh*,�?�Itq`a��7�d]#��	O��Gg�E�f�R�� �T���Ffb�u��^b���D:D�W\U�c�`�g6ӝ�Ȥ�����e _<%�{�����5N�bF�2 �ᧁ��=Y� "sAf���nY�J,^z���x���f����$�N�H�	��I㽁�Gf���M	���v4;�DY�4�)i�g�w�0�=��j7�u�[_�3V�c8��t�	9Av���Գx��8�����%\?�g5���Jf�Z��F����.�V�F�v
c�`fj������0F���ʂu��C+�%�f�����:����������-����kC���hW2�1�F�%��+;�>p��3x�1څ�14��S�$��>��j#�Ac*+�|E����g#������0�ɇ3����H�=�F�a-���H�M�R��ncIʾ Y���y" ��x[e!�n�o�l936�*���
�����|a-��6��A/�h\�o��_٪�O
1��2�T%�es�*��F(1��VP*�U�C�b�G5�n#���r�/HN���Zcj�������-y�Ȫ\n�FaO��i[�����s�Y��������aa�0�:R^�:�D��q�r��޲
9��XY���O�|�'��ظ�x�IX��F��|+��Ki�;⦺qT���|���_���#��z�Aܖ#�X�N~�H�rb-�)���V%Ǔq^�6B` ��x���z�h��� ���x8������=Ia����l�^�q��������A6��2�n��*ū�!
�|�- =�M�}��%��`ú���H����K�,Zu���(¿�DX>v�;|/�{v2Lp����id����&J����Q�\��<v�p�O����|)��yd�B���SY��T��N�Xf_�v{���F�C�`D8��zق�p��z%S5�R�s�/հA�R������~���u��%�O6�[���eH�gg���Riϝtp�0��O��{�� ���sC���
m�&p�Q����O�X���W�(�PpHQ�)3NFG1�����X�#�^�hѥ_����hM7��eX�.�
�9�4 ��t�[Y�����7̪P�V=�������'�2"AJ�]>q��p��I����z#�Wd�Xx ,��%[abݥ�}�r��lW�\���[?fh���{�rZ�46�̽�x6b#z(��k�q����b3�tXM�w�M�2ؙ!?<[�Л��Fڬ�t���!���yX[�jm�c�B�\�x��b�ūz�)��(#ӻ�D0��As�g�����*������y�ςF9.;�	ӷg��20��0JV�s�m����+���E��G�E m#���ARb�O
 {���q��M�y��n�&�
���&#��5=/������G Z�i��L��Nd���X�Ы�F��@��>=f	`_TK㋳��I+�n��j�����Ñ������T�G�z6�k�>�|�|%�plv�.������n�O�"絘C�<(��z[�BҶi ��s��k�}�cK�l\)ž������j_���^A�}�mw��X4���G�>�t��F��#I�^u�(ţ�RlS��|��$*�߰a�<�0����z�� �3��^xp�< d���$����~$�	N��c�h�ē'�Cb��KD�eD�b<���7�9�",���u8O\,ӌ�8 �]Ԥ;�<¤�A�mD��OjA[u��M��#�eĞ~�HZ C���G9����mu ôC��H��>�&;4��I��$~�K��ř��Pِ2š�a$���B��K���b ���3l�K�:op�w�:��n�2���!�c�{��1-A����w@���\�s����Y�O��}`��RtHw��p����s�E
���g]���0�ѵ�yd!Av1p46�jZ]dI�UkEi?����a��=5J���b��Rֱ�$�[t���0��� ���� �r��Fxa���X�tF��EC�rV5��1X(��ZԕZx�P�f8IHx�}8k<�1��u��@�{[���浵<�~�H����p$Լ�e��	�S�y�̾�Qg	�B�ٞ�X	��#��p܋g��0��b�i�QLW�lb�αg����{eĩϹ��0r���7[ѯ&�y3��&�vݜ�OYƌa�xg[��$�E$�=Q����ȒR��c�^��Ɠ�RZ�=n}LS[�B���&P��^���Z/U<O� `��n��"�0x+��6I�,�����0� qbU>��q�����-Ȉ)�B&�dȥ͔��f�Y�P��,ذ�WI�̕@�c,kY���o�Y�;TFc*l�l%]�t��
���/l�|��m0�Z[����h�b	X��Q&=��!BG�?a�$�ƅ��אţ%�)�D�+�\�v��Z�C60MŇ(��1�X�,�:g�#���������Ύ<�ݎ��PΆ���섌}&�Ӊ�x�b�����LB����x�m��ǧZF�&���P Uȴ �B�A-���pؑ-����c��AS��l�V+�G{�>�UZ6�fSX��U}��R�9����]5�	(����-G��tК�6�Z�[V�FZ�0���	q���SN�g���2;�@�7����p�c!Y����qX�\.^�N,���-�t}����
�$�x� AA��E��o�.�]��hdr~J0�C1��j� �a�
�#�U�+�Q|��.�*����\/d7ѳ�=4��y��MX�Cj/ӣ���Ḱ~a��YT���O��b6��a��؀Pb��6(��8tqz&��Y,6��I��\� д�
�`ȹ�"��r��Ā�/D�^D>�Y�5�` K��@�h���~Y��N���1j��P���F �뚹Ќ� �i�lo����N6yjk�m�l�*�#<�p�r��X�iXM$�Y�$$UV�b���F������sñ1�$���s����X�Ž���+���c�g}� n�ʳ��x�dm�b�Ҿ�a����;o��v�#�j��$jm��Y�A�b�沠�@��I��F9[6�r�3Єj���R�P���о�%M;�����m$S5���!x`?ފ�[YK�{���TGl}H�V-`��`o�ք�Ǐ���gbL�z�'��^��o�Y�=�H���ݝ�|�H�8�*���>!�شE�i�E1�j��ȗ��IQ��Qrotr
����"g�kX~�ؓ;�}l�ކC���ɄҘ�M���K�e�(�D0��:G�%Ϣ4�����1�����!�|��С3X��D4�	r�S3Z)��Ч�����~b��� ���цT<>_��;*��c��=�1�<Yoĵ����AГ��A��h� 2�\И�����S�N�N�)M e.3*yq�_��h�掴�K�/1sg���ɷ�a ���!�Y�^����҈�3�3G��q	TVK�$m���!};	g���u�������5gw1�V˒N��R3] ��#�:���΀8k���r�_c�F��2$>��:۝:�8���;0�yQp�������t-z��)̰e��K�0���.� ���}�P	��[I0�תfO��*���vC��V�=u�	P^$!Md�ym����o�0�7iK=(S,F���g��r8Jx?e@P�Bclz�c�V]7E�3%J-���i�g�����&�Pp���E���8�8Wb��k�q����ٳtܡ�M*��@L��`�h�b�sk0�0N�vܡ���o�jm�<�m�<�W1E�6��>�,Y�"/�:��C�V���`¦ogd$��@#��]�W�
j}��^�L�8ro5"���58��s��@����T����L�샓pg�� ���a-d�	mB�ZF�V�*��A,M��~�_�} �|�D%��\��`2��~��dGG2S�q;}�sTȑ�?l�1���rb�38=(z�?�{����n�~`�Y��۳ec��Da�w���_I=�p������
��@kϪY~JUO���(W�;���H�����;����_�1�ǘĀ"�%������x��Pf���avn���4���{@V�N>�ƁZ� k�V��� ���쮙#+�DD�3��H�5�	�k���Q%"��}�}:Яƴ��!�B�5��zF�]8TP�J�r)���<9��%Rd'ڋ�0^u@�xc�1��er�}BAi�g����[+�C5쉹kȣ��Z����|a��7�@����3�#7��e�29�⥜=B�!�R�k{Vb��QO20b5J2Co�9G&�ѡ$n�(��*]#ȝf$W񊋫H I�{�Q�� �?[U{�Ri�]p��Ʉ���:�2��ꎆ�tN��]"��>�0>:�|����	�M `NY׬rp%+�q�� �z���w����u1��:'y&b��`��������J�ѠL�>}�����S9��)���_����N֘��aI�A�M&O+r`�������
��:�@����;���H=ɥ_Y��� �__�d���0h�cs�BA���H<�tB*r��)�ʝy����۬HZ���ӽ@M��Lj��t����4�@�\P0����K�įTq[�l��AN�
X
T�"#�ʺ)Y��P�d������Q9�f��4V��?�Y�5u����M��s%F>�=n*!uw� �u�SB{���f��f��X�RH1��ci��k�Nwķ��ҡ��^#�{T�u>��d�{��<�G�:B��
kSy0a���jMLE�l?�Czs���f�N\Ўm���t|�='Kĳ�%�̒�^"���L|�58P�\U��P � V�+G���$����1	?ЏfY�^��%���y?(�8�aPA��#�)�Χns��+�vYFB�v�� ��\bs`���T�(u��'"/�Ǎ�0D9�yb�2'���N@��.iĨ�,12���eۘ[�
e��jy����)��$���_�6o�������y��C�T��^�`V�ֻ��{�)G{�`<v�B�U����I��XF�.���g��K��X֭c	�bU�X5/r#ul{�wMK���\��^�r��S:�3�n�d�aڬ��P�� ���{m<����Zh�@
��ua��tj���L'<���DNP��d9B�Y�H]�XzB�k_2A#L| �X�z+���H�'GO.��7�h�4!�Q�<��7�@�{�i�0s��RX�'�!�ޱ#�br�HKPd�F6� �#�F�f��,t��y�F �B5�|Hy�-d *>.��^���Y('viLG���y����Ӵgb�����C�K.���v\l��{�,�^�J�ʗ�x��D��i�vT�	- ���^%��bo��#lޠ��u�m����b
���Px�{�̰�9�*u��B�J8�(8�c��"J��-�K�HlR��M5�_���qL�D^��7u�O��`�<轧bmL��<{�{=�X0���H�	�F(��ސf7q�:H�h3ӌ��"���p����c}���d�=q��|v�?ۡ'��\���>�����p7�F�� �d9��Q�,~�jN��tv+���T��w���=�������s!;F�t�ý�M ��ki{��;�2�3H���Lz�HYb��7q��p���{��>D��iH&� �
0ՁE	}��sϱ�p��+��I[	�(��:Fa��cnj�!�� ���B`�z_FrS{Y��_"aQI�-��d���=7���&�10İ'LW��a�T7f��Eޮ9�ȓ�����S)=VPi�hF� ����R�r�}�$�H�S!�2��m�a�Z.���^��_I3_K�ضe�$(����9z�w$8I�; 	� h�^2�������vo߼���V5��Q��F�Z�i��h|?����z��w`LҦjX��%quO,��|�2���n���N��^��I3��z>�T�.��N['qp�dh�hF��,�srl����Kȱͻ3`���Ϝ}ت��%n�~$x.<�ֿoj��mԌ}O}v��F��/��Kb}s�DO�kle��Zۯt��)�:1EQ�.�$2������q��N8�g����ieϳQ{��
e�y���]�5��� ��_[ Y��L�K��݃�p�w~h� �ϑ�g�F��f�bGi�>�׺P.ӿ��X�-*e���Bֺg��9C�M�O���K��IC��g�q����'�6]�X׼��p]�͐�]/.�zYU"ؼ����ۺL�*N�����8���Yi���e��G'�g���A���D�(�F��{�=r	�$�W��7Lu�ԯQT��៟:���_̮3�pBF�f������ P
�K��+x�b+�����?�����~�s��m�C�LĤ��,��=�h�>z��7�o1�
.e`F>�O�ߵ�c��r��~䫽?���ޱ���ƒ��X��֣�	��|*?���b�]��OFbB�Mnb��Ԫ�~��>}L�rcظv2��y�Í� ���N���Ϝ3��)�=���"��3{�����J�� ��#��d���_�Wr���Ě_�r��S]�A]	@;pO��N[.�?g@����2��<��O���Ac�q�Y������U:�ZS��#;	 ���ؽ0��bF|���^��MAh��g�|a�1��+��W�l]��:{��JAI�J�>0�M��$Ym$��õǦ��W#**�
4�n5���A�ԙ���lu%A�{M=i�9���4`ֺ6ck�;Ӗ�L�������-��f{�{�V@��}f��9	��LKA"�Ɛh�i�Ɉz�`��Z�J�9�g�7b&�Z-h�T�U_��28�lN�����-�#1��D���n�� H'��8��q&D~D��� X���`�Ho�J$�b�PlH�j_�3,{U�3��C��M��D�%�%ݛй�D���4	8J��j���l}��@ݣ�J��s|c�]�2P���A��	;`+���r���<�W�g#��wk�/��A���#m��b#^�oa����[J�.� ��h��s�E�w+���ɷ�ge��}~wK����D.>e�˸��E�㖆���1��E�Rv\����˦!�ʧ�v�\>v���ǚ�{�U��a���*1
Qa�,�� "/*CQ�߯��-��'{(��{��!���������� A�������������ؼ6�)�{�T0���o*M������Mm�l:KFp��9n:������++�������=c��8����:P	3N,2�?��яN��dkY�s:KN,`�Zq���G�tBM�>�0
`1�#x����f|��ˑ,��+~զ�v��%(;��O�y����i9��hl�u�Ҳ�-�%K�玸N���\���[�B����X���;���V����s���>� f������&da������Վ*[�eKd��,�ً���ۯ9;_j�}���!�)��� �~ė�����N�ŋ�H>|��j`�2|�i='�8����\�rN�/�Ӊ^�y'*�o/يaG8��2�i�����T������={"�_�����͖�#ЂU,�����P�r�,�$ ���NG3?�(�b���P8ۙ>�.��'�aa]�;����_~E?�/)��Qؗ_})Gz�x���'�z�Z�]�c�[�}!n�����#y�?��g���\�~+?��;�_^�d�vN��r-�J�����'���<��%i@/߾�7�}/7���u�H2���b/�찱���gd���j �i�o���+�Y����m�0��:��=�C$0kqq��E��^-l�D�޷������R���@�
�$6Q����\wL�t4X.A!�g�X���\q5��z2�Ĺ���u�����#څ�o^���Odz{%W����������m���π}ᄎ�B���G��^�t_b*��ƀt�S���p�~�x��ګ%Ǫ���SS5	&I��h��#����Z�_˝��u��б�yd	����T��1��-_۸S�d(�$-e;7^zO����p"-�4����T�x��N�S�^�9CS~����284�����Nݲ��"�j��#�����`��uC��-_��5¹QC��ڵ	؄ \�b�X���E\XO����0��٧�u���A`��Ֆ�8��c3($�U�ao�Q{�R>2��cb$!������=kl��˛u����8n���%蜗Nr�
�D�����Z[:�N�����p��;�k�N�9Ƅ2��eO��L��rT���2�(�&H��~9p�NpL�ٹ����)@~t�Fd�� ��� �
'w?}��Օd#����Zd�޲4FAN�1���� {p^��`�=ϡm�!̸.//E>+	�{��h���b5�h�t��ǯ_�����.�~o�س��NT�Б'B�o�]ɳ~�����X��Xf�9�eia�lN,:pFL�#F��O=�m��7V�%�p��#�h D� �ހ��y�N�<W������u.;u�k]�<�̤@)yL#kl��܁tf�{ԓx��o�d�Uj6��F���[�L�FW߿���ecR�2�a�9�� ʃ����_� @�xV�:T����y���}���ehḱ3G9X�2�hg����jG��� ��� S�*x1{��~I����J��-�#����s8�[��H�4I����W�5�E_r�+�1�V�����^���HGG�)����]Y���#)�@���{U��w(�W�9��F�]g����<L"Նq���I2U�^j�2:7A����|	�ޟ��W%�f�����ܣ2d�����T��=���Cɛ�;�?�60&�k��*�P�⽢�&������o����!�8���x~����@H�q_�>�:�PUV-y���g�?k������>_�FW|�"G�6�Ȃ�U��^$��Ļ���j�ڥ#3R�07��b�#�hPMd8�q�VV2��"r�aP]rFZ�=�9�;%�=���z*N%lW0��lƗc���5��E�M(����
2��j#�fl�bC�	�`Dm���8J���[Pז�8�C�Q%."��F3�7��eK(��F���� l���^F�Ї+�qt0榟��bw���$.	��r%�P�\�u�I��L�2�k��q/e������`����w�ZU]V@�����xzѸ0b�f����Й�-���ڈ��w��w ��Ɉ�H�m����	lx�œ���0���$X���NcdrvN����F�25����hkD�����F�K�?�|�،�Ya!� �<7�� ��л�i\;�=Z	1�>�/����Z�1&
���V��~AC�i �ڤA�¬6�+<�6����"��C����]˶@d����7�A$��*��Bqe*�}��H#�Q��q1M����ée��	���k�Y�Pq�m1�Z��hK�Ԟ����o�E��шz�x&�:����|��X�&r-T]���_���:��c��� �IK8 �~�S8��������_Юu�k�����&Lp	)f�v	4 A���QOiem�/fs2[�4�0B����ƼB����mc(��yŎ����D�D3\p/��n���p������aO=��t���f|��C% |�a_?������PA&�u�/f�֓�(�1�����B�/\à�d%hdf(W�KnB̫��Ll�ļr,�j�⦺�3
$�HN[�
EX�h?�ǠU�Fso5��Q��t[MN���� ,l|!"5+��}𗶨a:i�Nᬒ֐����׆�%����1���x!ﯯ��d3Б�|��BFj4������������t��plM߿�(>b`��s⺾���^�i����_��5��mL���l�����͔>nVi���g>�@0@ ÑcR~�.�����}��ڢ�IG:0}Hw��k�ƘNN��UD���9�jԠ���Y�#�tהV�jF�����[�s�篡¥��*�N�_�V����,�B�	�Gd�(��Ȣ�α7<7|wW�k�+H�l�u�?y,G�%B��;�K̀���slw[b@&�!�8w_\�c��k����cL��0�������,����K=�\J�9,i��cd� �r���;��*�y6T�`|jH��%Q�a�"���J��H5d� h�48�h�3�|��r���� �Ղ�Z�m�<d��K�_䊎�@�#� W��[V�0Ǟ� �7Ki��B�������)F��΋��w���e�{�1�����&�w��@b���U}']{���MXU�n��*�X����9�����p����l�	4�!�L1��󍷌�)��`*T<M��|~[bA�X6�HlPɯ8�?�x�s|��2Ic���EuÀ@E
�a0އ�O�BfJ�+ �<A��(�b��=̜�����������y[:��s��A��1�����4�o���� "���G��R�j��`풦Ey���ͩn�v�3�>�N�Hd��+S5��Ǘp�\bABe�@/ف[�jK��E��#�Ք#ML!���.�&5� ��*��n��A����f5������Q�\Y=h�O�`j�Q�Cv�����з۩:��e�;��l$�"��$j��-4���l��`��|��;��w�Yf���t�n���u]�l|D�up:��k�4����N�����Śe�Bq�r�:F�V���jV��3��Z���y�*t�����B�<7��e��XF��Pg9��eW(���5�ƞBf�ڇ�*�Ի�h���˺��ܹ��PHh4��q?_�c��\����[ �0l�,չ�t�kt� F;j�#S�|�:�"T�����'G'��k�i�?��d�늠
`� :�x��D0) �M�ZQ�-huS:-�"CL�i��"���Gh�Y�� �p �졅@�y�!�ވ��EwX�fy���+b��y�����yY;MmP�{W���`�'o�C���HZ�#!	@[⣚gޘ�OJ2�,a��Cn�0��cV8���O�˚ct�'���zv�k)����@0jm���`���~����MzdI�+�kf>��1G���ER$
Dj	�F-� i���?@
� ��'���� ����Ԣ���̬��/F����tϹ����ef�U)QNF�Ȉp7��>���X*�Zp&4]uT���P�i�#pB��}�����T|�r��Os��c��=v�ר���M����y�/=f�^���ݍ>�cc����h�Xe#����{$&$�qN4P�Q�w��+��K���>�i���O��;�8��g�l��xh��Ԩ�����;���<��mNRu�� 'D����[��%,��������}�U��:����5z'�X��s��2��r�I����h���M�C��)���RFަ_.��ō÷�A#�0J��θY�>He(�!�_-� �\�0��$;ז��ʉB��Zc�dM�5+u����8�1fD9l�i��U� ܀�p���<C��6'�29��8Ñ����X�\;=x8 �P&����!��C�����@Ύ�w|}��T���C��jkо��x"��L��9ս��Y�p8���{��2�h�:�������on���r��4���������^�P.e�5�a$���9��r���:�Aw ˛i��ɪՑ�~ލ:�\1'���e��>>x�T�sBg�*�/��R�x�Z�����l���:-�F�&���a�k���/d���׫��P�z��c���%[*ս�<�x��~��G�j����FƟ}&�� �����72o�4hړ�JU?�@ƼV�- ����I�d�K��Nn{�f��@"P���hHp�o��I�굄�9��R���#����P�El=�����=2Y������]�k��W~M���N=uFŠ� +��:�.���P9��?���@Yo�� {j�{+�{!.&�8�HcB���d�`�o��#����%K2�o�^y�����[v�g��c�v����ܞ��W'~Y/aˤCp��1���`��1�ў��~B�����ޯ�>�:�D�@�
���c|�V�U�-���8��{��{�����J�0��a����w�x��<�ǟ~*�r�՟�7��P%B�m�=nɼL�)@�h[1��iݣ�4�d_�׽���>;`��^�J�#CLYe���Q�	q
���	�&hѸ6�2n��Ѧ��H=�^��"M�zMM]�<�ݠ-?�^;Ђ�<��Av�v3�nǦ�ʹ���-y����ݲ�w��;�.����R��6�F ���2r��3 ��T�l	F,*+7#�Y�=s��\��'+	6d&���?�S�e�Υ��[�qx�ɉ��\+i�cw}����Ї�6����",5Z��B�P���9��=PYo3��~~}��{2!�E����`���ŚC���8>��@��􁆃��Bw��v3�ʵ!��Ut0�2RG�S8��f�kȓ�J�!d(z��,��焬q�K����f�Cub��f��LR#�A�>!��ٺ�2fa�[�4=*SPh� k�����^�|��]��1���ZFj,9���k��{*�� ��
��}���f���$�ܪ�B% W2r��T�\V�P�z]�����~��d�;3�%2H�O8F	`+��1��Éܷ�,�wF��R��\�JS�B� ��;�5D{'� eltjt�-p������Z�,>�.�͡����Y�uj�%d|hgp�c�!�0늜��!����vD�ٔ��SG����C�fL��^����cPQ���)�ϲ-V�f�BXI�����>���^ysے[uD`EK@�\�K�5��[�c�Ї�������$�AL�M}�e���v�q�U@o���q�0�j�z���n���FF���R������?]d�>�u`�c���%~��Ul)`�s��I���z.s�ENuo�5��9^A$542%R�nY*}�/��7�gz��y����ʃ�lx� V���W���p?�s̴�ǅ"pf_�����99���ڡ��g ԯ{�ԁ)�A�*�s�I
}N�L����wlj����	�	��1*/ԐXؤ�	�Fۓ����#z�z� ����[�fe��h3I��@�8h��,�>�>�9�������;PJ� ,�8����׿�u�%���r�z�����koX���-@ؖ�����a	����<+��&[e�!c��'�a\�2�cA�P0Y�q��t�ԩ�=.U�T�gr� ի���+��c��̾N$����de�oF�RC3gHɻC��xڳ���A���82�� P�kB%����i'Nw�Ue  B�u�/�?f$��ȟϲ~]if�/�h���u/dQ�����t&��sݟp�w�>��[�o���Ϲh��{E5(��z����$�J��R��!�'_��f�Aā�IdB=٢���^���Woh`J��|p�*z��t`�V��1f�u0�u��2��Jz���=�W����"[A_x�γ{�F.q^�,�ta�����u�(����b�����^�[w���V�����$�!A^��8_Tu�+J�wf�B!׍����9m������Ku*���3��є�}S]��0F��q��
}n��#ݻ��$
j9��[�mkPqu{%��>[G�AO�s��N,T�A^6�]=ִە����r($E�p|��:�Z�&�R�1����one���b�]�%tw��P��D�tQY��ZΖ�J"��~��Y��d�=�燪��Νl�I�q���ǰBf33�= �a�@���G8w��;��r%y��l���m�jͩ�m�p�č�����������Ak��4m}b���0�#z�h�=u�q�H"�������e��5���8;��f�C�ϟ����y#��!ʍ��8�D�M��g��$��l���VG��Z*|>:���粷ߔ�J��2M�|�8�8��@2ٸ�1Ӧ��0ژhKx����:p����q����wcl-s�Gsø�����R�kS��A�oF�غ0���m�gy��?�)����]�]����,~�\�{���A�[���-�o��2��@,6<�����	j�;S�~-�?��ր�Dt��"LɎ�L�$��U�.Pa�9f�d��4rp���%�"FO�(	z�
Wb�5�ޮX0�2V�D%B�t%,�G��%���i0:)3+�!���N5+q�\���C�3�����ǏcC�j�G60<�$�Ȑ�����}�{u#����'+C��T]��5��SQF��lv#�>{d~�qfS���#�U1����J6�XW#vBC�# �=i���t籁�2 v�{@tBx�X$r���!��j$��z,5��V�k�k�ǀ����Bb7{��0�VӉ5����|~j@�A��D��j02�����U����D�ƈ�z,�8y�ND�c4b��)���"����"��x�q3j��@����f�A7��M�*K���FV�D������*/�V���P9@�$�����P��D���@B��x�A�f�S=w�̃q(}���11U�@"̐��>���I1'bɫ�h��1�8��c*��l2������猦��9nrSt<��[�@��CWu#�l���5 �(�Yj�`���y��G��~�9���!�S��6+�*��@��ƀ�,��-�� ��޻H8&#RPO�z|G�y<K�S����W�l�7�!S�qb�C�F��>���OX����J��mysߒEj�.�����uB-0�m��g�&�����B�$�ր4��NW&z�_5�K͋G�fn��?�"�,i�=U���᳍�� C��	�=�z��h�����C׬2��4��!y
�MϤd�1@����	`+dW±��F�l>�6u�HS��;.hR�l��������2�w#�w�x��';Y�n6�e@)�Λ����[�f�1�53���9��; c�y����+�ҧC�l#N�k:Kb��I?R��07_l��bB6�F���p��M�,U�Ԅ�aL1ۼ�]�,2yRN������q�#0 ^D��R:AS�7�q<�!��M��'�bT.J���g�9�U'��	KfȀ|�!��=yoMe(��!�0G9[�v�=Ae
*K �z���K�e[[]{Ȧ���O�0#4��hƥY�:h�sJ�S��\9f�'�ͮC��/�f�a�bF��Pi	Ң���{�}̙a5@��C��Lq�6�N���֠���:�B�J�K�-�Y��h�`�	�)�mS81��b�l�,��,�{���٦e [�3�J���]ץV�r�D�YL(�1��h@qlpAb���Y:�"�M9 ��>��+`��zźV�(:�	��	�9 �]J%1s�-�)�-Xb_�~B �)�Fc�՚Mr\��E#��:� �S+���tA�fR��z�p�qֈV� �Ѭ�<��z��;Xu�P��'E�7��w�R3�4sE??6�L��RG�B�'lHjj�Xo���L3�Y�3b,7ޚ���d��r�x��
y�2����T��i@�X3�>J�iH�^�*P�^�~j��26*��W3�T�:�g�A�)\/�2����1�HbA�U
CgK��F�=��	�؈�^��Ӈ�=:�y�(/_�����:E�ܖ+�[Pu�m��	�^���l��XiLm�����1f�f���;�kк���T��z���,ù�
��d�&N&��" ��N`H~R��k�6薽n:��/�p�	�'��͹ܣ(�hvc��E�qjQ��_�����5�ہ~��S�zg�v�\���7ߒ�z'���l�g�׻�ݿv�蛟�!?v����3��og�'��2���lJ�
�-h2�/�x�92I9$k���m(~�x<c4Ae�� ����SlN�e��1B�ODo�
��zF��mj�՜�0� ���Ōt:�$��Ɗ���:y�4b���:a�c]���l���I">�w�c7����܃��g��ʛ+u�Ճ�����W�A�
��M�%�UF[#Ҡ�H�: �����Q�½��2��l�l�pg�� á̈�)f���4:�jMJz�% Rb�+��2~�l���i���,dY�0Ymҿ�=�Y"/p�@+���k�2!�zrE�ΰ��cOf���gcA�{�2�FǛzc�����_v�B'�"&��;=^I�)44$�ɑ�d���A{��ʿȌ@3�q/���> ������j��=J��Y9f=��
d�xVc6V8��li.V����\Q3fV�V�Q���QrBDͦ�.�̀�/Ju:�S�:b�.*�9��g,��=�IQ����N*���Ý��: ��\�v)���]g����"��P�V��|.C�B,b��ݯ��mT��=�7Z���um(�X�hޥ����ǹ����LkB6��9Q�� � ����v�L+G
��ʣ�,2�Ț���'N=�Y��Q�6���ǙM�J�h���K��T�����1I� �D��/�Ֆ�tE|p\����4&Kǃ�W!�d|��@%1'o�7D�m>�l�B��L"]u�����E���4�Qٌxm	m5�=`�h����9�3b-�1�s�P~���¡�qƕl7cZ�4&��^�~�g��'�˥9�,N\�<`��g5��}g�=���*�{��w{曒�{�f�Zl���|WJ��B�c��4 8�>�sD�PW���t� �bv�5�3j��q�cǢ�1��yN��&��$6c�ގ���	�Q�;��0qjt�K�aM��zf<���k�_�g�_�9�\b?O���hR^
��SՈ�h��rH{
w�^�ԃgl��[���r�qh�5��&*�XHd��j�?<�\�Fl@��7x�{�.Ȉ�����sñ�Vf|Q�EY��?d���f�4�Ȋ��FD�l[�a�� 87�,�4`�j�f�Q�D %��o ��IL�[�'x)U7����=<d� �x��Ǭ�Y��)�2�9�8(Vfd��u-8�4$=�b�24xLr���`�Ŀڊ�l�L�(�^3������߃G�\���X��h`�ׯN�Adq~�[�jt��e�+�;�1�- �ح��&D^���)�2ܫ���E�.RK���`�%�jHd��]����q"3]�Dh��糦�YP�U�O0Z+�LƲ��:hP��-J�:�fh��Ѣ�6&
. d�`D��{�ZN�F�b�I��Vs�s�.7@���%�j�ɏ@�n��ha))�AG~���$|!6�h��=>�;Р��$��	�Ԥ�Y����ܧ'b�mͲ؀:FR���������ݧ(}[�$��9u��Ʀ���rxr�YzY�c�����$@XG�mİBۅN7��O͂gT��#�N�1�`S,0���3c�ԟ/�5�����>r��8/ֿ�<�V����D�'	���衇k���N
3p%8:�p�!s����]���+�ˮЁ��-��>�������!�y+�������o��X���Wl�7�B#ӏ��b��J�@��cV*��d1J�q>r�������*���<��:'����_cbB(��l�ɖ���ز�|Eɏ��dn��b*b1�5�D�:����b!����O"0�;��m�܆�p��ox[B�m
W�8&�8r���e'N;H��1��K���1Li��'9͎��H�P�0�
�~�q�����F_�UH�$nЋ/7��|e�Ki!Ì�vd���x ppb�3�,K�QMH5��S�k@1��G��F��	�p��͟�CG&9�kV�Nh��	3����,�c�I�B����a%�	�d��*J����4�q�2���)�!{DߣP��p<�}A����S;�-	?��qϔU��;!��Ya��%I?�b2lD� &vA1�w���J�X%�1(	���!���0~��|��J B˩��|�*
�@��TO}8�D!8Z��A���^,�=�j&b���	�P���_��2XAG��10X_�=�z�n=r��s�����<p��JD�#0DymD��ߌ���krϔ\E�u��G�	���
GM��� ��c��I��j�,�r"H]�	��0�d�E��o�G� <r`X��V�I��8G:��o2��PqEV��ei�����ђ�VO~��\_߱ECƱ)ƻ)njU'T�n�v����qb�>���	�r6ST��a�$�Ƅ?��(�V�d+4R ���������8����������{�)�Ǳ]�GS�Ad#����ό{���Ć׮S����4w�ž�>���4g�goc�~�7Z��24�����E}���+u�Ր�4��B�$u;,o�`'�)^/[��mb~;فPr��&D��L2��Wɕ���e6�� �Y�"o�F������xZ�K���8#7���.�N,&��62�k�)��|c���M	�:�9ݖ�PҶ_��S�؂�\��#:F7m�����)��0��������W��Y�Ԫ��lu�ا#�����d�e�t��}��}R?R���2o�?���T�Pn�ZCpVβ�d�9;�� i���5K��y�j{U=V�����p�h�0�[.:RC5������8f7bM�Y���BM���+e��>�����ƿ���>0��$�� �"����T�Z�}ᾮ�"�R��G���hV�Պ9r䫳?�:��T�'�<�h��(װu?��� �J�j��PA��mat�S�5���H���Ye8�Rj�;a9�C�"(��d6p� ��EC�h|`�7�2ڵ�< '9�Մ|�>��q��=�֩�#ľR��&{��nC�Rf�g6]H�ӓ��}��,�c}���,��4u��T��,+{#�[dBM �dԆdC�����iD�\�407�� jh+�t_A�`WX9 m�r����K_��Ν}fw,\�8�ZD.��;��#s4뵧��`��m`�F�J�g�WR�oJ�y ��c����/���+��b��׭��5�	����JSL���+'�,�} [��n���W�į2>I��LUjMNLj@ K&˔62L�/�=\��1��t�yJ��!;u�;B,��"�,�g���At:���9;�S��Y�Vc�^?���9��w�������رv�I���r�E�~�H`h�d��h�b�E�g^�����pB��lӱ<�#�L3�3��&+������
9�C�]�q�jp�q��C�d���a8���kJP�~qk����Љ�Gf�5"`�/�U5��.ҷX��y����pZA�f���2�=��F�֓��ݪA[huT7GY��4���P��_S�T�PDruC�s�1����`�.��$E$4�}����a�P��f����0 23��n(��k ��A���X�uv~(�w]�_��]���!��ɔKux�Z�=��7kj�T}���L�+��t��,_��HeZ���C��0�v�oo�oi�3yT
2Wǌ�����ʺ,��3˙h��cf#VL�ԤV��r���Z��C#`��vG����+9����Z��P�{���> �' U p�G`����4�~�a�����L��-��4�ы��k2Q ��o��'nǃ#�~�N{<��
 *@A��_�3��0�ґ(pF�u9���T�:Q� ^��Zd��=���kp��q���H��Q,k@��
&��{��O�k���$�<�g�D`F���W^��˅��"8���v��~C�E��׵�P�Y�X�{a�j��!J�N�\\Q-tS;gs8]v&ڨW2��ߺ�v�.�k����Ԝ:�c��� G7<~,q�,�|������}�bN���:�.�*�7�{h���j)��Y�/�XgϽb� �o����/�YKcN�_L��:
�0��@!�����s""� b�X��t�\��h9�'���iSwe�Ζ��	�H�w����.7�.�9�-�[Y�˼��/����fSf�7Z�(�1;����I�}�$򽜝�n �V{���d ��e2�01^��K��:�>��ڄ��m��||u.Ȟ�m�n7��(�/�#f�Q.1iB�|�� k���U �̘g�E�Ԩ��C7.E�j0���Sp���̦�:�߁�osO�E��.N^0���p��.�3�B1���=����
�K d�UYu�r��ٱ�5{��2����F�:Ѽ��������񃣦�]<���c�F\wW UAI�Z)���L�ݧTf�s/��#y��y��D��XAO._�˰7�s���do��;�k����G#��.�����}ι߼iե:�cu��'RԌ������,4��6*R?ؗ�Ϟ�#�%��d<�:��A�����'7���Lc	����>���N�?��9J�{�%��U`[���K��tL{{������k4�ƵRb:��#i6�չDrw{#�7��>??���S���+���ܕ�s��Q�?>l�C��z�����=����(+{��yẄZ�1�� g3O��3Z ���`��wO|CA�q�e��������m=^V����ʽfʯ�[f�1�8#Υ^@AњA�~sO?�Kn��⼁ S�1IQ*dV�ӥ�����o���$9�T(��g�I�|g����(���N�YG��҂�p� Ĩ� `���Ԭ��9v4������;$�}��l4���മ������o]ƬRf�=��piȒ{❡�u���A���́3�v�i�}��u~�����;yc����k�N�рѷ%ɔR>�K�J����ٜ!:kkZ3�oU;?Nl��㳬�k��ԟk�5L�P���g����"c̏W�p�/`�H�P��S<� �
X~�n��%�q�;A8tF��VZ�S��:�ݾ�;�gble��/�nJ���M+w��=4���������������j�7 Z�c�Eg)���* %6��tF���V�*  ��W�>�R��C5hp��hև�ё���Y־L��f�ˈJS������	��qb�t���[�F>���!�˰�Z�-G@��^�.�,��=�����0�`b�9p
f��<��'�=��)ʝC��hp��`�Dv��e��jJ���{��2v���_լ���tГ�:�a��Nl�k֒n�,'g59V�=��rw�&2"��˥��������w̞u��*O��yONO�՘.������b�4��b�u�ǻ���G���,|&����X|"߾x!���6��(�OF��x�{m\�b��8|�!-27�lK9���t�rߺ�s��*r��TG����\^~sIB�U�����jv�μuG�Zb>�1�������/'Ǉ���/�D�Ț���3 ��Zmy��R�����_��$��ѣ4�����z�gt�#:d� ����E0P�5����^��6ՠ@'�`���K�U��N���F��ӗ<��~d����,^�&������ق����X�j88Udk5=�z	���\0��<8��{�2���EoS
������#p�aW
����&h��ձ�5`-���eS��8���*h�a��u��0���Q�ؕ�K|�Ћ�:#H8=;c�z�bP�6��f~�����p� ��?�=��\��v�=�TB,@�M��9t���S�[U40^e P������,�|�h~����'q�	�E:��da-��|���veu��ڭ������Е�]o=ݱK���B%G�:[�ɚRxn0:i�h���Kw��;�'۔?�I���{�W�A��d��G�ӭC��oLa�m�:1��D��'�P�sLI\	~��ſG�Ew�����';���3���7�c/F���+Mv���lH�1�/&���:�"<p	%�d���X�����Z�5=`�Xa  hA�J��9�L,Z�0�xзȜC;/�����&3�m̹�,Q�(��t�O v�H���7�"�	0;���`�&��޽�04 S�3(&��OD�L̂<��r��p���$�q%��q���Lt��V�z��<?� �����l���ԡԉ��a�9�A�dN�J:�qJp�fá�e���{jXa�`4��o���wMp���:�>g6����;�!b�Y�4!�C��@���l��J�~��X��r�������0�D�Fjh�8��_M@%����%��Y')J�S��{R�=0� ��ՀC��N��q�UGf�d���i��Rg�'H���)�|��0xX/u?����ٱ\�щ�XJ\ʸi��5'{�F{�k��;�+�����P��4R!]ɚ��yJn�;p�w�1�6�������`\I�*z�(��g{^Cs� ��Ki�n�p��`V���r��k���|����Z���O>����c��g�+~ʷy��G����ru����؟�<��s���C�&t���93���㣃���g�y���^���IM�F���D�X�����c�����7���g]:pm��<�'�O�l�M˪h!��x�������f�\$>��OO蘑�B�kQ(2���@�H���ދ
NQ�����K������>[�DV��$&�Z"��/���O��Ρe\F9{M,�:�H�65p��^�����:t�08 �g4&A�(TՎ���t-ƺV�7���S��L�M\>�ɞE�'q����L�l sn��>b�ZP��$���lmF�C���k�J�{�DYK�^��H���2�kC��D�,�֜���w�6 \�K�zA� OrN����G�|�i�����d��f׻�^?���w���q~��C�(=��ye,%���GVbL3_ <]C��q�b?���فf��F����t���}M�
s��O�1H�.Q	@O\��ޗ1��XE(V�D��=Ůe�9�2��������ul���]�ׄq��QFE�� ���1��
ңD�3�X�����"�C��r��V�
�y�^�#� �F����A�^_:cUh<��N���=pr��� 6��k8��`��^��9����5�N0��_��-v�!K�ݠա_��GKc���wƐ�X�N����V�^�ٗ��:��e# v�6^Up�?����$^s���\�%�OB��8���@���Z+�1�j�LjS���('��s�2�����i)��w}kfڔ��'Y4��6�- x��v5�5u�A 1cf\��l��[&^�,v�j�F5�.n[Z��[���)q��M�ӵ����͕��Ԍk��f���Vg,7�{*�!PA����D�����\_��m���C9;9�����/�G��5�� DE���F~���@>x���H�{���JkC�[��&��_�zɱ��44p���Y���[�ݓ�^��ACN4(C��~>��h��ۀ��#]�=�OO����K�?�D�i��6d	պ���~�A�
�y��z�:Fa�M7&b8�%.�7�+�Yo�r*s{c���3{�����]��4�q������RW��<hARN�=�X�єJ�N�T�Vĉ���mk��k�A��}6�����L�v���t,}�pt`^�(�$*u�l|�������	�9\I/HL����_�w�l�L�+b�V��m���r�fړ��w�~�t�C(y�����������u�?�h�w��cY��� �,.���Ai�����0��l��b��rj ����^]K����cj��0x R	��k��GjD����(
'�F1hf1������]��-��h�+Y�
��|�()����5�9~����{�\��yγG�Cغ���UVRF���Q���X`qǉ1B�|��@�@�qc0���ɒ\�xp������A��vvv&��Ȓ1��0�E'���(�΢\��-F��f�ϟ�Ǟz��*4Kf���j��:�X��9����y��f�5������� �[�[�k�����{cP�S�� B��"�Q�1�d�����$F����r��ƉՐ�T̀��Z��_w�a_�[�j��d����;��i���u�֗�P6@:2�a/'+f�h0 �hAJ�8J�%u�j�ɖ=Rv�3�Q6?)�+|�1*����/��w�k�3���\��]����S��L���.��{����i]:] *�\��Y��i�Bb�d��}���+u�xyL����Z�wW�n�h `�7�]����S"Rno��k ;Չ6�6%1�hvz-Wo4���)b�(��O>�6��a_?�\g_��kz�6��n�Cl�Ç��������7�fͩ���>8�3�8��v)|�p3�܄[���NZ�Ȧ\�=a~�%��(��Ǆ	Z L�p6}��`�=a��5��v!����ǤO�����mF��y�;�]v�&�ދ��qY�ۧ"��I�.+��	Jq?��o�rO�`FԌ�Y-3�L���|/ۿ�#6&8A��=J0���I��dK�+Lo/��51��{�0A�����{?�<ޱ[���Ȇ�p�_,�6��^"2��X���O�?��K�-DN�[,[�K���"����;�F��r;6�P6F�z�yL����]��Ѝ�sA�6��͉:�[��r���<2�q��߬~�\삡��@�B���2ZkJg��E�[Y	�3IKpa�@np���<�1Jl�$�@pC���q[�yT�ui��IM�f�O�%A{�N����ԙ�43o����f��s��B���ǇC?>9#���յ��6�R �B���`��O������Z��rrq�=���翐/�|-�фhe��
��Z4k��3���վ�{�CRɶZm����&�_B 8d����H�Nf <��������^����pBpZ��5[��g��2�P�v��{��ɳ���W_�7�~G�������c��Z]��sZ<�`���ű���!�ŷ/�H0$�.^��ν|��Ş>=�8���)CO3���[��"��n�nt����Cy�����uI�zz~.}�!���k���P��V�(0���'c����a����@ۿzyɬ�� ｗ�T^��������w�m�\�!�u;�{���b�����Ot��0�I�9�ա �J�� 0"p���td㉇�71��.-~��z����s����Avwo�F%;������D��|f�R6�IY���	�$O���/�b�k����i��\<�ǚ��� |��%i������4�Nu,�`�`��XZ��&2�6�b3
&3�)�	Y���W�h.���I�¦��a6����uM` �p"�g7��=|�o���
�{qMR�	G�2������4@r�8t{�7?��W��ء��Ev?p���������G���a��rE��b�dѿlESP`��i��mӓ�l�S�~���[��ـ�������q���?�����Ei3�,��s�9g��kS�s����3x�s4�.B�\˅*�T�� ��Se�?{���0{�9b,J��1��m�k���\1��`���R�2��B^b�ȲA��m.�U"����'��ђ졐�l�#�~H#r��ƞ��t�Ԩ7dO3�S5���@��8q. ��N:[*9�5�����\��Gr�������%�;u�.5T+&z�&��z�`��hH���)P�˘�h��~�ËG�TFÉ��>��77�.W�h�;�1�!T6ԉ5�1�ի�.�0��J>��7�������Iw��Y�G���ك�6(lr���/��Z��+]��x^z����?$ �?z.�jI������f�
IBu37٫�W� 2z�l6/Ϟ=c%���_�^��ֵ�y���Gl4��7t�x�N��q�/��N���kҚ����jh�>�GMih@����� �5k}�䑬�D�n�����&���;׷W��3�Oώ����P�+�X�b�K*[H�ΐ����;����9��:�gB�ac׃�E	�ZFۣ(<��U����CC@�_�u���;��ݽ�*%VU�����/^����:fd�h+��A�:�AWt�k%�Cuu����o���O��Y��c�/d��������YC��:wŠ/�_؋`�C��Dw��
��&x��z����z��)f�.x�Ls�4��1m
��'G�V����
d¤(���L�+�Fe�q�4}�_���7�vw�)ZE��C��}�%U6�%>@��s�Mg~��;��v�c��Ȅ��N�s��L�c��T[��}�����g&�b}x�5�!�V�ǿXb�AqFc���w��]8�ʹw���:���r��{�[�7�6�x�l���g�X.6�s/EK���Ã��l�{���nJ<?�3'�d���	�?.^��/	"*��EI�Y
Cԫ9}�*>}��G,��^�˛�;u5�32�8O�	c���� ��ɵ�F���@u��R�ٌ��6_I"�L��>|-�@/ޙ�Z��i
�!P@�����'a�P���<��ֽ|��~�Z�G�r�����.�}��*�����=�s�H�����k�ײjpr�I�4@	�=��:C0�i`7���6�����i�����f!S�b,�Rנ�+�޽L�3��X�ʒ�x���+	T4��i\Q�c	��c�V��p6�;�)��_~� i��宭;/GGJ ��x�� e�N-a)������� �AM� �j�C�`
�Lh��W��~�����8�
<լ�[���Ŏ~iN�� ]A�嗟�J!�<M��T���x�i}N e.ȝfA�}���ܶ��U��쑰@���+�+g2�S�B�q%߽x����8qS�f��{~�q>�k2�Cl�{�р�J����lM~xVh��I\+��K,+�Z�'��1 :�a�NK���s��P�r�ڟ��ry���:hTu<����z�<~�g��� N�?�J��
� �(�s�L��7�����O�����+�\^�w��t=n�9O�Zp��w�U}f����c9:9d5����p�)���_��Օ���A<�q^ϯƊF)(�QN>��S�:���k��W\gO<A�@��u�e�'b� *�a_^��V���I���a�	T�wƼ́��rjI��(G��Ʋ��������4���+��aUb&DXO��<��>�}�G�	�=�b&~�v���ﾼ�����������ޚzr�ձk+�n�HJM^�ZD�;Iy��~��߆�����,=x�)�Ŭ��w��<����%�;}0��������SOM��ds�V���eYV�*��He��NR�8ٔ�wK�~w䍧��u��@��B�ǜ:JN<%���Äq�H\o��aIi&wvz$4����s]��.8��j���n�d6��O����[P�Kc�:��YNT4�U���C�ּ[	�k���:p#�@XJZ:��:�R�*��#��Gk}@�~T����b��٣�����{�h�Q���\ B�$hi����}�~|@-��R�&U��e�2)Hވ:��$7�
y�k2J&R�
R��?.N�̋������(P9�y�OC�������b,)2�3����4��C�հf�*2Y��@�Q�xL]T��ah8ΒY��0~d0�0G���,q����4��[_�=^#�ȫö��WA84�Ejl��2h���{�=B�b��,����4�hwt�]�}� lZr���y�(��H��n27��Nw*���f�g6��8ɲZ��F<�9x�G�6���gH�2�c�MW�)����̰��R���|8l�R�e_2�#�ffH4��������l0�U�Hb���[�o��@����v�	 	b�,?s�p~h���]S�B�d����(���j�#e��(	�����+������@�k���������0��0j������7���g�Y*VnEƎ*A��cU k��R�P&k�w|�ͷ���J�EcNL�; :j�;��JQN5�E����ve�p�H��� Q��J;�t,�#"0�%���>7��,ypb؂�U;���]A/=c㲨Z��K/Y�;�K#�6u��|%�W��_�÷1k��F`�6D���H<P|�"0-9�`:LY�	�~��Z/T���qb�|��bjN9u���9�Nl������|!�/'��47[.��l�Y'�U�^ͪ�bZ��G�^�h)�D4.@X'o�n�-��z�ֵ6:�."���a��`¡p�lB���Y��@f�__HY3�r�)O.�rq�'��}�5���RɧR�t�$�ǧR)7Y��@���q��;Ｎ�(��	�Įr������!3^�Ƹ��e�r���nm�%9s%{� $`�Vh�G77RnTe�&���<{��|����7W2V�T�ϲt' 1]% � 3!���S�i�	��~Cڗ7����fj��%}pq�R?z҃N_�{yi6���PV�Tߓh4$> F�#��Z���<�c��	^�\>e6S�В@_�{a�i�|�c�8/8'�9a��Jo������9�@��װ�z��|mҏN|�����S@P���<������1�OqAk�r���z�5`�y���e4xbc���jD`�X�q�̨S�#��e�!-x� �G���h`�QR�����iA3aJ�2X��l��/����$� ����]�1L��x�* ��r*9Egb��$J�A��'�
t��F��,�3T����s�1�4q9�c�cUe)�+
�|�k� =vT:��C͵��u#>��n��;p��uZ�r ���z)�������W9�P�{������޵� ��k�{p?�Q,����#� �����՝`c��/KV�q<#=�[T��AK�X�h�^�g-Ԁ�%/^��뛖��ۃ�g�<��z�-��#����ͱcfC�<듃�*;���ت��?�,@գ�Eɦ�
��sr<�U\��	�t�����[�]R�ο��z��Q�%t�������`.D�1`H�$���F}�^/�|�D,kԉ/<P%�	�8f�b��٫�?ayY�F��ãF�T+�����{pp|uqq�*
��hM��OƝ��\���l��=�����G�`9@�B@|j����#@!�I�n�t���'�sFF@���b�E�eøϖ�CqZ�W���LU�ч��͇rԬ�Q�$�ZN��e�+eȩM5fp6�A/D�����C�v4�S�ѭ�f� ����He6���P�$_`�<b�<�u�(%-l���P�\�9�H,�'��<���ԞP�ˤE�}�F36�|WSA4�}ʹKR��t�%�,�/��L���,��r���b d�XR�+�$,�D�5�ݫm�@3�R����K�iP�`�@���qGr�����F2���QF����FSY!@倔��e��"P@ ��k&��4xl���D��r6��Q��5(ZiVW)չ_&j8A`n
qI��Ζ��t3Ku`�5��ѓ�'X �"�1����I��|����gd��C��X㾑���BY�,��z��O/0n�AUz��k�A*�Dh�s���{���"j�	�yT0 <�!�	�ipƃѱGX?��Q�u��ܦ�?���|�ςAX���,�Zx�l���&�8B��	�٪ժ�rZS���^��:�3�9��}����7@�O�< n
j��Y�*��)�Ԭ{Yo[������|�Ya��J'۔�Z��:��!\�v8�^wJ�[�[�q�D7��Y���T�����]�kf���p0��p�{iA�t��Q�.����޴�R� o�3T�{�N�����RW=�3�?p4��:»���b�4�*��ww���� gT����[*ur��#��J�'>L[�	��-:s���*E�U�0�����Q�|.�Q/("d#�s�B�|�����4���ۤf�3��,�p1�;�#ڎ,�ytG��'k�����<�5�({���o��U�h��<�mEe�� 3*��7?�)2؝%�@~��2�Uɽ���~��aЏ�a�Z���ړ�Щ&�iV�����3]6�5;��F��f�,V+��g_<~����?��T*ݿ���xkP���7�����������/��0͕���a.;��c/`)fc��#;%K�(Z9[�����u�X26n�/pH��W㙡OH@R�և*�� =n��s���<h6����SR��ԑ�W4���A�!�^K4^IIӻr�He4dd��� �����N��]���J#��u��4�����9�i�y8؏tc#qlP�hE���C��gX�ܵ�+:��jf1-e��v��T2�D������k61}[��V�iM�/JWj�������
4�>߯�f�P_}��DP�b�ݳE(���*˕"EQ�[MG2Q����g$����b$lǨQ����F�}:D�["D�t�Z�\��Pk͵�:V�R�j�LPx�G���78 OJ-jQ�����w E=7��1홬���o��G�Q�$����Qc_�j�ѷN��&�%j�Lw��tֱWű1����m֪20J�<�9O'�ý�2 Z8jS������ *EgQm��<���[����̠7k���.�0��jV�Q`$Q:61&ü��mbU�ؘ��^���k��� Q!+�L��\kc>�x���AYl�b����\.؈�Q?3���¾>��%�l�p��9)G�;K�uhT� g�wⳖ�#}�$��RAn刧�M�:_��25��.0}�L�}\��|�M������h�V'~��o.� 1��h�X_ ,I�;Ko4���-�oʍBl�$��@[��&�}��1g�QA��c���a�N4HC ��N<��p ]|D"^�����;���iY���{�����,^�1�46�Չ4o��n��'d��4Hl��$1�Vi3v	���`?��61��IH�M�Qrs ����r�m�r'�0s�J��_��C���W�g��kV4�͗��督�#�Ǉ���F��~E�U�m�?\�ft���F�����ֿ�{&���>H�����8.��)�����bf(�/�*�s�_�\�<F&e��H8�d;��_D0���$4E��:D�\��
��Ƀ�p����.��Ek�c,�\Rg;������� ��]�u͌���rUn�RTf� V�LW#�PU��u�3�8���^�g�Ayk'����y�9��NQlh��ŲVb�y0� �H��-h@x�Wk��e�p1ϫ׸�d�E�>O�kf�Yk�:fL�
�/ԋX��Q�>�W/^m'{'�t�Cu�_��g��N�ప�VC}�>,+HG��{E)Y ���o߰�#�y��zM��s_06$	��O�>�����5���^��P��V���C�X�jz��u��yu�Z�]_�A ��T�ܐ�n �(�
���ɍ^�]�k����@4#��s�k@��H>Z'z~l����5�Yu�*B�E3���cr�ÀQH�	�.& J\�&����9����ϰ�a�}�������z}�}�`�u�pA�&�x�a�c��{�(����F3cI�x(T���*$�x�D3w��L�S�{
^�S,f�,�G��b��=��jU)�߀���@[D/彪��y6@Xv5(Nf+��b�0
�j�X*d7F���G?~��2a�s�ۢ�H���R)�y����C�R5�T�ZҠ|��:�0��k�D?��ya���B�f[�Q��J)Ǭd5ԕw�O�C�� ei� Wc9��-�6���?^}�8FN�z]�3Ña���u�����=u�zo�n�6"	�S"�,���r�]�dG��[������ �5��B����Y������x�A���
���Z��F,��n�Zd{N�|�l2{w�M���T-P�A;1���_o�������8�+�	�~c�����o��o�����0��
Ǻ`7���U����S}���W�W��8I\*�r��	�/t3�lZh�7G���r��nT_,W|0r�=N,#�c��M_Ŕ�'ik�͢�����
����'���(�3�$�횑:�!z��uc}����@� �H�X�iA֐+J�P�5��l8����l���,��mt3��M��A��)����^�I)���U��
t̴c=��n3�F���wcE
�6u1�Z7!��F{2�\�4����b�U��Q�**�p�)؟�	�`{���8gG:SG����-�o2Q�4�K��a���s%�t4[�Ԩ�� ���F�,����P�|ݺe�Q�!9>�g���s��W�yͲ�R�(�����������g�е����[�i�9K���8;:���︾Ӡ�ӢHNv�)�gGb̫���tX �!�/3 �o�$V�	������/�7�ܟw,q t���h��9�Ѿq�CQ웗�m';�[�xO��$K�Z�&#T;�=��W/ 캺�G�����@��ƴmA��^eO��/��mY^]���N��q��S�����X��y!0�8N�ۓ\�3�@&t!���_pd�B�PR���e�h(�������u�!���NJ׉ci{۱�d L��R)��XG� �6�
�@��}*���A:Ē
`]LS���e��"��	�c�b�S�C��s���V�sc��=�7��d[�{���P�x�vZ����Jރ��9���(t�ųg�_`��z~��F�b��T��t�D��T��w� �,��3����Ή��.;l)��`��h���hgC=����"$G���0o<L������wԿ�pm�á$�d���h>H��5�]"����=���O�<�
�Om�<�d5��?<�>�����������?�����O��[5�����;��+���t�MV�^��J8_Qw8Uc��N[#ܵ�,���`�}�儊]���+��D6+U��ðE�	�$.��xH�J8ԸN|� 0� �ѿ[�ĝ%�$�D��I%S�y�0�}ז�=�L^ �����ܚ�3L$TP�޵���"S+�<?8s��Q���O�b��>�	+�AٕjC��5
M}	��e�P�)S���FAY2U��q?+�^*ե�p^�l��ȡf�<��3uT��7 dC�h������R<<"�z�y��?.�^{�Z��y�kV̗�T��G,��'W�z��?{����c���йF�X���ۯ�ۯ^J4��<���|�����"��թ��r�25X�(�rsu)���4��j� j�3u�S�Op�`�U˔\5����Q�7�����jP>���5�ٗ�ܲ�v뎙(g�5Ӝ��/� �(ٝf�O�Z��O�DN�������ӹ��je�&����fM����~�����V����5Q�Z�Nh�����u�Fd���u򇍆�Ìh0�Ⱥ pr~z���.�AW._~��)�'O�ɣ�OXR�{T��E�6=����z��\���Y9�N�O��> �*z��9�)Y��� c����~ �
&tON�9Nԡ��g��O�p��yq���Q�C�t_����t��{��B��,]j�Ə8y24X�'�#o{�U>��x)��U-������Sy���é��纮iv�{m���{�싧����<8�`�U��S N�q�j]'/ՉM9f���^oY?����W��X���__���0���� ��t}�rvr ��y���t�]��RD� ��!�E
�G����ðo�j��Ñ+p#ItԞM!�:�o즡����t(����=s��Q&/��Y���f��qI7����ر�I7���(=�x�G �-A�.�I�n��~��M<o�����(��5���}������/������W��O���D�����z���&a�dC�80x��x�W�En�X���\$}{�c��$��K�c ��-�0�{�^�gFPy̜/^�F��2�_�X`�/��*%H#	�:��آjF��������FT�r��P�jp�����$v���6:4��#�K2�ࡶ�΍-9-a5��Kg҅i���H�<�m#F	�; }��2sA�P����̙�j�Y�؀izdk�����{��A�2���P�:ٜ��D=�@�Q����#�FO� �L��-�Ӂ>כeyWd��PQ��������B����1��YP��P��f��=�������d�^\�LV M�q�qW�[]?�u�}�����9��4�l�]3���u|�`�$�ɖ:d�������Ԡb���w�B�%f !��9H�	����ɱ�����`�`)��}u`hP��0�ueܟ0h�e����J.�9�y�o�� eHK���jГ�:wT�
pX�&żw6��띃�(�]��b��{7 ��@���H�>���P���T��2p�ȂA\E�ʱ�����V�V�U���d0���w~v"=��;���; �-:����=�=Q�����v����-�o�赵��qG����c��alj���t��X�����>���9�������c�/^]��ptM���K̄��4h�Qu�����^�"�y�� �ToP�zpq����A�4[p����@�)����|��k-qZb�{�6�=u����]�8�\⽤~S��G�@Qbq�����m����MI��(�̪xbS�a�X.gO 1P�zM��-!n,,u�»ʗ��ɞC��v"`��8u�s����5��n��0�%��=-]���/Χ�G��w�G�?���������J~����C�9h��5g{�d��Y�{+`v�C.�z��f��ל��D����WW��.�8'>@�8	���14�Q�	�Li�۔ji�XK��ܨ�І��D�&aB�K�y<��6t:7|�#L� �y��e��L�G<�B�+���?�#�0fT?����c8}�䈱D��(!i/�`@�j��i_��a$w�[i��2<���R�{U��`�����}��D�zc �@a�����������i��5�ٗG�|�AK^��@�CC��ý�:��Ͷ��t  ��G51!�����i $GU/W��C�E���4�Yލl1#�bQ�vFa8�C5����p�rA�%�8M. M{z�U=V�2�h,/��/���R��a�׮ϋ8��*_茮1�Ä���^��[`�&8���~�ZjVp��`#l��k�1$���?��A�eݔFʉ��&C�4S]PR��N�\ �ghea�!��������u�]�wC�i����~]&��"!�#F6JeL[��F �yd �r�������(��ǁ�^�}GA�Fþ�#�R1�R��f�h���\��͕�o,Ş�$���=H{�{m���Ϩ�K����7��D��@��������'��^���q�\���|$ӡf�o�r}u��U�>�������v[=r!�!����Z���Z:�7$B'ó�C�;8�-�0�A�N�ZMK�ꂑ���z.����1i0}���"A��`��n�Vi�BciC9���9���7l�a�FoD�4�l-�:���� �����I��*؛���(�2xb��w�8>+������L}��޻�,*�L�܈���l�'q?DT�[~�P���{��(����?��ӿ��?�����G��� ������O֡G�*��w�R�敬��� {;@)2b��k�L��:zҝ��o��a�Wܜ����=�n�:��y�:Bj�:M�(%��3-b�3ǈ��`�v�t��������c3�D�ڌ>��@��l�6�<��׫��k�7fi��02��8*Y�ΆۙN*{�o�)[a4e�L��|4�t5V7��7���ci��'^P%�Kfں"t| �������2��~J�6��0_�Yk���S��g(�P&���P2_J��Þ)x-��9�jmON�����������|8>T�#�ja$�P�Y)���kv��f�g����9�l��Os�^D�g�艑��Rm�%���D�*F��Nҥa"�&j���&���л-h�gI�
�cE���NȀ+r�x��XҀaO�I�T�:Ќ�s����(h���7�e@��h���Tʳ̌s�c��J���g
�k �MJ4��ƞ�%��9<�8њ�mI�9=!��r,���g"j�G{�R�Ţ���s���p�초��l�r|��D}��D����x��{�[�f�O���	~T�y�q�ǚ��:��ajԡ0�B�}8�%���g�L�Μ�U�,HdP�^�l:�^{�=b����Yq�0�<*KX;���5��:r{s){iP3��aW�sJZ]�>��އ b��՛׺n6*Pޓ�O�z��A�cl����l�yD�w���G�������j��* ���	�x!�А���h���]r�K�Q 4>���zT�L����d��b#������F���������iyH�a��L���.m���d�cp���(�����/���G?�����W��d�:� J�L�H�#+��_Ɂ|:'�jF R�	+4ǆ�ځX8��»�:�l%"u��t����u3́�O���wFl�ȳ�F���B(<�E��qs�ě¨�,��L47#d#S>[�~�0aQl(����/�,�λ���b�ȡ���8�8ȴ������
�wZ���?C��zA@6�0��6��	6)M�Mv�檜��p}����"�HI�eՁ�5���22���3}�;]��ɒ��z�>�^CD7��_-`��o&�<�0S�L57���G�{��c��1��j����7K�����qÈk9�X	6N'�Z>?o��򖘤���ȝ���89u}Dk^9	oܞ[2WQ3�M���J$yp�.d#Ɛ�d]��7�1�s�>	V_�������L��]�S�d4���5�c�ߕ{�ν���߹��#��o|�}Y"�?����^��+�ً9���>���۷��B6�Z��<xGkͱ�^<{�.帰	�q K�F{{$�w�F(�#�����$a��π��)|���[B�c4t�D�7���2�c�կ�}E��*q��\ǭ�Dk���]�0o��r�x���w�K_����nʉ}��F�!��c����6�1��r�������p�#�im7l����>��vYO��z���4z`�#�_����-H�d�sl�v��Tg�X*d0�i��8y iU�,�Cu�"G8b;��ڿ5v{7o���+�Xma����\���$�<;9�6ZAY������e#�.tW�E(�4��,����v�did4od.`̃nt��݆�;��o����auD��!J���g�����uz��}wtx��S����=|��e\��*N�i#�ߙ�˚xt�]w|��3y^ H�������y�+� � �}��Q�cz�Il~�@��ƽ)��A���se�����T�yϥ��Y �������ב�~=V-i1���GL�=>�>����ӽ.$�>�]}�U�ӟc,WL�K{e����鋿��o}��~�������[k�CU�~d9r�m/R���]�-�)��D.�<�l�U����N��u:����-̥g!���N�*��]"��&��W%1�"�'��KҴ^{��q��L���O��z�
N.յ�WK�-c��ԁ�;I^��A{�S�	�BH�t�(sSE:*0��C���0&�A�-�@U�:����5��G�Y,y�_|��]�rC�d��d����R�{��1	�p�^�#��+�>_0�*A�����˳K*��X�m�5���{l{iv+w�{!��%���4�*K�+��}�����2�a��o}�=��!�$ՂP��S���{��D���������wu:q=�FH���������5�1�qEJF��?��8 ���F�?JD8��Ϟ�=zp������UN�B�����=���ĝJd���DHɊ�CQ�~�}��_a�Ս��������?����}��>GG���w%N�$)�A��|փ�!2W3Zݞ�|�.Oϕq,����S�;������D������|�>���:X�����W�IV���7����w���������?�k����Š���y]����n��{7��]�) r��T�����{���c>��# ����cBg���OH�#���~�% �3>@ZZ����+w��5��,'��89:��1�FV�ރ=���y�5��}ā-���t� � `P�/xxS���=���dyE=~#H�!���-�2c�.!���'�vw�-�W����Q!���`�!!#]�O�2��G��hN��&��Y���v���+�L����I��#��ܳ<��	M�T9�z��$7���?���D�ዒȼV�j�Z��HD�PB	���
�&U�������c(�� ����sTgDȐxL������{'��#�11�J��l�(�}��巾�w��G���?�{~��c���4��%�Be�笢��~S
A2�{Z��kR����L��Z�6��!e���� r��9Bp ���T>S��A����J:Y�]��(�<�?�  ��r�u�L+l�-�Q��E�v���ڏ�X=�V�>�A��E����W'v�S�<hɂBk2�UK,dkSO��!����A7��ѝ
���&m���<�[�a�a=��L�"jE�d���;@k�<4W�K����-�b4��rr�p�%��j�|"pU��1B���i_~��(���D4��O���DH���;�ϝ�eF.���#H\��[����={>u�����D����*e:\DL�o�/=��������N8� wz�QF@*���B��5h�t�9��������܍�"VʦHq`??��H��ݛ7�BVӹ^={�~"D� q"����B���T��t��ɶ�د���������c�D�C:}Wg����@=�ƍ}�c�|>���G�n!�l�MO��T"C܋]9�}��͒�&td<��,+����Z��s��M�LEM�7͜��0}�u���tI�uD� ^�Ƭ��xbp�O�3q:��QȺ�c�� d<��9�l,FL�����;���n?��O��OS���8� s�����/+���2�Y�խ��~˽zy�>{��[Ŋb��0w|���AN���3A���5�r�?wǇ��v�c=#��yp�}w��;lÍM�!L��C�S�_���]-�up&����ذ�_�����;��@PI��Ha�L��DgQ0C�i#9���4�=���6��P�ap�k����^��}7�{��)�wٜ��C����dTm�SSΗ��U�2��y�AD��h��7�W����T���QX��z�����:�]e�W�|�	
�8M�������?�>i�u��]rl[��x���$��N][��h(�������t��������(̑(���l4r�6�$j�)�s(c�p�h��������r�g���,��|#<OXyګ>�kmq���%�o���t,#��m9��HU��WUz
+�h[������Ή�ƿ�ܺͿ�=�`b���Тt,�B"�ir���Ȍ�ヌHe��0@���m���4`�g?��^�Q�!#e��}��%7I��!��U�17^��T�-�bU�K��l(�{#wG��-0���oC~2���b8_�����RM�1[P�����rz�v*f-����ѩ��:���;H�ǌ�gV�L��u���)S�h���8�z���	�HOf���lȦGZ"�1����Ģ�|��[H�r�I�Z�$��8>%�*�_ҸN�'�\���C�"EH�B�T����q�!��$/�j�1X�3ݴ���]R�-�9�'��88�ɕD��<�3j���%-��FLN�{��W������>���)L�����/_��W/^0�z��[w�;}�,w|���Wtn�#�/Q08l���/��;1���1�c��������ػAG)��/�ܳg�ܓ�/���ݽ�h�r����{a��]��Hv9���g��?������,)�}D��9p���}�_r�,(����/�x"����F�d��ZE�� "YSְ�5�����'��~���$�B'��� �S��x�$�.�B8�3K:Rr��]�\28=���ݾI�7tX�ݙ\_�D��1DG�T�k�� ���7_p� ��p�8�������y��km�z��Z���ٍ�^���׬}��o�����|qlo�}�◿4��~���=x�ݏ>����w�+����Ț2�^��*�'��`N��M^+��e�T�:yG�d
�ʦ���kG���k5�̦���	@�����Б(8��k�=u�;�ςF��S�
5RE��˺��e�>g���z>��������$�6��tL�N�Y��E]��5{��;�zF���(U��7��n�ξ{yyNNA���x�98����cW�5d�R*�f�W�QS�9'I�4"�ʗ�&��L�Od��~�{�m�k"�p�3�VG�R���W� ��+�v]l�.alҘI�e�kqC�gdH����w#��шEfA��R@��n�a����w����I]J}�l�ۣ�N�I�l�Q�m���熇�����;�x�JE_��`y��=7���d�\0��|�1�H�C�K����
����{�*g]#*BGDN��J�eO7Pnī>]\�c��s��	��P��h�id�/�s��-}1�b��D����z#���1>9%L�49��n���g'G�&�J�j��-k>3 Zy>;��*W�i1�Hl����_hHL�È$FH�¸��/���f⌝����pP���H��QNOt�0G�ʱ�:-�@������2�!E^�M(M�{������k���s:�6����%��`Ē���86�ԉ��A����׌V�{�o�bcP��>y�"eL
�A���}��/�������S������)��3`�Q
}�W?��}��)��vvI��f�"u��zB�2(�q�N/c/y^��F�'ְO��(G�A��*<7h�[�ӈL�b6�Gz})NZI��h;D.o!룄���Ld7ю���\!1m�Yd�9�M���1�B��^v/]3�]��z����%�N9>�4|$�w�}�߾��/��������s�5�uU��[���t5nch���z1M1��گN��6R���1�M���x}��k�N��ʡAv��T�b�ϼ}HQ��9u�}HY������tZ�w�t���X�o��~u5�{�����������׆ԅ�3y�-IN=&e�ה@�i��bP}n�`�&H�H׃$�|З�-a(y>�  X6��F��:@Ld:��A�r���c0�\>��ۙD�5S�;/	���3|.R�Qp,y�<�wd�G1�9�m�WC��/�<���r=�C�1���@�-w��Ǎı�D>�_�c٬����߱9^�O���z��~�+_s��@��U18O�?u��C������G�X����{�޻QߕH��'���󗲩\�!�cr����Ky��=�G���:�s�셫�������q�����q;��������K�y RQr$�� 9mm�=0��<m��/��keN;@���Mq0a0�r�mt0 s�P������
���iԐ��6���SYI�X����x�Q��=_�$c�S�ƶұ8]Vj1�I��h��Ӡ��z�½H]�쐁��p8�
��s���D�8�Óc�.�ϓ��(]eR��&�D�p8���=���1��P����HE�>�F�7n��-Y�ۜpq��%3�GՖ��܏���WS�� ��"�jF�����3�!�b�������Ni܆����F�.��T�<�O����Pӡ̡��LYiI���ʝa.�������8�ǯ�����/�T�F�B5r�P�D'H�5Z9}f�Z7���y�uxS��W��C����{vK�[�����U!�OÎ�r����?��_~��o��}N���A6�@���Zp��������|��ˠ�Vwk�t;�ꃷ�s�*�X��rn��Tv+΀�����C�$�4 ��'c��j5�����M*Ԛ�F�5k՞j宥��Gw�ͪ�cK��բN����ѭ��ب����d%DN�p��;̶=^|ZPPD�3�Mi�q�$R�0�0�x�����P�r�Y����6���fɣ�4��^!��X���ׇ�X���R���c=a͟#jQ�TK�e��"�F���\[l"U�eǦ69�r�cў�l�B6�9D8p����w��>�����E�:t��aS�!����pT ��@y'Vdl��Pf�!Sk�v��!��L"D;s|q�r����>�{� @1M"��=��n���ћ��lI�A����9�=�;�oiD&��80�h}��a�,\Mj�7nw|��{��������K��'�Eݹvc���A�9�=�l����өc�����WV�$�ZWt�
)TLKK�S�2I�L���>3e��#|�_��w8k������jN�C�f4��r��<�+>�c@fw5�^m�A�*�}o�Ò�m["�ݝmw��C��顼pN�v��V��,8r��<|t���|V���/9���e�j�.TT�����c0�H�߼������Ϗܜ��o�ހ����Ȑ���_A��ƻ}]άW妘?0_�8aM�!���\ʚ^�Ã�~�G��%8�b"�Sβ�5�i��G��^Ț��\z|�j(="Ǿ%�
�
�������"<x�b�Hs'�Θbdiʛ��v�} �5u˻r��Z'`�R�8�7o�U���_��������o�A�f�6k�YKV#�C�ed�ǒc��(em$���711"��$P8M�"�����ԨYN�Ѩ�u�:͛֍4�jh˨�2��L�M'�HG���L#e�{�.E��Wd7�,kX(6�w�\�r�9a���´J9E׹ ~=۠��@՛��s�T<uz�m˃�	6��΀��۪*yH���*Hh�5��I>r�l�q��M崴1@�锺���gɓbΑQ��v�2���.0����u��8>�G�$p�M���ڨ�Ndcr��Es����=�b4#�W�S�e�!#�i~m�f��0´""�����	��ծ��� q�P0����87���� M	�G)W�����ME�B��c��@��cQ��ٝJ�I������г>�q��p���]14۷oR�s"��v������8N��F�ʵ��8_���W�1x}9��RdEU�41#ө23���u.��\�W��%�������xT����!tfi)�m��9�蹖�#\#1N�����q�Ǟ\��Ϙ�f�KH�J�����XD���B FU�H���ug�� �>��l[��{i���]lm�K1��x��~2�m��'����Š�r�^��p����j:i$[��0�>S]�m1l�4�ors���r_@���:�pJ�p_p/n߹�z5� <[X�W��t���+��� �R���亁��΄2�yP.�1�S��|NB�J�H�#��ﶃg�t������핁�Tu�cU׫R��Ěp���|�]�
�^ςm��c"��ehw*5iOk��ՌO��`ᔴ�E�>�~�@��P���gpJF�as��'�<������9�[kз2_��!�CM'�`(�-#��$+D Tc�62З0�H�8��q-m(��S�� V�F�ڷ�2`���jq[��M��6�u��f���dL˦��p��j���
1�ԓ����v��y�P��>�l���Ag�k}��YZ�!�/&[iOfF/�2/����'l=!yn6q��#FQ���>��ƀ1�}z��Q 6'�ks��k[<��b�����]�&9,�DE�W�g!B��a;�T������6��$��-���\7�b�ιǹ�r�8h�CWe��K�%wC��X��C~�|;�-�� ��^N�`QxN���7v���tb�8����\�3��\������a��^�`��=���-
�d�F��trf8[����܇K�J��BŃJF�3�!^���\�Ԁt|.��.�X6���W{�&՜�d��q���D� �4ދ��[�)�i�Q!�\R��A�B���ř+��\��ѯ�	��&���6)�LOQ�X���͝k�ı���_�Cq�앫/��ǥ�-�.��C����ƃ[�SeAF����nzt��ߙ��\�^�J&��FQ����79<p[�>�,�Oe�=Y�`g�sB�#�`�I�yt[��		��ݒ��#�b�pVR�?��B�oș�b���/e�^�)u��W�k7�<�,$n�λ����;��4�#(�>f	Ӂ\�N5��F��i۪g6B� <��R��;��s�����l�Jp=:���S݀U` ��W�Y��l�2pʘ`�n����ā���A}^��+6ً�<ܢ���n�=�w�2��Ԩ�}X?_�N.��(���UT������*뒥W~3%1c'ym�^b��N�!��y9���G��/>�ڇ�����Z��R����X�Q���WŖ�&�TwĆ�$*%yᎠ^�%T�V��&�j�st"�j�E�oVt��u8	1&�~��^,"ܘ�][\Z��;�4u_����6����Ȼ#ԥ���ԛLoΒn*(���T�ז��,���6b�~�;��<x�4����2�c����|hX��������\�,U�#o�iN3�*�b^���eP�Q�	Yh��L�(Z�@ĢS�)KߧL����N���5�+� ��l�wI�'c}o������l�荆��^tQ �"T%ѧ�zd����� 8yQ�(� �ƚ)%�'K6�b&N�l�،�g���Ҽ�t� �ɵC��:S�#���#[�"�cf|�9{z2QD��'�Ӗ2����D�4责0���i�(��^�
&V��`TiOԬB�B��0t'粑�y����!oVN��'�W���@Ք��朧T;�#dI������J��o����dS�"��x>��� �	�����=;E�!�c���cw~t@��v�A"lht���da����=�^�ctw (���,x��HM��Hr��J����٧;"gd����{����:ǡ�r�x��m>s�a��-r{d��A�&�"O��H���a���¡��A��u/�s��|�e����=g��T�O3�]{���.�9K��Ю����:+2�Q����~�y|K��Ut �8NQ����.
w���r��d��ж���,����0�`�+ɭL)xU\E�ʪn��B+������>��?c~�>�x{z���Zby�1_<�:[l�c� CR�PQ<�l�1�ɠ+�<U��ֆ�p����h>����צ�#oߦ��5�*T��|���ug�sa��p����둽[{��:��S���ʬ+8��c��c��]��d�֏�C�����<ޥ��
�1_��I ZK��k�뒦s��=:}ɥ |u\DK��>W<Ų	���..�@��1t�dם��
}��\�N"USk^����mBuVd�-gM#��Ө37�u�$HUM�QN�\���0yd�g��ϘZ��͠�u�p����l�RS�8bLg߅����#k���ڥ�k׺!놛כ�c�u����,�16s��ѝ�r���5:F��̇J���|@�C.fW���7z��NYJ(�fW8��̑k4zf�=����Fv�B�ܷ�����N�x�e?}�
���t����I|&���kR�f���0em-O		]�Q(#j�B�C"��=S.�n8;�96�V��R�!�)]*9z��@1�#�5�éD�'�309e�}�B�w�:;\.�x�e��\�y����0�3N�\���D�y��D&��B��|�������X�}C��h�yΐ׶�F�c�1	�;�����{⅌�Jc�A���QɊ�O�rf
]�g���:CC��hVm��u�6��9Π֎��,�� �emm����PZ�N�y����s �<xJ$0�9R��q���r�(YrE���ƷF=nm����,o>x��O����;������5���6C\����T���%:��Io���t�p"4\��X*�ͱMI�T\G:�j*����s+�װ*۶�:���Kͺ�:c��_k���j76*�G�(˞�,?�C뱦�x�J�%z�Z��Cw�o�f�h�?�RJ?&G~�6+l��5�I��-}����k�����S��$bӊ:��GMo[�#S�^�C����>�M)f��5�{�V���I�x�Mم�f�E�5K��z5۠�i�3�q��
8M��A׷�����̽�y)�u�����a�i��܂�6���6��m����:d�����n69�ҍWG���!��+������<KY�>6n���Y#��k7I�l��D��fa�VJI�������M��f��!btK��5��'| .O}�z��'�艶� + au67�9�M�8���ҝX�$_!���G���)x^�5�dh���A��g;a;!K]�s�"	�ICE��t���>DNXNY�Y¡�J���ا�H̸� ���9Q�EZ.N���d�#���kY�Fd���3��P����"��}=������h�]�S2�Q��5��ĒE��u�ൢ���J�c*hs�b�Ѳ�9~���M���l80�J"3�}�I:�lX\u'��dɅ�4ߑ�:Ɉœ�6Ȓ���p��e�}w>�S��NYK�B��SY1$�]<�0��G�M�m�~4�V_�Y+JK�m:5��1�5�c������̿�CW�O���pq����d���Z)C�C���itJ�V<�N��ӯ���jd�Qph���2^�����^��6R7�6����k��#�t��GU�"���K5m�Q3�����p�7�����c�ku�6[�x�`�����O�:,әQIK�؜���R�.뫞|����oKC�v��ա�~����j!񩧴�4Ȉ$<f�qT*���QW�kN�3|�%�`�v��/=ۺX+,���(�]ͧ��rD 8f�Y35��&ًٍ�Ff*�n)���H����sl�o�pc���G�Cw����q̬D�G�bXO�XB�Щ@S��F��0�����4�f%B�;�W8��=��+ǎz*��x��Q�d���-�(�9G��Ź�8�N��� FhZ�:�/q��r��cw��Z�$�WJ D&��]b2�*]m���F�)r�h�f�D��aЋt5�S�Lj���cyu5���#��Ȣv��>�r�5�UJC�zV@�ʒ�|k��Ԇl�-Pǹ�ԕk�'˺1��;��RD�>�$���	�>/4�-��A��i��x僈ӵ��h�S^x����s8��������M�t]B�]�r�3Yו�z+!0�A�cKK*�yv��2�|W�l����k����щmzy�|�dlڥ�SSȃ�T�"#��t6�g�N�-d)�cZ���~�଀������b���2�C�>��\7ʵ������2�A���/����_���S�!xk��b+Luo��U�>W6h�� 
�ol�Mjc��NǱ$!&3��`�T�n��>E0��R�9>t�C�Z��58odF Y�+1�zy�����PB2DmOfW�^��ʀ9�@�'�`��}�2U׏ǯW'����ڂ��%Md�.M�iL'���?C}����B9zXε���O�0�ԷFZ�x�5H�ǰv��*��Z]�&�ب�K���~
�];�V�E�ƅ�;2Hg"!Pc�6$jQn�<���,`�W�!@�)1�l[��KՑ���c"I�X���\�D圫Ʌ�@�\蔯�8C�T��adS3)ݫ����Ф�.j��;_�~61�>�`Gݨh�B��*}F�i��ѷ�W����TUvs�z���Wy"�Z+�D@�\Y��y�>��zy���y2���q��fx4U�i���Xn$�>�[���g��z���:Ճ�����.� ���Ag��+�d�&K�08U"��$����rR0�;�ݺ�Ê��5u�jۣx�^�-��4"���2E����@�p�� 1T�И,pY�3��k�i<�-xw���pk�3���i��g����3]^vY4��+F�jɡ���>I�?;>v#���a�U��da0h� �Q��'V�O&	�6ũN�_q��u��rUb�9��G�tw���P���#��x�)*{���#��<�W�?�R�WGY,�+=�,���9�N�ΐ0�.��0�6�g{<��"�����m�Z����l0>rÝ��cVf}�(نB�9z�����eM�5�\#�.�:�;��:�6�H�<X �AW-�U�휻f>�%���̵ѨK_Q�>έD\���3�>l�pt��~|ڈ�7H��cڀ�uc��qw�NV^��R=�Jd7�4[�'(#�$�\�,��F��ӅDmT�w�M-h_6��:���'�]�w��+�Хk���Hfքi�Հ�Q����ߦ�{1�:�uE�����eж�S˳،=�����Ts�pe�˵� �?/W�{�@d�ǠuC�C�\�RH�@I{7v(pM]yp�N����q�n`��Y7`G����҂�֓��*��N0��ҡq���M,�D<�����u^�IZ���H��6nT�X���@�6��{T����-8 =u�rn��pgi��N��\�5I��)ypK��P�i�\4��.�Y7��tW�_H�6�BAb����y2�+��k��q^��Zǆ�9
���k�0�R$��G�U�A=��9�*e�R��k�ٷk�j�����{o��z�)�W��t[��݀3���8�)蜇-y�z�&��RIz����-�8�X���HcM��:KQI�u�B����3��<��m�����S����:i�ϱ���R�.^�i�f����Ylu�g»�(��ر��;����Н��N���Q2[�)~�i]��M��#�H]58F��������2R�����kI!gi/2*��gn�/kF]Ȱ�"��9�Z���?�Ǔ�_<����I�{��*�!-Oj�.r��9��X��a�ū�*�s�䩃��I�x��IA��x����7M� EJ�_3�-�n�0�u-��(�G�22y�𻾉Jʖ�K_�Y���w;Br��w�zw�_�����֒�[c�?�Js�d ����<1-���c�ߧA�F�\ L����5_�3�ˁ�����������-c��M2�e�{)΄o/��q���\[k�!rs	+�N��T��+ί�����3�Sk��Zɥ}���{�a�Q/��]@���"�Ǻ^������>�m�!�N+�1E��1��#7��+Ԁ�=�p�C$��h��KN��H�u�(�9���9G���L��F�����蔷����иC����fNT!���\\;�Z�y�B&�~�,n�Z�dƀ�0�9;�,��K��>2;Y�Jv�@)F/�t|04�cj?�LUeԛ���,�@�(7��u�x�<e\+�Ti�?O��Kin\�&ݷ<�77��Q9�|�꯵Kk]KUAWZִ��O���8q3q�~��Ύ���)�GfPNd�<uӃ,-���T;��a��ph#��W��}&4#�0h���S���ʹ���^�*����<��� d��	>v\�6jֵ�k1�v�x���N^|���f�Z�ܕ�x�ao��к9��Έ��'����)Gvܩ�@�g�H�%"l�:�@����v�{��,~>�X��%�e�A6�nO��.d��i�c�ʲ��yo�AO$��~�'�nW�|Y.���,�������P���T��|��j��*���g� ,j1�~�e�<�Y�.V�r!�a{5��Q�5\�-�E�k�P��.ŀ��8�2��lB|Ұ=�:�����{���Z�]�5���{%n��Y~OM��ˇ��NP�B]F���&Ƽ��Pi,�������!�lx�<4=�TsY��9��5�o�񑜃*��_�2�j���ҹW�Ѩ�����f��hx|�����lxC�+�M/?.z���hx�+zK�TAC�Z.�����%��\̫ͦ�ފU����ecm�y���{�L�n:G�u�t����0�C{����_
])ŷ%�v�agΊ�/��/�s&�s����~d�,Ҭ��ef����a��S��j_�ǁH��(��W��~1��6�f�r�h����>���6A�`���R�ب��Y�BVw�hݴYg!��P�����A�-�� п��=J�K��&�b����"[�r�����^�/`P��'�V��9�H�Y�Y�=e�x0�zrlì!/��y���[Jl�=Ҭ�f�(�I�;�8Z���"�~=�]yA}�!�TK!���,\y����t<�K>�� OY9M郠�+V�A?}��J�G:�����ډ�U�B�!Ե�J}.��v���>�h)������sKp�Lbp+����M�uH|�uQU�~���5��{L��^�F�� �ӌv��`Ĉ{_���y�N��2���s7���r1#��-�W8�̊����$��~}�a�~��2Y�� o,��#�h[u,����q*�r�nC���_����܏�3�?��,��v���k^�����o���c�}���x�{�����{qvz�'{�ѣp��k?Z��|k.�@��:�ݚ��l��dTUw/��ë*l�o���e��C�O�~&NT�b>�-��
�����F!�{�/@Hhą���H��8.N��tD�1%��y��(��Ļ���j�'�|E(�K�А���:3(�k}����!�U�vS,3�A w�2�}U��lP��6ٙ��Gj""�"x��\���A��U�ܡ�k�콼C��#�B��Y��Se��dU�w���J�S^_�LT�V�&1	#.Opi�#^��u���[s�49��sOgHB�Z���*������b� 6�Ź�Ϛ}��~b&�ԢֵZG	�^�W�E)ౖt�=����hX�Q<sun�m�m,�?��O���JJ�ڦe��5M�� i�m�ڐ���j4�c�W����&�4��������Aي���N��ik�g�V�F�:�p-����wt�~^{L>�����WϽf2��ؤ,�:7�q:��3-�^Y��hGE������*����ћ	˚9vd�� �r�E��g��Ǆ��X孫�\L��d�UCA�&IƲ}1u-Za��Ǭ�_�Cӳ�Gkg�=v7}wK�6Jl ���l$�\�Wy���[o�3x�mc���DHil��	~q��P}���{0���@�O|kǻgiܪ�V��r'�}��Z�v�|:���~�g�_Ȟ���Zl��k��-{~!��{�K�?��tB%�$������dk�W��3��2��k�)$V�*z�W∅&u�I4X�*��U������M�M����l��Ǿ8C9�mה���{>�2�ǲ�%��5u	���X���O�W̽�|^��l���A����)��|E]��3�CGѱ+��JЁ�K��Rf��jX��Xl���s��%��ɀ���O��P�8�tn��VٖF3E����<Ķ;
f%Ok<ݚAo|��1���	������+�NI�M2ډ�.���q�|���c*X�����P"���F�g��K���;�M�ԛ�� ��=ZbQ��r^�;a xts1Г�v�gwS���D�39֙8nS���YC���*E��)���ޞ��{C��j��@@��n�/_��[%�����8l��������nC`�`�[Br�Z��s-1��k�d��a���۷�����O?������׾u+\4M6̮�ԊY�3�۞/�n�r��ޱ.��]���o�|YYY�u1���K1�5����D�.��~V@174=1Z1Z=dr<UO�~ˡÁ�z!&�#�G�H:8v�J���(��۠Ma��Q���,x%�#�A�V6����@.J#�c�{�t�[k#�G�lRd�D{m�3Ӑ��r�"G󁫃��րjDn
y@����4E�j��>m�k�4�P'�A�<����(��Jl�l�t��t>��P@�)r_�{~�5n�� ����,d�ȍ����5~VUaZ�~*��A��U����e8���^������/�R9<yF
DQd��G�_x���Vы�a�C\�1����{�MU�z��Z��9���?��W�����M܆���`�a-lc��u��X�.�
�oo����!��z�5{�l�A���^OKű'=1t��H��_z	��sW�~(�e>��Yޫ� �c{ ���f\�,�*�<d�U_���P���X��U��h$��?�=��%߷�N����<���24 �i�&�Q<�ss��T
�e��ZB�:��W��z��2f��ȳ��P��b�Ai����\�Z�j�1�k����y~5�*..����yqy9,U�NE-.X�E�ܽ3yx�>k�=y��e�W<�&���b���e��>Л͎�W,�~矸M�t��`x��6f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a`�`0��t��`06 f���`� �A7�a�-Y��R"    IEND�B`�PK
     eO�ZN�ɴ<  <  /   images/f4826ebb-d8ab-4c3e-8d6e-ffd2265d28af.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��+  ;�IDATx��i���u�|���[��n-���t����MI���&%v8��b+@N,�����P~����ȑ-S�D���9C�>=�����յ׭��~�=�y�۔lL�8�?��FMUݺ�[�s�s���}���q��S����� '�85�	;NrS����� '�85�	;NrS����� '�85�	;NrS����� '�85�	;NrS����� '�x�A�n��߇�-B��!f��0�0DE��ݝ90���#�B~0D�G0B]��iZ��! �hРC��׃�?<�\S��P����"D*����:��:���������H���� Թ4����n"��"�5�����7��c����"��W����fX6,+S^3Mh���k	�����|=��0&�c�S��a��)C��>�Y-Dv��_� �����
��F���5�G���A=;xX}���^�!�6���n%>��J��/�zOk�wy_�?��9�h�C���O��?{h�E��{�ӼǑ��c����F<X����6iP1�<Gl x]�C>l�H�RX������#���k��_���s=� F:�/���ܧ?�wK�ʧ'�l��5?R���\^��L&�/����U5���)N*�ʰ�_tMgD��#�3��+#��8��[>���t8�tF�Q�F�QG��%ݛ�t͙�����~R���bșxG��".P��(�W�:�i�Qdh��y�v��Ȟ����N'����"�PB׉��T�ӗ�a�yA�;�_�W��0�u�U�n���L�*r8�n�20b(���{�L����G�|�S��O���o�?��n�h:���&�G.�����N�GOIFP��'H�M:=�F�c�g��8嶑*y:�̖K�a�T��}؀��N�y�NQ�TMf���%�i���q��=�.F����	��:!"�vݝm��y������M�$S(�=��;7Q\]´7���\���7n`��g��ob�n�����{{�kW0�1�?���?�WFG��g�h+����8�r�����
wz�Cާ��$M&X����C������������
�G.B����%�^��E#�Asy#��O���1�=�}f��*�|�̐L�ن`�=+�v�F�X°׃Qȡie�/OQLe1<����ak4n��;�P������,�Ri�r���q��G��k��ΐYL#V�M�XY�n:�^*��̢U ��Qf��#FG4����B>���C�R�����b�R���s��G!;q��h�2��a���.�Zy8{G4��/:C�C�Ȭ��B>޼�a/��������X����eI��1=��)]$E��2�� &TCb��q��F�@*����oj��!o��|��$��qPް��S���x����6�8��t:Č��yS���� �g�ar�NG$I��)rF�ȅOo�
(,/`�׎��F��*6�}T�Yx�{;�]:��N�d���/��l��\Ƅ0rB��;�����A�V����EXt��;w�`x>��#��ٓ�4&*9�����ɨ���\z�2�g�I���O��J���pф��v|C�<
��ʦi󛆐�#��p�ͻH��Tz�x���ǫ���h*Y��c$���	���l�h�1"�'0��+J����
�$�ww0奦���A)mt�@D��e���O��|�eq�^�cr�Fpɦ�I6\�ڡ���	aU�G�;`�����&·OO?h5�N%1���Ǩ-t�0Y͡�m"K\
I�3����H�0�Ex-��]]�co���1�����m�������A��~�x�A&<O�gdBw	U=�!��&��G��Ņ'C���򹋈��ڷnar���N"��!�A4�gk��ҫS�(s��MP^��7Y����{���z���|��Ã6鱋K��^��!���YBC����w��yg��,����#��f�J>KX:l�"�5x}~O�I�C"�L�?��L�#�d��{��s�^���j���-]Ĉ9���h�Э*��#�Jr��y1��e���5��Nb<~8�Dn �"�eFN�מy��1��q���_@�7�s0�F9b9���_Ƥ�a��q!�2%eL�C��8�"CVD��E�������F���fhvY��%zW�;�y����|_H���.�
��1���CFb��#/���9��F�ΰ�\AJ�3�̅��|*`��ӻ}dmBU}	��K3b��%b��RSzD8����;p-]^3d�I}Mb�x̜�gVd���P%~a6٭v��O��3K	�(�h��J�0�����������L
{�*�w��{���\�B��9���ҙud��g��2P3�՛�����hc���V�g��D6�a"v������-@1?����-)�LL�PG��Vg�h��N��!<���9z��b���B��qLû��ã=F��~.��M��;����	z�4���բ����	lGMY�b���d`B�2 �-
���d\G�M°�D"�4��^C��X<��W�O��&�3�~8�8��J frE��c<u�����N�p)Qt��kXx�z�PACQF�%B$p9 �tK[;�籷��(I�H�6Ș҄�ь��g=�x�2i��7��4����چ��$���2��-yM�eBU�BR��|FVR,1 ]�y?>U���(��c�h�HA��:��3I*n:ԄѿD8c�K&�"��*�f�$F��³8���C�}�1�!_(��ix�C�T��4���	���~ǃ!�g��Y����������M����rm���%���1��� l�x+����ş�h4P�<5���2�_&����9��ugK��*Z�sp�����=T���|��b�=��e���=�#d�1�&���:��sumG�?t��D�jU���3�]qİ|�n�F~y�@c���/`��m�Ϭ(G8�1D�R�����:�ϓ����_�;����>�J(IP+/`�9Tc�"�UEC������4�N�C�궎yC&��V1!v��Ґ���yQ[=��)Q�jKb"��*ƢH�r�I�:��z����������le��r�a��G4�g>�2���=Ia�h�m��*��12�sĐ�U���j��2�{v� w�G=aJ��b3�gХCTI�#�bt4F���`��k5�	���`�'��A>��dγ]�wo��T�"i��1��`�e����s�,.�4@)h�l�fK͋y�w<;p�g����녺�!�0IϺ-�V3�y�o�2	R����ƈ������.��	?�V*�YZ4"� ��(戯�Ԇ��(y�:Y^�����xR�mzq��(C�G��<B�M�J��f�&̈^(��t�2َF���/ǿKm���	�f��4ŮO�3�}�{�d��@iC��kJr�i���H�������
�w��t��1��XH��	�&r���!�󤐦�6Ԗk(�\
�̂�\�D����DSXЩ�IL�L=.�i�Z�b�W"EEI|x�5�w�!%עΉ�~�|m�ƫ�z��%IS=zx� ]�Bu�B��IC�S�؂���s��D��{�`�p&����� L$it���SP��$��k��4�#�w�TR�5�H��\F�Ign���S�� ��W������dp� �qU{̯$�y���a�ؤ�����ùK��֋/~��뿈��>�ϼw=�=�o�d���>әEiz���>���7a��V�<�����K/�v��!���*.L(���.UR������%E1�!B�=T5=iV� {1���!��m&���&uc�?�s�y[G�44$���ƻ�0�\�������������JX���D��1��)��woR|�02��A�51�;d��9����B��6�kPW�1����߹�D�����!������>]s��a�\�Q{�f��}w��?C�s���q������=�˿��?X�$�YT?�,~��/m���+��a@���uq���Kf����w��y&��e:oH�'��@<�\��w�/jD_#E~/F��ᓮ&j̚H�329��pz��Z0WW��f��ށ�j�'�COۭ.9(#�~���@U]�՟���A�����!���kob��J�:u~M��C4��/�Q�*��m��,qF�nIјN��e�c@���%H��;G���q�a���HA(,ꈟw��;(K9�N�������?1�_���������o|�����?�A7��]�}�ߜ�=_�;� �?G�H�����w���/�q��>,^ؒH���&�g���.�j��7TL�^�o��4a1���_�)�&�D���?8�F֥�x�*�ڮbv�J��:;�x��Kx�������g?��g�Eq���At�hs��2J=��/��*#G�|F���)v���Pz���L���0��yB��E&�"�U�"�=
t	K�*��Ǚ�s����O����SO��2��H�F�w�� �ެ	D�#�
~�+�c
=���-���'3�r�E�h�<�X��ikFS�l!Ǫ�Xt|�<���>�ɧ!��3�;�o~�7�c��*o�0d{
��Ej�1�|砝��G��.(f�T��>s��Q{��O!�XĻ��g#�/��E���K���O�jE��7�����G��,��d���S9�V �ʮM%���g�]A�w@ş��g���W�l��Ŷ��
k�e�[ ��Afd9�����J|�D�����>F-�AG�U�}��P�\�M�	H[�!�Qs�9ap�B���Éd|ry]�|��m���!Y�)���ј	��|P;��r��62�@��ʰ�D�x/�!E1V:��;���^��ͭ-�.^���M<����gq�05��EOu`KH0:�"s#�fRǌ�P���),_�����{�KU�AU�/Ą�1�}�/_~�r��q�3�/~�g��}̓#2�5�X����J���";z�Y��4�EoMRg����I+���DΤ��<����V47HY�q��0���}^��.�|pa�D�T�F��G�
����C*���po��)E�G�S��d�o5���ɀ	>)�<4�䏲�f*�b�\�׿��?�1|j�,�'��p���LVW�=��"s�<K�Hzo�ȥ���xc�CD�!�8:>V�OS��<J��2)d���)����8ɐ0�Fb#�s�h��V�yi4�0s)���%��T$��e�t�^n��C2�0!nX0�fe.d���Aїۥ����-��	U�zJ�-��TC�#A�L��a$I?`��p �1�TI#K-3���������&�M�U@�胙J�;��.��k��P�zט�J������ �X��=w����u�_�x��)泣���d��1���A��u&���k8����ߣX�拘���Տ>�[o]GAꊥ����VOչ�}�̷�|i���r?��)"��Q!�H�-����Z� �y� �BQ�=��)_v!���"�� Ao��Z̈��q�Q�d�)�)���R��#em�����t�r��u��D�z���7mӰY�i�37��l0��p-[M�j�@m���#̪)fF�����(���kҽ��G��	g	T�ϑ^�0}�%&qo�%!�t��l�v��s�aJ1��ƻ�9S%>�*L ֗�4s?�Az#1Bfĕ�KY	���6��sy��%&�	<���X\_Aqm���V�{V_F#��N.�葋sp�L��ή!y�.`�BRځd� �aKPl0���.���a��K(����#�q����n$
=~�~���L�l��w�>n ��p�+`R\�4A9�"my��|5���d/R��M{}�	�/���}4F��$�zh�|�L���>���/9�����o���A|gת%�vU���#?�A���ɔ����J�hu�� V˕<s����)��T�����!L�.����b�^�+v���`1��+��2�w$�\����A"�;S�j_5Ƞ��ˀ$(�d2��w�	㭷���Æv�m�!b�l�~��/���u��y�޾�W�f[��̼�?$��b������0u�LO�	<��C*��^}"���]�WJ�&#�N�\%����;��/���|&#��d�#�GBD�mG4H&W���n���ٿn�~�+��_n��o���{��<��߸����n�VG�ZR���8zǄ�J"��g�}u�&Rdk>��ǐi�����Ņvi��HS��dh�X�x�4?fr��u�'�u��m顋��WI��\��d%:���M5͜z��M�c�oA�����e4��Nɍ�|LX�!��"�F�3�B����%�GU$�U\E)T�I~L,Ցȥ��H�l�g�2gi���
�	�&Q���$�,%mg����^��zv��Ͼ���'ΒQ��XE�Q��;7Q+՘�������K�[��	C���q���ŀz搴�I%�r�����_��p��ҧש��f�ܩ�>VL���ۄ�!s���P�B:��x�v^�N(��%M�TDXr��@&RbZL2"��O��Z�1Ҽ�TR�4:�]f:#H�X��9TW&Y%�M��p��)u:�E Tk���s�OJ�<��#������u)��y�:-��T��Q�K�p}�����?�˿����{I-����ֈ�}���"޸�*u@�堐�ㄛ
�h��
�R��}�!a�&PF	�N����D����g���b	1�Z侸J�>t�d<YB���[8�q.������"��e��ES�F���Q��}1B���8����F{�*����ڙ�$����F<���~,�E�s�3�$���E#��u�n��A��W+Q�."�M���n���iS�:CT�9X��t��5���� rH��C�����I�ӅQN��R�G��$x��EZ�{&�J
f8���F>X�N/8��z| ���߽�ョ轓W���lw���2�EhI/��^W�X�L4�=�~��H�G�d[�o
MC
�"e�	��KD�/���_u60���<�sǎ�����8�0�S��,�D/S�L�)ޛ!s:d[�.y�P�|��O�G/S۬�:a|�rUc��~����Z{��tc�����l=xN]�duS��P�&k_�h�ȼ@�9L؎jv���� � mHQo���AZ�H$�IM)����$fk���k��<�H�6G%Ufd����,����z���;tӾ��	k�DS�Uɗ���R�ej9
1�gU_Iޟj��
�wI�Ұ�D��ʴܫÜG�!s83&�
#6�J�����$.�:}�����#�L����Q�*RHtz���w��tT��ad���G�xM���[�����O��3p�Szj���꛷��#,�L�G�4��/a�D
���^��XRl^S	UbF|L�U��r�RT�HZ�]�M>+!i#M�~��q�$��w붚��P#�#�V���c¤k*��!�9�i�����W���+ƚ���^ ��s#���@&�(/�2�7��0%��.2$%��#�VRX�z[�0�}�NUDvu��Zr��v�[�U�)j4�(��$��jdZ�"�p�(-��c��V����}z�����2Q��e����KLd���������2���"Nؑ��e��JF2e��\i��YҨ���FRџ��*&4T���0P*I��	F��ڗ"�Ӝ��H�����3�Q<�<��y�#��y9��xL�326͝`��3�:�+E��ǯ�����Z�!^�h����Ϩ(��4�|nU�,UTm7����?�A4�s�O�t�2)�xa
�J	�vqkRяU�H�[���#�gW�Y��m��0i�5�	"R+ac���HCK~R�m|zvij�ls$lD�"�ǞB��B�ׁv��g�M#^����=�|=#�A�?�4U��d����gDi�I�P1�Xg���u"��!��#�t�?g���	i,a\����LY�HB�X��v�<<霑�eB�����ǟ�G�����(�i�,������"ewYya4"槩v{�mUê/T�6�"���z�1�KhO�(0��ݱ��S��Y���JˋН>��=U 	�!�ߢ��$���V�ˇ���%|�����Mz�W_��+T�OOgH~���ϛ#$��H$�����%���B�*`^V����R�	�|^���ǪD+I:��+����*�6��vp~i	�W_Q�w��ԭ��4��[G4~���A�ټ~���XL��W�#��b�̫� rsT�"�	�L���=G�K����X]�P!n���x%���vژ!J}�],�p�!q��ȑά�p�FCy/3썻���w�!y��7�n��x��"����x4�'.\Eb�6"&Q�-�<J(1�g0�6�9
ÅɌ�G�Cģ(w�5�9J
���t���(P���|1�4i��C��J��B��L�k��WT��������8�R�~���T	�f�Ҕ��M�/~�!O��n�r4C	��`���F(eh��.��C�)��$JM,S�<Tɡ���^�Uk?� ^jf1���B`����&q�q�܋S��z0��d7)�C��Y v?%����R�PI] )��ii<��l�
�y�`>y&{��)��8(Yn�!C����/��i3�U�DqU�9D�Mj#:�nX�Z�2=,�JS�D �D���
)���\�7-MZ*5SD�AF�`���#U�ђUd�k�2l]j��$/������X)b�0L��Nh�k�{8�K௬�[1L9���jzΘP���J����"�u�+5L��I�^xog�l���� &5�"�W��UT��>������	�C[��x�<�ב�-�y��P��ڜL3��2�&�@	D�#K4I��Tk0�	��]�@Q]�!T����}WU
\�`�gSg�2�L�ћ�WΓ2�|/�Y�(㘊��޻���pUO��)��)j�L�C[&�!T}��D/W�����k�Z�
f����Æ,><�V���%:5��[����N�	�I�0q�V��]-a�T��� �ns@�%�*��.)��,E�$�4#U�L=7�Z�M���Ǭ߇vo5����u���z/Z��VWE��X����t��ӌ^�v6�f}�R�E�� $m��jI�ނB��\�����>��b>�Խv��7
�aߛi�OR'�hw�*!J���dZՈ��9��n��v�G�z�����M<�M�+���]�C���mv�^}�P�h=T�{.6_}K�%h��8��Z�;UK	����j��b^�Md+����%��=�S�����4��zø�&��2�� 7e!zM�u$Ru�x�a��o��љ�`�7�������aŀ"$øF�\>#�j*���6޼Av8�nU��A�3����x1G��Iˈ�%��;��c�����p��g֗Q�7�ѥ�*뤍ӭm����ڠLve��,�U�H�<Tg�09;�|Q���*B<7Tsa�T��,��!t�4(P(N�3L9�5��B��9������.��
�V�0.�x�Ψ\C���~�j��H�sIKMdY�.`@��ҡ4�+K�E`FqG�\E��qQ&&�36�1�h�]Go����#�� 㓎��f>�AT��t2RZ7oÿuW�K�#��R*Y����L�kKT�L�C͍t���-&���^����L�W��.��V!���R��"�5Iz����Ge�}
>�Ռ��5l
�`uM��Z�|Y�5��c4�eѥ�UE\X�Jh	�¢(�+LQ MMM�%�ߪ&Y��l>Kݤ���j1�)�]_SQ�܍&	��P#�Nuu�����������i!rhU�%�ǳ�.���U:� ��a�~ܫ'� y� �G�%�2=[#L]�{3�4�ɻ{R��╬9l2 T������ϥ�Tۿ�s�dC>�s{S�m<F�(̖�H?�(~���]�����) ��'I)����)%��,֡3�MRR��э��>����$�VP�̧������r����f���v�'�ݺ��o!w�t>��,�T��V�#�p|�6�+Yd/\�����C����u�J�&��J�2��#�E9i|0����Vr��U�SE�@av��J��Rd�ΣX4Z=�Q�Q��S���=�����`���<��d��'�aqa����ԄA�/}���K�I��!G�0H|o���piV�01b�y+��� �A��i�a��Zq����M��y�4BYK��u4a��1Y��,��KHs�S�L���m����tߺ��l�Q���<�8D�m�k�1���NC.�`%C<{���eBߘ��$]�S��g��x�Ɗ�>I]����Vr�޺�V9o|�	静��2Z��TY:����0#bw-�'�̡Z.&h.K�f7o���M�8ʆ<���7z�_�BA�^�$���`�!4i����!FB�ϩ��H������4���23��^V�Q��X3U����4������a�Z��B�{wa���o X��������32j��W�١���4�Ut>A)�ɺ��͍Mx�!��]_ì�`��M��&�0cI1���]pl�/}�F�P��/��o}�O�@i��E��������SSaF�R��7HqOX�fᐉ:G��K�����(���ImPyO6�U�OS�#hpd�yN�����Z0��H�����J�T��L�i�ۂކ̑�nF����T)�ϝ�c'���� 6�rF�X���"������:�O?IH9��o}��Od�S?�R��z�\D�~��_W������<&,����P�d�$G��"K��	�dcF�_*S�MԄݔ�[ғ�gn�}ꁑ8��_�X���m�ՕU$S�3�<�����g>����������l܂�;.x�4U�Z�(�X��[$�^�=�I�F��].�{���A�QV#T"N�H�y�����h��J�`>��&�@
y���U��vP�!ͨ1�w��F*G�2���1J��^
5�cɂM��;}�����G.c���e��1��\���L��]B�́�׎�c�da�a���uM�V��E�O@T���+�y�58�w��D�Na������*����5�}�x�>�� �Gm}����#�~�P*��pos�W�>�(��k�q���IW�h�ҥ�NI{%�˶$R�0���]ܤ�'9hE&�z2����j��)��.����Q<Z�P�4�W6f$kƍ
)�p+�%��x��*�~��!��߸��S��"T�d����^]^���>�W�T@��c����k�c�c����W��ω\F�D�@jNG����+t^}�h�����6���>&F�%��.=!���51�|���(N�uX�β��e�HM�������0���G&3���Ts��(��}6p\Y�g�j���rx�g�B�u|RU5-��`�Ɓ�f������g��9�+oj�k8ÑR��Wi��!�|*e~~��Gq���H�F���8��G�`��B�*?b�9�[���Ul�ɷQ^��jU��=,����x�j�պ��L"m���t��=D�P�磧�E�]ե|
Ǉ��X{dr2��jk'���K��4
�c��E
���E�$����u��8�k�'�*Q�ͨ�Rd�I#^&�:U}�S6H��"���=[�W�����D1�t�\���,�����v�X��Vh�4��;��"�|._��Yإb-� 1������n��
�c�ˬ.f�j]I��RLJux���K�jR.���g�����J�������&B(�¢���ۿ�M	��d?�GZ܋�6�QU|]5�MU�{��B`yWT�QU�b�7�DuN�H�׮�帄�E�Y�c����[��GqO����f�/�T�ԆG�){>I����+W�(TK��$I��L�{�MF���K��%H-����)�Ӯj:X^\Pk 3����f�s�7�2R��S/R`3�/�Q��#$I��/Ug~w�8�ɜ��T��T�ly�����˥�Z~⚚,n��$���\^QV���c�H��a���J���F�L&�"n҃Z�ϋ��0me�N�q���?�[ދ?�D��{��`�I�s.�Ii�$�x�#��#��C���$��T�R���*�,NAʺ;I��l&g�xM�TP%Ȟ3@Ph�S�3�	�.u%iבylK���,��/�Pʸ��D�54�8e��Ҕ�;2�c&��t��Y0أ��2q{��YF�(�Q���B���2Pa��juD�<��`F�������e���H�M�*����Q\&��@�qF�EK4��M�9*P�Rd�)s��"i�"��@�D�E���)!�R��}�g������p�U���
�O�)�ʨ�AT��PR^ �7 �ӻdi�,޼��P�2Le�?W��z�H� ��6��`��D��WϮc���zw��z��l�{@�O����Qg�%3A}0V3\��}v��J�/)�x���x0Cz���L��n�ƒ�b
�0���\WMT���F�::���H_��d�2�F�R�tHUOVY'8���1��Y�1�����6f�nR��������%^3E���u��}!)�Q8yp��#DZyd��0R�1%���5��b0�[R��/Y�$Ƅ��wXT�Mb��YT���c�J�@Fd��L��2�4�T]��:R<]����lB��Ȫ%5�Ц�R��5�*䘗�ԓt�"��Ȝ�l�����J^-�+��$ZÙ��A��.�m7�t����$e�rR���V�aȈ�Q.�����e���Tycz��4Z�b1�������=��6YPBHNw�Q�*sg��3|}F�5���7H�7�sڑ,��$dK<*�jKKpi �k��������n�/��!�JY,3��e��D���801�A�)Kՙd7�G��;B�����<>��ۂ�](W�<:FN֕��z�>Vjˌ��� `�^�!>CC%��N�5�cN=ϞYF�q�j1�s���"6�q&}%3ɿ/�-[i��z�"z���$�%�#\ZYÝ�C�IЖH2�P*f1"Q�'���{���r��)&���8��%��㝬���|j����F4��,˴�(�=�-+6�Kq����d<j��0�\��g�^���{���T�]�d��@����2����w6�8���y��}C��P�1���y���/���!��.�T˥�(�tܹ���戄�����j��t��5A�Qqtcm��r}[�l+��+��#�)��9B�NA�ּ���,�����i0��d|%���&�fL=��3+Ut��TU{�V��A�";�����U�G�=S-(j�Du��Q W���V���t�L�	��f"K�cf����4,����7�
��m��ge��o*Ŝi���k�O_6{���]�fc�jU��<�!�{C�	"h5�� ,���U�5��Ř�ՒU��D-\U]����#���d �*��d/���g��o�H����",R^#�B�+�;d�)�d��2�i@AX�f�$���,ߗH%T���PB��(�%I��&�&��8؄V���0R�4/�s� 7q|U��L�����t��Ĝ��й��;}>�4�	NG�ykj����s�Ɠ�*!�^�V�7�/�G��t�D�?"؍��3�T����"�ƥ�}="������
CRm4A�L�<�9���L�R\�=�Κ�Pޞ��1��oRoXjg���{��y�͐/V��tP 5.>f�%b�t䩿�*Et�M%��reYA��4l�%I�,���*����PZ� A��80HE�j��YJ�"�<Y ����'��!§?��WU����/�y�X(���l�4��=��P�g3��.�"�`�Z��1��nS��v$�Z��?��O~��ͷw'��m��Ν�?|�έ[�{����z$�^nXƾ��a�.PeY�P\��3���3�X��<�m�;;�.�/,��������C���=��;�޿B/M2�䘋��j=��dSmr#�)
-���"���� CR�F�O>��7Q��L�>��v�'{�}[��j�w7�J�v�/�E�R���,R�w����ϝ��ΎZQIf�m�1����/�1��w^��T�a=){ժqQ�Vڑ�s�j�Xz�WW����w߸u��/������y�C
c��p���`�)l���zb��*��}���yĺB�d1\����ָ}Ӈ�yG�_Q�3:�����Z����5"cIq +���Zb��ڸ���hCf����������k�l!u��ZU-�09֐�)#��C�xH:�k���Y�M��Nb��P��D�i[u���H�v���HW3���Lv	��������e�Z˲qC���y��z�>)��Z)����~�7�����w������y�yO�$�T�ٍ�r�o�h��0��΄j�����5�Hc�S��H&+�Q=ޏEڪ�i�P���s��>�����0��
2�>YMZ��e���sy�Y�o������'�r5���P���Ŝ����}ǐ4���Bo`FE���=��BV��YE�J�u+!�1%=lG�91T��[5)� ��eٲ�>ОZ��PZ-h~��U�N�M�0Q� �%�te-!�r&�K�"^k�0�*�F}U�b��ƣ���'�g�ׯ��k���x_���B�9�/��"�d�J�H�Re����'�����jT4����-�ąI�+J(��BC��4Eo������4V�R�(=ZG���s���$OQ�`�?���q���XvM6�������v'��ڄX��.;÷,q �\�u=�Nh�%�6q=c%������-{ZG>�?
5ɚ4gdf�*Kˬ.G���ړ�}��o�0����W�x'�0���?r�.?�����@���?��E����/���̴KQǤ8�P�eն�Ö�#��"��T�Q͹�U�ПqT��l�)h�_��Dj^�W��ܯ;��'�g9d/,�JD�͓���U�=�C°L)���W����d�_�������,��&��dy���H�w��k!H&��^���n��t�=Yd����1t�m����E��:^����_y������?��9aǩAN�qj�v���9aǩAN�qj�v���9aǩAN�qj�v���9aǩAN�qj�v���9a��������Tv    IEND�B`�PK
     eO�Zj���� �� /   images/3281a32a-bb08-42cb-a591-9481e2c9eb0d.png�PNG

   IHDR     �   ��"�   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx�\}��U�i���x�b�$g��gq	�����C��lq$!	H�{2��dܥݻߩ���^ _2����[u�����߰qb�$R�4�V��:e~,.7��C��o����L�q����	#�Σ��W�G0�Gw_?L��ʊq�{b��p� �ӏ�s�C(cA6���\t扰�rhh�����N����xN�~K�?r�C�gr��Ќ�+W�dw��u�?����z��n������܎L֊T:�ʀ�W��E��;���y�Rd��L�đ��4�
�k�5;���"c���������i��q{��CF:>��">�v3v��w���.A0�Ӈ�~����#�3i�����ĵ�H�awy���/��_�t�g�8��\�ǃ�KW᧥kO&a�Z��f�q�0fx-f^z	������+��(�y�x�8��ca�����x�d��	��X�N���<�29'~۰+7mF�̯��pﭷ`���r���^G(����O'c<Ǝ��D9s�nt�x�����̳?����\�e3�WI%�i����%>�Mi<x�m���,<��W���a���v����P8��qq�9W��s�bs"�L���BM�GN;S&������X�r�At��p�-py� �s��!���l<��|��ѣ�{�V���È���3��@-�=��G����CQQ>�a1>�n���sIȯ�� ��{OL�2�2V>w�]��u����ݸ�_W��, o�ps�Ű{\�8\\C�D�ꪐ�����=�"l|R�8}*�8x?��f���V�~��33��F�:QY^M[�a��8��x����'���+_�3؃7�y�^̧.}>o9b�hq0Q[�<��<�ݝx����܂��7?�����b�k��Y�<�8���=����<?ÄRʲ��;a�0XW�� ���/�o �.�U���(�i
ך� KeF��7[PR1_��)T��� �YP����щ�_���~�#�#gEgW'ZG��"Ge3[2ȥ�ؾ�;���pv~���@��	����x9�k,�O��Zln��f�y��b<�mݨ��+�KȀ��E�r�N?%F��]=�`l6��(��N"��m݆Dڂ�8y��#7c��fL�����ISeEB�C0;�!�XPZ]��7<[�y~�-N��6d9��wv�P巣��
�7�N�e�qX�50��[����\K�uX���pV�l�t��	"�N �� ��Åɒ�"��p��Y������V*
�k�Z��Յ�Y���6��J#�0�Tv*�)m�8����hV~�h�9�M�a�a�o�P|�|���zb�)�D��=~�H��9��6��O�r]qظ?���N`dm��A<��uP��dx�&�	i�6�s��~Aqq-A=M瓀��D8�F�oüE�1mڝ�>��xa&0�-4��n"ö�Hd�]LY3�ԣ��PRR���.�Ƅ$u(�J��A6;B�4��>��}|��!�|━��I �a�������9$@�pX�� �t��x��]�\3n�*���Z��>��~^4��`\�a�d��L��3s⏵1eʾ(���E��~.!���l�"�O�Acn��BYI)36m�N���s�y;|<���>�z�U���y!��t����4�W�|DA5���J]�e�
ЩA���;���������"Ը<��gf�R��9:�ݣBrҳX�Wlio���@O� b�?�N ��Qn&M���!����G���F57�������lE��A.���߭T�<��B/�I��ts�$�����0�0��7B���r����u�k��#����-"���	(\�m� �T���PQY�,�DE���ٴ�>J3mW[+�E%H%S��f�L�Qc�Nu聈��R�l+A�L��z�{��,�Ž����9Y&��CAt���f�ш��n��j�A��+)�R��,��뷹��rDFz0�5O�0!�ዡ���9�_�W/h�IQ��A�er��5�j��CA�����3mG"ßoF���f(��V2�A�F���,;�$���	4�$z��E啺���nEGgƑ���*���f�R�Y���� �JG%��iD'�����{v$�y�K�̬�-��$�?��,�-�e���YZ�!@@�{�襬�o\��2Iqm6�G����r�G���|��o�e����gE�4*�,z^b�Vꪓ,�M���>יJ[	����Ee���h'&:�b�GD�)o�Dv�E��$(�<FO� /Yj�l���sq:'L���Qd����+�%Mg�$�9\\C��ɉ!:kS�J���}Ɛ�й�ZQA�&��'3,��r\W�rJ�RikV�p]m���6��D���ڀ�u]M-��ǿ�9Tə�<��Y��� J���V���d�Y>ڒ�*������M�L�����A�� J;HQ�!
�a��H���[12�Z�en�(������3�g�a;3IU���r"���sa|�E^�PÝ<q"Z�"4|��	\�1:āS�QD��HN,��<י'��Q�bт�R032�i�jLVD*܋ �C�.��Fb����E�;��(���?���q��b��
c�P�s��hH��
�����0$��P�L/�G��p���hL�6*�x|�	z?�D*�T�@�4��M!'�4�!xI���i(P�T�	�#k����Y�A	=DfQ4��C�@��:jX�U=?���M��&P��aTM���J��yY��,P*Mp��F��?67�C���9���e��ͦ�}Dx��g�$l�L���!��	?��+��a�F�.�*�a2�<1�~ʱ�4�H�(l
V~�	z�l������sm��\���+���6yꎕ:�u#��	+���ǩoee�
��6�߯a��]��2?*|E�L04���<��E���	:-���fS8 k�0�:��:����9d�4t�tQ�6���H9���\�K�	VC�
xЗ�	�����-�0���L����F�f�F6"�'�K'���@���d|6�W̤PDg�e(:�Պo{�~�Z�*�:�R�ښ8�GNǦ���zNV�1S���1���{z���i�N�oV�8*OQ1*��@7õC��"Ip�a�����k2����z�DK"���b"Xyȡ�a8	(�LH=�z?~�br��7L�0��aQ2�?/B�o/�ux�p�wuPA�������nWAجB�8����.���� %����](ƑG����(EO�=�$r�Y]�>���;f�t��.`\N�"�oP	��bTVWb��N8�9�X}f��f���#���:�T�8�-zAz.2OFa"���~�4��OWy9R;�ճ�z����DW^}5~��&R8'���N<��f�=v���W��w���\��S>o�����Ko}ȃ�Ȇ$�]p�Y����&h�KzY*�x����S	:��>���J+&u&`�H��]8��c��\O��KUQtt�V���s�3_�[H��O�3#�x8픓Ѿk+Մ�v��;��d	�9w�@�԰o��n��>�c�����?�D��
F1� =�������D�dn�8��~ ��dm��S&��b��3���I�kǎ��T���=�X���_��٧���+�#�p��-bHGwn��V������A�C��ǔ--Z��jLC��������\�83KwƉ�͘NґFqQF������AQO��6m�ǸQUhmn����<�>C �e�?�%/<��͛0�л�}7m�aU>�����Fȴ�&�;{�tb����H0�E���_�24�&t�vq�6:4�ϯ�_���q�J�7q�y�L<9�u�n�B��.��������	et~Eu#��#�2�Ӥ�+����#w݌xd���
��}:~��l��+A���O�S�Bf�$q�c�����9r�*���0/>��STԌ"M�!Q��|�?\p�H�;�Xllh���{��FBC�'y �w�b~]�Bo�CF�q4i�J\ؼy-^}�Y�v�}ߖsdQWQ�G��V.������i�0� �.+|��xs�{��ҋ��%m<r�}���VS���^dba�~��]�����;|�*z�4�Fcߴi�9�p��0v�h����P�kKaxA�?���(��Yz�M�v�B�c���f}��7|�	�S;��V���x�w45`�5��~�F�x��|�x{�l����HE^~�U�~�������?�ƍ��n�W_�O�	�i��U^���~��G�-Gen�݅��N(���f<��#�斻�N��ϵ��'^��_c����R��������Ex��q���Qk�·�q�5�� �'C�\D`~��ǰ~�r�hRf2�o~��@��Ш����u2�F/���ì��-[�a�N̘~��<�7��������Gh�tR� +�g�D�^��zZw7��g�Ͽ���7)��;
?��,��}����g��{f+����V�='�)qоq��C��_��qN:��|�t��e�t&�w?�0�G�F����o_q1ޘ�>n��lX��=�_|��<�ټcF������� ![5�_u-��gV�H�s&2�o���e�� �������[�q���L3�KoK:ic��8��P{HHސ�x�����m�І�q���ҡ����-@1���Գ�];�!�>��PA��HI8�u��D����S�׾4m^�[�:�r6�D2؏��u�v:�/��!�[sJ�����6�]�uӵ�Q�l���
{�p���ڄ֝;����[/c7��։�?��ԏ�۶ҋ��È����Ӫhy�yno1���+�{�Mh�߉;n��nC}}=ʩܧ�r*�����p��0�w�I� M�k�̟|�-.��\z�����&:{K�D#ݭ߰��G*^���K��&��àa��Ko��M�]�]�p�A���Į�V�M��]��|8>,X���kӜ�i*~�y�5\t�h�r�yӍX���wnǮ�z\;�x)�-�O (ŋ���ʚ�F�@�@����w?/��iRy��}�������Dۮ*&��kTJ9�<)��O.O�3�Ͼ�1q�l�~�=j3i������̊1{���^f��R���{�;p]_͝�Ӧaxu9V/[�7�{��2eK��z�RƳ5�A�|�`!�SFomRoeu�XQ|��w8�S�n�|�s�U>l$ʊ��N���"�TTb�o�a�U�ʕ�_��	�d?o}�	�=�T�3\��'�s�^�w���u�.2��y.:���`	��19%����?�;o�������]��j�{Zvn��o�E9�������ڍ��nxi2[�4�x�=�,�u&c���3�#P~꩗�Ut
�h
���ʆ�0ܢ{�g�KH�]x��Y�񆫱� S[�ž��g�Ѽ�WRs:L2�[��ƌG\ئ�^���eYM���3�v�q��3a���fq�jxLQ4�Z�2�Sow'>�i1_C�O�T�N���r%�w�������X[�ƊS�FH�ݸ����R\}�(����_�E�J9�d�x��qQ6�ɓ��A����-H�Zr���*j��λ�]��X)��$�%�P�g0��xw����B���� ��b@���˅�n��#�#0�������<���ԎF\���1�&^H� �{�<p��XMe+'}?r���0|�j�ī֭ES[�A�
W�o�~�~7��7ߛ���>#�k�;:�J��q��������Ͻ�&=c�kѸ�������N������CFgO=Y��i���v�T�`���o��_�p(�I�lF�q;�eU��q�b�5�b�� �3�W��������EY�-��%A'Yf���n�7l�{�?��������-_��]RR�>��$2Z�bd>�$fwrq ����7 �G]�p(�*���QW�Y���X֦
� �1����ղ��W������BA����T���jw�\��m�.|�`|�5%��K�dRs'��4����wBd�[��S�m�3̒�Ɋ5�PTQ��+��hn(�sO.��W�.���E�J3G2ՋhXM*1n<�ڛ<�bDDw(GQT�%���K�CqU�y�U<r�mh޹�pE�Ś�ih��f2�]��c�*SJ�Yr`�xn�G��P�.C��N��R^d�τ#�G�~^�D�LS�������#�dg��
�����)'���a��������ڎ�d9�5jE�&C)�MqOŔ�7?.���ä�#�K����J9}��|lml�=T"�L�I�)٥����1x��pљ����
��/ri{B��˽7�����D#V�ʉm&@vT�9_��1CC8�!]�:줬�&�㡧^F��qI&�$a�YTY�[�9�fgk?n��\���4���Z�r�]���;��|��v��C�o�� .S�~�捐`�*IK�Y��f�)�t.ɯ-dù��qi�F<l^�u3v���7m���h6\J|�\����y&����~��<�Pѐ�Y�&��6�x��w�z���5����>��$4)��h�/\����GkJ)mJ�L`�w��!�@�uR]o�r_B�����?%����EK�.�>ƈX��j�]֐��ʉ�R�$��\�D�Á��5�b�E{�|��[Ƶ�Uv����*7)���8J�x�/qġ����b")B3�r��b0��C���V!��`����N#vы~D�7z�������B�n�5��o C(S�c�ʙŬuw@IX�r6t�����z��K��i,M�-(*.Q%�Rɥ*��\��K��y&�2~��we�6�3�������s���ErF"�0��&� �$鱙g��c/�َ KkO�,^��r�ϳ�gw�(Ô�����G����ɀ�Fʈ�ת�<�1*b%��T?d͒W�������|�Lz;RY��P���'U^Ҋf��$	/U��.XT��X�M.�3�~�b|=7��I_�A�0B�2��!�&��������	t�:˰����D�d����i�;e�.������De��u��ʨN���/[�KVm"�(&��I���Q.^:Lb��I�#vbA����ѧ��jS�����=d�NX�o�f�Ŝ�f+��N*m�K��P�(��7���L�����׮�gIiv^�XV.*z^bV�0��T�B�L��q����T�"�M+8P��@$F%O�$}I�A�-�ʙ'�ک+֬����H�5���?A���<����?QZY��Q������ǟ���g;����!�oAR�\��EA�U���ʤ��� ��%+��J����sZ)�*H2-БS%�Ӗ
�U�Ǫ������+�e
�/ !	?�ǭ=V�Y��'�u�����(t�+����9#/VTYM�;���⹉\��99UN��ن��.'uu��]�hdd��5R��3�Tc���<�K�UU �g8F��I��-Veo��Y�|I0��i����ɨ�s�m�"��ky]V�c6�����7�-=SQw�Ӣ%x�߭� �ͨޙU��(uŢ�)��Ur
���Y�O[�n~M0 ���Ye~�%�p|�؃��@����w�oK��HZ
��@�=CF�p��� �KSV[ጲ��0lL�Q����j����x�҄e��I��3�m+uè���Y�t���|���N��C�'M;��
��D�ϼ� 0I�A7ٛ�,���&�qQ���E��k7�����k)I(��I6lT�ͺI����"ᆋ�!Yy�S`5ʏ�B�Jb*�R��.�Ac�U;���f����Ũ3�:�'���2��ܜ _��;���<4/�8Xz)�п���/��@j&�{)�Y�\�N�ZőhV>����#��uj�C�����}���HBN�H��/W���r
�)ਚ����j#���Bi,A�� Ȩ��3$�E��:{����F=��*�z��תa��z�$Ȫ f�[���6���n �(�$ĥr!{u�ͩ�v$Z�F�lH�`𦬂����(�i���yp��S��UPA�?)���_�%����U/D[�b"�"�J��f������YM���ѽiQ�̪�V9I?
�]s�]d�oΉ#2�� �v:�X$̳p(�MI���;Tc�O�������2i\�KG.u�4_J��>���H])i�M%�!����	*K��X�p����{���}�-ϳ �.R	����VGb8T�f)�`$y/�n�N�	�,v�����+o�8#���@+�$CO��:� �#��!���C���"|s�Y�b1s

��&1��QX��.��MJ���K���u�OT�gУʢ����B��a(z�Gj�͉��
`a`��C�r����:G���ƺBA-V���pp���R"�7bA��e�i�y���Z�㉧�&�v2Z���`M� �wE�a���3�ҭ��L6ax9�)$n��LB?3�5����a懃}��b�A�&�!
�?�W��O!�j��=����)�'M6�O+
�&S�+��9�O)�*�I_���F���g	�Z��L�h,�`A���oi8��T�l�pf���>i�2��B����:KՃ�ʷc��v�ƇB�-f�[�L}2����n��㥭ږ.�+)�ͩaI� ͆�bݫ��{��h�.�Y
M|z����D/�4V�%�eQIԋ.h����/��Io
�.@]u-�b��X,�MW�3�:F#T7��j2��A]�kkŉGM�p���Q�?��`W�ft�lh�f�U���( �XK� *��&M��@/�K�4d�"h�h#�sgn[I��Ϋm[4,uJ(�s�����~ꟴ'İ�QIkK'��p�6Q������Y��R*�Ԫmj(�����#���ady�8��Ӵ��A��h�"�z�����ݭ�Rz��s� �t҇�����%���̸����Â�K�9���IcN��6��f$�N�����e000��:Obw['��ڍ�Ē/�U�Vv�	�"��X��Ǝ��;S����*ҜO>FG�^�T}�R�?T;/�N腒�Ə������0¹�v�Ο�P[����mf���KȒ2�;/(�}��$��^T���z	�����@cK��/'F`��nY>CCJ<9��q8�J���*CKK�V{�{�0�7Q1l�2Ga\r��[�����Ey���Y?�`�R+{�L`��%��Wc��C�+K��"��]	��(��?�N�Hx�j���D�)�����N_�*;�ic��i�o^�1�����[��`�n'���QZV�O��
�{z4Գ2����9��vh���������0�vӀ�#�3H9J����/�UT���j8abH����8��o�x5m*�<�d�g(��Ҳr�?��a�t^��
�B�H܂���V���~y��t)���գ�����|��1A�M��H�JsTf�`��q�7���F:\�k����8�������~�"�����5M'-*�c��Z�U�z�Ll�}&�;F� ;��P\]��}�=�Ykgə��K�%�Ij�6��ɇ�ӚR{rS���k��كC?����e��^il�j�$BC8餇pӭw��-Q�+J�r؄s���v<������T�t(J�:�)jܒ�ϊ�ќ��H(�"I�i���&��w*����h��S�������=D�h�Rz�5��[3��1ދ��nAwW��2�����+�0y�x|��w|_�H��X��k�DD_*�W^Y��h��c%���pљ��'��;�}�߯�P9���@�����FT�c����B�׮Qd�Q�{q����A��QZ"����A��7m�݂g�z;�"�0ɞ�#AJ+]ȇ�cS��jQ���g�	���J�c�����l<�=�U�+�Ńx���q�������Ϸ��8�ps���p�1���5���)�	������|�wD,�ҹ&�٥睡q��.ӵ
�
9��S�2p�^R����}�q�;��&]�MM�g߹e#�~�	���Hx�ڼ�Ef���X�S�<����@*���Nn�[i�8 3��i'�g7��o�T�&���QGO����0ς *�!��D*���
�i��.��'�3��~e*(��b/9�l���;����h��-�9��776�7_C����C:�DR�)�Rb"�Go��K�������h�F�����k.��k����Ő���^]]��h��o��z�?��D��%wg�:`��Y��u�^H9��O@��I^+�3J�3��G���v<��F�G�h��b���Ԋ��l��؁��m/ϐ�IB,ǿn��?P�1=n�z�-۷���g��gf)�
Ӑ�F16+�g<�=�ߊ��.�p|���BRL�*�|�΃���R)�"����blN�Q鸔�T"z_� ��N���s�p��x�g�-�v(tи/���o��zݨ��,ٌR2�z�tt�����އ�N�]�&P���Т��}6��x��� PJ*�ʡ��~z�s�g���砤ʉ�_� �pQ����	GI��irqq�~M*�$z�v��'�ǃ�?��X/'I��&ո����{nGg�.�y|h����Y��`���������z�X���I#L23$��ÿf^�%P�$#-Ò���<��5��^R�K�)?�/PA��*ݓd[�28|�}q�ԃ��ݡ_{�r7YV%%.$��7^u�}�u�M�R�S�+� .��:t�����xsh��AEe5�����6�=��īo�'�U���������3�?�PO'|
���������y�	b�^y��5!��� ��!���:�p����&h��bt�C�n�@Iy%�N��aJ������'����II˅��e���<�T|<��-aĩ�ø�p$���4ji䪧cK�t��u$8�W�}�mMP®Rl�و�[a􈑘^U��ZoK^~�I�{�ct:9M�.$"C8����פa��m��r=��>tlڅ1#F��g՛�SȆ��W��](+�b2�������9]���\��n�j��8��+�.[	�A<��C�� �%L�A��u4�瞦<[QSY��L���.$��{��4ꡟ����m]�%��#j1��}��ȕ�ﾝ
��D+���ZLh�f">�G�ʫjk�g��j��!��i���MaLU���-fl��U�{���
*������q��*����{`��2���f����ċ�2��1<7���s��MZ~��q,[�E��e7뽕��rz�!\q�9x���
��D���a�}�I��n�p�;�1�b�}�o��RhS��Pw���q����Ͽ��^S�(R	0�B{�a�C��u�T`��F�}(�9q��S���q�*�8��[��Ho���:=�m/��<�����>�[���(&�;`�^N	@=�@D(��H�1¥�Oy�0	�WZ���lܸD�Q��v頯`�o�M�^���z���4dLţ8z�T+򣻣]��!�Ο}� ��,�����3�z"d}����̋��|F�Q.��Y�p�����Ć��X��7m�J�+�=~�2	E��9s��s%f}��6JI���pѹgR��PZ�g(���훰d�H��'�?�d(#���/�C/����`�������eG"�Yk��K/�?���|���$0���ܓ� ������W_��!���n����b���03������BIi�^i���L������3����sR)~$ҏ[���ɝ#	���[z��ST�;[����x�k/Ng.��\���z�?K�Ϥ������ ����/ǂ���\�H1�����f�PW[�SO>l�b$��<�8������,-�Ƌ�~��]�bo ��W�_V����+.`�kV�s�9gk;�T:�\x�?����!�|��/��epT+(���V|��"<��ݴ��6� �@�h�²?V�^zx�ӎn"�Pt�R�<��iT�8��y�O���T�b銵�輳�ȭ�>�e��r%�qur�e��C��ݾ"��旬\��[���l�{��U睅�P��w`��h����5�=x�)|V����o��w���&�p�r='�Ҏ�r����s��۟x�u�%li��ah�nGi�K���(��L���M"8��i���#e���i;��_��K����w�|�&4<�TXa;��q��'h��p*�$��lݩ!�0�1�Fik��o����o���i@߳���~z������v��B/�R��W�SƩp�@9�S9���W50I,�	�ݟ~�+�q�^V6̍�T��Q�W�8p�I3��,ؾ��2��W[W���3O:ڨf�MM�4�!g�&0eF� C�ҊZ,_�	���\��)�W��j�P=9h�	F�^Q�$/B���r��B���K�̫c��+4���l�o<���x��1!H��QG`��HE�J���Va0؇�#����<��pH������U���/q��HG�w/|���i^����Zإz�'�gp��!K
h���щ){N�cϿ���y��I(>v�H���^�G�P��(Hc�u��w��#?���Q� Ue�x��Y����d�R�.�-%`�f52��#��J���H-Y�9���������q�9���x�?�8C�>mw���x�4C���F�
R�˱bS�Y�LY��|���3l�6���z=�>r��p��F2��	0LK3��{V9[>��w0YL&�.��Ly�_%^|u6��հnݶ��v�q>$�a���ኋ�@v0MO�VW��֬F�� Q��/�G�~DG�A?�G�����;z1��O�_O/ً�Аz|OY�&u�U@;�v_8���15ʦv�Sgel�q}��w8�����-?�"���ۭ:㠼���C�c��e+�4�p;m�i�4V޴�A��̼�"Є�o.퀔
��f�k�=4�ˉ������N���ҡX멘{��^���`�&�-)} �ĔR�$���[�3�nk�R�u8Mck�E�c��;i,�����j�FX�($�&q}0EC�w�}���I��.�{He��Q���Ҝ�V����2����~��Dh8%Ux�����I{<^����Q�J#<����u3��7q�bX�"�Z?.\B�nזo�P_?�<�y�����O�ɡS����
%�U��9����J���0n�1��C��ړ��=���7L7>��H���Fe.N`�̾\K_�n��>�,�[|�o+Vb��c��?�#��+���,�ZawR�VpI~�щtu����`���Y�D"���[ޅ!�k���NJ� ~/�CTIý��b��=�pm*�ѼK�C�߲��`J%����Sn3�]v�t�)C;�(m�@ Ji!Ʉ��J*�;��V��X�V��9Ȫ��:���cC�:��G��q�� A�G�؂}��)�VUhk}��='Y��8��?}�\c�ܙ3_���٫�6o�LĄ������\g�Z u�� ��wW�|��eI�����I�I�N9�p�jsy5a�W<�GX�h�b\�[�\H���h��bu��)3:\DҴ��(�$�z��r;v5btM@��c��m�Ɛn��K������Mj��9��Q���ooߌ�G�Ӈ�8䐃�l�Z���:��0d�C�����.�lFeEzLJUh���I(A��g(��[Sx�$���b�ɘ�sW���F�S&���8��Ƀ;2S6�����@O�AX2��$�U�u���
�BO��r�ی�-��q����F#�?I�&��L�S��ոw���WkBM�ANzi	�D�Hy��n��=?Gr򧓟���-A�S�wr��Ɍ��RPA
f鬴���ܓI�R��SXJ�`N_	�].������/׆�࿉�K�1Ig��ؾ�ԇ�Q7r�5�%M�ș�t&a2�"e��T��
K�V�I$̓�&eU�x���R�C�Y*⬆z��܀��;
%�"=KI\�M\i�ƹ��N�+G ���n�j�~���K��GE	Yd�T
��CF�2r�UV�!�z�����SD�qi����D�aF)��(�\�l:M&'�~M#�9��`�YBc3٩o�Ϣ���b�k���Q�H�J��/��.�I��G�A�a'0ɐ�T"���!�W�QJávg���HU����Ґ�&�ePA6��y�qASdZ(!hұ�3(��э��^,��T�	��Ր=����.�����K��2���ҒP��b���ҕ'I&�e�� �)Ԥ%+Mҹ�Go(W�3��8�w�� ���v&Z�!+Sh�2��^����u��Ӫ����n�=;��>�]�l}J���,��c����d�63�r�zY*�16/�٥|l2�-�}��^*� �ej`R~��CS��TfC��q���am}#�j�01*��D����� ��cq���C�֘Tht���k6ʥ�%�� )��Z�e��;:F@��� )�On�r�*a)L:�n���&�si���A:�>-9%���� �t��F'��	���CR����n�V���F�V�+�]�0�������3����( �6�զݶ�e��R�Qf)��?o�K�/�6tu��Og�P	�҅.,�èQ{����]N�Y�hl��������K�T���:	`��$���/�h�Z2R���'dJ��̌)cX˺�L2zN�d)�qqq1=��U�kY\l@ �l�* �::���fe\D�O���tFM#h�Ɍ��=��bd�f�N.����;��e����m�&-� �&�LDz.&���`J(S�=�	�f��/�a҄	�Z�ɾ#:�O���!����'Kr�������,�Y�ۦ՘)���e��)@������
h��GI����x6���J�9�L\��\$�4Sa��X�����ssi���K/p9�p)R�Ѥ�TH��!��"�uD�!�̽&�ç_ϥp�������{���ı��h�f%���q�2�M�	2�B<TmU9����著�)�N#;�ho��q���q�wi��+�̦�?֬�H�����&i����:�^��qw�t�l4%�l�cU�~�&��R�e8�6r׀��+�zy�y�

E���TBf�X�9 VW�!&1�ɩl���z](VJ��U���p|��A�����q\C����n��i%���Qmu%�m�J�`,ӹ�v�O�,#����iS����h�$iB�(�J���v�J��$a���9��\Dv&���ܣC�-1f��Y��E�./Ş�Fi󙰯��aF(��=B����yg��'^�X�zm?�J�y��밻qB�|����}�~���Ӛ��܊��ܓ!��ki��NV��[g^�H�?]�e:�N�lebW7CAi*q�'������[��#�Ѡ�:l�NZ��L�IR���n܌	cGs��1~t:�|�G����/ԇ뮿
���4d.�M;-%���v�>�s�)�v���W�C���E��Ҳ��^�,]�ݼN���(F�S?c*�m� U52�8�>�O\t�'�p,�d�N�η�+o�2�����^ڗ��)�;q����u)�M�\'�|�=2ZӦ��2���
]�;p�ݷ�cw���h�٤=�i������q�(M{���p�Y�z�z�B��d���'�KG�e)�-;v�[Z�t"��3�Ӌ"��A��s�~�]���Gj߄x�H�|�-���{ы��d�ƣ=Ҧ��Ԍ=FTb`��?x���v-muvv�K
Z�0�䓎� A'/M+�2��2NP���^����5���w1<)�a�B=�v>�!ո�uh�Q����i�e�
6ҭ��veʮ��7^w���;�l��s<�p�0���r�ܶ~~v[W�*��O�>0���ظv5���x��9Za�<%�m�q�ݷބ��Vi�w�������'��R�����c����5+q�y�㳯��u2��EeSKZ~��g`צ�6b6��9��G�0aG1�P�ގv\v�y���:zN��\<˦�5���܀�a#�حw�-������������b��_�ٜ�p�]���@�4���<���BGS=c�$c�e�/��6�f}����q�a��av�X�j!�
:�0��+�Ǯ��>QST������:���a��_��OE�r�y�y���7,\��,ӥS����vw����y���[�T)8'�R]W6ol��yp�QDZ���H/�)ĕ_��]�S��	���6��:�%X�bƏ�����}w��_~ŜϿ"h;0Y���܎�]�z�A��4�e�R��i��qm{C#�M��8�D��}9��e����~���=�kI�N�?����T-�QZ	�����}7���-45o�m�^���Ė���H���~v�[G�3��^�%��Ѯ����������+��2���Ӱ�����hnk��݌��O��ŋP����W�'*K���w��btPI�Wo(�o~���JR+q2�0��G��s�<+[���}|�	�E�Z$��8x
vl�c�O�/̂]nij7��q�O<�,��z�jc���ӂ��^��p�=7aż��W�� ��~|b�y i����$e�b��_��Oa������ߗ����j��5�]����oѶq̛ﾏ�.� ]m�������c��Fxh�'�pj�c)0�������I+��&����q֙��G/�'���S1o�2z�|��]r�v���P�r���wQ��~�鹁ީ��9bD5jo�u�5���_t�ı�q���aê�uX���g*��_
���p?=�8��$��Ji����|��g��t��3����e�r2�b<��,�f�JK��ko��fj�TC�r�-�bѯK���>�����V��c	>�~�5Jx w52��d����'�mZ�7ᩇ��U�@��>}:Fו�k�zu|��W��	�O�҅�lߵ��B[6�oGM��C���u�&;p��G�Jo�#�k��^AYu-d	�[�ѳ2�ĜO���k�A�������O;�(��hڲ�l��0��W^�-�э*!������tn�`�3���/8_[���S�A���q�����x��:��8&4���ᵷp٥b��[���=�m�Rhݵ����K.�%�Ոf�{B6���_�O��Uj��0nx%^}��]d	��hmځ�}ɯ��qw�v�˟�fI+jG�ƅ���>t#z�v�+���I�H�'���ж���^��<��t��Xam�5��«�q��7!�{7l~�{�5zu��q'�m�eq��۴G4���p������A6�C!��f.J+j�9��%���@c� ��n>N<f:��ő{��?�?Bۋ�h���72^���w>D���.B�g��i�`��Z<�����b��^Ɖ�6]���'�#7X77u�ǟ������.|FŰ��变1}*)�k�D�D��"� ��[�5\w�G���ϑ�j�E>C���u����oƥ�8������Y�OCOo7�I#�=��k��λ0�i��Tr��b�i��+P�Ͼ������!�R���9V���HZ(W��C�v_7E�r���,Ui-�!:��m�ia��G ��NjzHZ��\�hO�����/���J�CUr�i�F��+o���C�u��i��M�D�s���[W,Em�p���GH�]ZV3��H���Ͼ�=���ձ�����i�Q�Bh�}�浺i�l Ӣ�f��?'嘦�Ƹ���-Ź�����Q�5aҡ�؍��]6lm��K�QQ�ڌ�&�v?����sp�5�!�s�!��2^���$�a���zÇ7*/2�[BH� ����ï~�Y���M�ٽy+��$��E@F���g6��j�|���#���ɳME"��v�Jk�f�8�^���Ǩ5JM�T�|���s�N��Ͼ���/B�,�c�V��Ś ����Lw��W�V���d���%�}�l�2:淿�g�vJ�6�4lG%�����2���s-�/d�r�2b�p;וg�M�j+)������;����\Z�g�G���5��3/��ʚ:7���:n�d�]=����]�a��1�BAY��l}E�(q�=����y��hH��u��H_�0_�G:�%k�P��\t����Vc�!� �ߍHC�N-�0��1�|��O��C�_HZ�d$��"Y<�Cy�h���;���k�E���(#��k��ն6l��EQQ[�x&��2�W����eĊ5���ɨ#r+���.��W�I�Y����v: �p�Q�!s0d�q~�~�+.����;H�%t��w9�g?�չ��DZ����M¼$��ǟ{7�pѐ�ܥ��7�;+k7l�2���1��&;m������3�7����<y��f�
���e���2A�[R^�(hL��-a�0(�b��_~_p��a��P(�7-=dK��H*L
m!���/���/�䴽�/��.��V�8��j㿥t��ڑX��7�X�Vˬy�E�����jI�+K$y���p�5W��j�
"-�`X�ͼy�qni��F��nK��ZA%=����ǅg���F���>���V�~Z���Wk\m�"r��pwG�aq۱��~���]H��5xlh�`��s�G�H�C�D�����HL�����(�,÷������#G"i�y�a�&@Cc3\<Sɓȳuj�����t@�P���=Q�Z�K$n$ӗ4���s6�:_��/�4���q9���}�I���3F�iv��ə-Y�N���#"�z��Ԅ�F�Kq�C���{���Evۅ"�����������X�WFR�)�tQk�sN�8�s�~��y��3kv��V���^���+��k}��T�:��d ��nܤ�RI�kυ[�z����D�K�jº�z���`�07���P4�@y��+pj-�p�X��������<���:$8�����(�s/'"&�F)���ɤ��'R�vx�zUz���X�f;�<f�HW�G@n6�PEdD����C�
s�%��Yq?�+�(e���!�-K	��p�P��ˏ6�k�th�ށr��Ͻ���Kː�X�Pf�����K�L��ǵ���`_)�Y��V���ŖtR��W�a��2�`g�ޢ����vrƀ`�l+�6�+��^����A4�`H2���V}�["gg1�S!��J<��+���(�{��[�q_"�
�M:8��9���u��`�"�l\��'^~C'��=V��.�bq 2._@R�
I�/W��*�dRu.*�s~ZH��W�$=A)��G��+�|���zɮ���?���C��`���H�ڈ,=�N�"��hPv~FV�O�����v��t�ڜ�>5hl����6�I�[rsL�1��L�����^�)\�4�X(�4udg[�^h��*�	����� o�Tp��c�����B����h�ܤ�j�|��L3�����J)()�n�rʈ��Ȕd��65(��1�
�k�󋴡-���睈�VNŮRy��4�5�����&�FBc)�Ke��,�5f���zZF�T�����Zz��;�m��с�*IG��h@�c4��=��&���ieU⑤�譨�nҡ�G#M�øI��Eޘ;��1�y����/?�Hˈ�S���x�2o���S^[��p-ޘ�e$�$�WV�5pO�EH�$�\m��0ʵr=<o�7�rx�E(��$(�ht��~�Ѻ,W�u�[��br��r��Ϲ|����\�> ��gL`�Yc�2!o\���Y�ָߣ�c�P2eܴ�;@��l���K��,��J��c��詤�'�煵��8�LIs1��>�I��TY3�DR�4&/�����r;S����UY
���`Br�A&��eޠ�������O�h��!��ʧS�t8�;�k͊�Me���
���i�^�M+E���{��/��EN&��~b|�sN���.�����:�Ŭ���u��ZNg�?�Fש?^����uvja�xd�&2�6��uF��M'j�A�Ӿ������U�nȘ�\������`�(�W�,��%�h5Y7�M�?.�wH.ˣ���
�?ubEaR��Yfn�e~h�0Ǭ��dV�aMK��bR��&>@�A�P���F���Kf4:��ϯ�VjAތ�>�1#�L!�Xt���c��3��3��xe��D&wI��CF��ut��g�YSƸ$D ��Ò�J�l�d�{���ݘ3j�B��8���99In�J�� �":9�BH5Ȯ�L)��ZF��X���
�B4n���'r�=Vc�K��æ������L�:�?����'��arT� ����9��iͺ���V1�&T0"QT@r�a��y�g���t�ש��~��y>��W��~�_�:Uu�����4.HH(N���*J�]3�l�����HJd"
K�oq����]~�W'��^/C�#rF��f{>Ŋ�ټ��1M�H9f=��hh4�d:�\iC	�}�&�3`���n`���稠G��Ϸ7f�X2ݷ,�ғ+g�%O��ƘIS��t��_gQ��Ü0�x�h"A5�^�*m����i�� ��a���RW�D@��x0��H��b
m[l��5Ϊ�����Qj������V��V.�R��&�OTCx{�C�����0�Lp�������Rhgz�ax$���\��bθ�kڢ۔����^!O�]�-��fō��,A�*�����1��R�)����E��'�|�W�'�Qۤ��99y���2��$!�9�IEa������Q�,O:��P^�������}��y�
E��R&�ZL�UyȘ|���L��c�]��]�`H*���Ő��~��a*8�J&�w`i�1|�/_a��d��:2IC E��RhkiT�7Y~��t� ����<�i�7d-z`z�����hWjq�����qm�Eb:;�����b�_"4�]��Ei�؝�o�7K�=�gQ]S��B���tX�A����{*VB	�4�'���gi��:)���ꍈ|ԣ!�AT/�4�@[ƍ���D�����^�^ޡ��mGcY��jǦ5)�K��؄��|~w4��c<>���OA�K�2��4.��
icc3N�<��Q�����=r^{�m�-��-�������`�ӣ��A������44H�����}r��&%3�gdJ&2�JvA+��f<��}u�)s��}@�~����9�Ll!�E��kȧ�niJ�1`��`�ԓ4<�6�#)�����c��Ү�P�_��Z�ӿ,7]}��_�<*�����o����\���JV4�;e���x����YTȔ4�8�q����b�7�l�8����3���m��x���0��_�>�[�V��c/}�!X�}�)�R�kds4ƍ<y�!7?���l�;��`�p�_A1.��|���*��jK\@OQ{������j5.-nZE��62Q&�r҄18�	�[(),B4��\�e+W�U�T?��`�j�V%��I^|��p�I�a�钍J��V��)���'�K,���aoT����8�9�9/>�4Z��5��x�b�����|� uu:��X����#��[45��;n/.�\,rww Y�\�-il���_}�/O�E���)��UB1�$�3N���G�8��r���J4����̿_��/F����ɄALS�+0��>G��4~�1E.��vѧ��n؂����ʄg��qd9L����z�>]ט/%�%Ɗ0q�qx��WPTZ.�oH�sPɞ9v��b����v�8�FMA9|~����'���>��b��҆����)kЁ��`׷a�%e}����ˉSx�������ҹ/���* �Z��Ё미�u5R��X��C��ً�ϛ���^8܀U�a 8��<�D��,O��a���e����+D��JM
�r��xi�;��j�<$��5�N&��A�1��ш������Ᲊ!�u��p�s]�~��ga'3�I٩�(n��.	�Q��Agg���s�kj��?���뮚�����Vșu��"nBkC=��N%��)-CSr%y'�=�퓰z��/�1zwGfϚ�!����-*Nꎨ\F�ǁ\w6��#�VﯔK���
�x���w׍W�����5�M��V�fyN��=�Tt��ȅ�p�,D���	4��߿�y�}��]
�������!��oF(ԉ����su�������:)/A���p��M�2�C�p�fҨ��R�9�1Megk�XĤ�2�a���Y��>O���K
����P���l1H�]s!*wosVnƸ�N��W��%3O�Ɏ0M�]��S����wuu4㮛��)ڍ��`{W\C�`O�6���d�sg�EKT5*&��a�O�*!�,���W�1��Q_����$���s��Zp�M7�շޕ��W�O/�eON��M�D��c�F[�}����G�▃��%0t� ��t�rF�fC�XC���v��8�{+
|��)G�\�R��nٟ;����9첎s\iK&����+���^��s�ۀ�9��
t�n��4��Ot@�I�Ϭ^��=�c0n�pc�ɧey��X}�X�ʭ�{�l���k��Dy�2�u
�:z�s�GJS ��I1�Yw�\��v\}�X���^]���d�W�ɘ��%�kaO�34�W*F�/�ۍ�RA�����=���PVi:�c��	";u�8L�4NlNPPo/zű57�M\[8"w'���8I��q�v��=H�L���������%!fzd��U�c#gEq9L�F<�؃x���.��݉ެ��q� �'��H�s>n��d����hs`A��]<[�gk��3�wHrr<�i'��i'�Q&hi�1رw?���п���2�@i.'d�hW�/;K�UX3�WǺ�u�\�������0,�)/:���N��N�-iA%���o�й�v���f�{b����ߏ>�d�I h\�)D��t�����0*�շTI*�r��6m��;j�vC.[�
.֦j�A�li��b�Ϝv��p�3�"$ߙ�e#Id"����A��x��7PQ��h�4A�Kf_,�N��8�;A6�RR�0"F�������G��C�>Ֆ2��o�Qe.�ݬU�ˍ��IT�P�\9,�xD�C/�`/�U[�'�Do�SN��$\�:��SA]SKD�E'�'t�is���}���C�`#��SB��g�k�$<�$v�ݴQ���E�7HD��v2~�s�[�4����^j��|�E����4c��-;��㗐�'��a�v�M��_���Ee�CЄ81̜�SB,��Ⱥ.��dsWD�es����Cw܀�_{K��U�KH:u�D�G�y�:֮_���C�I��N��[��m��>O�"U*�$gÝU��n���9y�ؽm~��G99J��r�(�=��7;p��-���"�b��,�؆��v�Vd����a�_���]�b���sg���G��n��o�sv����tu����F#ah
�e���?c�έ:������'c옑�ml��i'�A�Fe�����ttw�s� �.��ù֬[���.�*�q���S�B��Ƀ�߆���M蒻��W��,	+�cI<;�5�ʻ�x�-�1ܬ������Q m�����M��gr�g�NJ$!�m�����)F�7q�┟y�Y�vX_y�S�	��Qw�v�XEN��J\���?���G�����/�Ԍ�����Q+��|^.<g��Rqt��e{g�'Zc&)&�k�R���N?��$�,Z,-*F+�S�g�}��J���8u��)bw
"��s#R�Հ\j�%���8t�^	8%ťȲ���0�e��;n�?�}�Pe�.	����Jj�IJV��?�Z;���e.���ꅿ�������I��C����x^x�:�^Y�C����;8�d7S�ۂ���SN��_��(z�qxC�PAf1�Q1�Խ�����z��lt�p�,�Aͷ\p�|*�E��r�B��;�\�#,kr������RSۑS��TĴ'(�p�̳��˯j��h���W̙#^�U;K��W�A�����ک����?��?ǉ��p����q�jxl9��y�	jh��q3��-��ګ��1D�/;�o&;\�{-��`&^��m�W�����Ç��%�#���'K�}�VtȻ��;zԱ���|%�u�6�OI_T�!7i��K����碭���%���?��erV���5(d�뚭2�q�<+�`f�8O<���C��m�N���Zq,&�v)�K�o%H4ۋQ��>Z��9�i���ư����3�@Z��ȁJ�����{�ӫ�X�����K�i���a�'r��1�S� V��%gL�k2���'�}{UI��BOX�lD�bV}�=��Jq�&��u�+AJUX�K���ҲR�ɻ^y���(�#@�~}���/�'�	e��܂j�v1n�$Ӭ�}p�)�])E�|wm{ }�>��V�C"�߮���3*��JγDu��O�7�Cog���e�1�\�'G3ݬ�P��?�\��P
�M�r�CH���]�F��O9Q�a\.yy>tŌI�(�t������.�7���e��ų�W��(b]�H�D1x@V��,oQqq�*�sΪkVn�ު.44v�LZk�A�.��rT����%�P&��
���-p�l��ExG�ġ���tq|ǯ��=p�%��9�ɠq����]�^���r�)�VZ���Ʀ��q�.8��,?_^R�]{`XE1���ݣ==�z\:L9�8_�Xv��5�^}�-�R�Y���~�X&���&뜔�|M�%�L���(�;�ZŘ�tfnD·T�D� �N-w�`X��NF1��eBa�"6�I����iv���%zY�~Y_^	�X�}��߷��Vj����"A!1���l	)}x�OPY�W�x��nm�ߺk7����<al��B�q�pSCJG7�K8a��b��-�'vA�:Ke߁�8�(���O8g�$%�Ժ�A�����z%IZ=X�lr�+����dT����u�2I�a�}*�s�{0�$G?���;�E��u�\��8a��`
<6�7����Ymc-F3���fqt����>+�\���L��Y�f���0r� �Y�J�K�>
�}Z-��y�U�8v������h�(�
��/�v����%!�"K�	S1�jQ펜<�����C�WR!h̎4:�8˗�����5��+�/�-�ݻD�l�\��G4|���.Î�YB�T�u���ښ6���7��6,^�+fN� �I�W_#	�k�"2I
$���wG�}O�v.�s��U�$;Q+2����k����Y8��~��Gנ����Kkoǥ�NW�j<pUҘ�Ne,���*��/ю,�W�v	��z=f�z"����jS&$���Un��>�Ƶ��H6�u��ĕ��,��U�q��z���|n�]�P���]�p��V�{�Qޔ8�Y�'��6�1P�蒍��üޘ�\y�X����_A"�7O�Nn�n����a�+!�e0A�ܐ���Yݱd2�U5uغc��\$Y)b�jGcK;��������_y_hh֎W&���b${<�~X��)�̨
�uZ(-�괴��*��mʛHjo�W���b !�o�v�:X�"I��1�����+"!f+ g�������Y�Io-��H�VZ�	�{U��G��Ɨ����A�5�Xu�0B�!�@�0˔6rS$�l�Я�@�,���Xz��Jvlҩ�k�);_�;�Ib��䒸r�-��"��6�ܠm�$��^��cQQ���G8d�,�2|�y�*[J%�6�w`��)!)g�8�D�h�y.����f�����YP�G�����W�UX��8s5�K�H�=��P��n���FLU��Zݢ�A��%9$t*#�)���^�İ���9-2q�՚P��U[A�3}X�Rf���f&+�B֌Sy6q�eIs�t���6I\!t�$(NB�!d$$��%��qw����8]l!=	�-�]ͼ��L���*��C�8�8,��������7��6��ꬌ<��d�x֘Zf�ٻ�Y�3I�2��2�Ę|VKg�A���D,�ve�%6�u�t�{�e�2k~q���4�1��0J�p���i�KKj���Z��ӕә2d�G��Β��]����Z$N�Y�Nw���q��RS��q�'A��Y����
��j1
�Z͊�ٓ`V����˨{�Z�g��dr, �?�c�0�*E`N���P�����h�W�J�'[�ru洆t9ٽyy:	�m�Vn��8m�áT5r2`�#�x�l:�5`o�I�0g��C62i�d@���,�	�95�\/Ow}��J;t��ͬ��9�G�1�y�4��̥~�����ĵ�-*��K��{!�Sލ����ܼ|E�&E)���9>��=������`'W%a8&&�m��)�F����r��+$3�ڤIbV����.��d1fژ9�X������1��'F�ߝ�.Wr-\�9֡���I&q;�%N!m��Y��JYQ�D�������:QJ8VM:��'�ǚ=����u�( ����%��T��:5�K&#,��)���]�f۽��v�9��g3�rr�>%�-ѫ���ޓ�[/)[��-vX.nBEL��ON~�����	r�t)�7�V�ʣG�U���cY����mR�ꐋi��TxgFB��V��6�K��3����~�TI%?�3tx2T��\iT�8s�V�bI�����":��Z���J�_��권�wR=�#ˁ|���v	��I���0{t�ҕ�U�|�w�l"/S�,�577����6�,����n��c���se���¸��J?��wg�U��P���nُ~���v�&�t������W��T�%"a��k6��a:w�}%,�� DnE�7����|NqI�z'����=�
�Nŵ4����Y""���^�
1q�KB!�#����u(RJ��r�é��ꛚq��S��oċZ�1֦��	��������jB]��{r�Pŉ�m*L�/�%����Vk"l�Y1f�`�ڵK�>,�`:e�V�mŋ�x�1M�4�j�٩�Q��lX�~���.)+��]�=b�H/,.�߉�?��]�cM,7��)n��SO��g���Na�E�nH���|���D,Yi
��<�-�"�ǃ��9M��)nDt���io9�ݪ��}�I8}�L�d��(2E��s����#��@��r�&�N�Q���u���GG����1�������8�n	������g��.�/d�VBC�@[f�p� ��q
�8��]�����	t���.�{�.KV(�R@y(�l'0vP1
sNv�
рg��#��D�=���a�:�[���ltu�UQ���\�뮿���CbU�x91r�"<����ddIHaL�z
~[��v1\��t�$1k�I�l��Ɖٝ��(�3HM$e0K�ĳ8��	J�EWT� A�	Gf�:	������i��d�/N�$H��Y���t�8l�}P�(�6uY�ĈĂ8��	hm�+�Ӣ̀�d>a�ۉ�lhC��-]8o��b�9��"T���z�P;0��͍��S�H��$5V�e���z3f<�|��IQ4�z�yn9�8�=�dԲ�.�f��e�)��.e���I�ڊ��/�5_�a�r?h���\��zt����Ï{��oFUm�;���|	��
�~�9Ĳ��!�7AY�w�v=���C�����5��1p�g[ŀ�đ8���Q�	7�����o+V�9�r���N��� �d*���+#*��Ƽ�llط#*�(>�G�Ͻ���lA²i#G����NAC����ٳ�l���s�WB�D��1�����w���%�"�	�9��Y֠A�I{W����$L�����n��ǏA��?���W�?�K�]�Y;��gLE��>���ҭ\�Z�)�v�m|��7�玹hk��3�=�"ĵ�aU[��=�6u"&U�P�����lۧa_�$�\�C���=P��ŀ�,\5c2�/�a1:l�lh��7���׋�4�����|��H)NK�׮�I'L@}�n��ޫ%�Z��6�m�B�ׁ�����������Jw�v$)'��v��ȑX&�٥Y��Q�K�}c�l��q�ų�[$qޅ��Ţ��������a�٧��^��`X��Z���#Y@¡�����.����̣�胏P�S(G��=����q�]g��t��p�s�����EE�QG�� _Q��� 6��-��%.�\��O>�C���;v�DoV��rѳ�X�i�u4���G������`D��n��D9@��.�V�[X��,�w���s.�X'��sƙ���{�F�_��&N8c�.F�U���͂\�ri)����;0�����zЧj��ر�F�Y$Ba�O>~voY'���ǟ�+�ë�g��@�^�#��歛�ȣ��e�a�\�d��Kp㵗c���p�7޸e��ˠMf'^��:n��|ڛ�#q���|��gh�/�u�sQSyP�CX�������wd�IsG�m܊~e�8�g3^}�,����F�$0�ܳQW�W�TW�.[)^ӭ�Gd��Q>�t��>�M�s�@�s����R< �rq;ۚ��E� x弆)�$�n�?�9�PZR�x���s3�ڻ�d?rH1���imCia)������p�r��D%�4O����ؿm���NT�yڶf=��&��ea{�Y���ބ+�'H/�eb���U+�T�ۨ�ÔA��Sw�@�1,N*.B�vK,��f�N��sp�"1�WT��^���}H�N�r��*|LEűY��P+�eL���%:���u6P��Z��G�~��N�����\�.�PYuXi��[����=
�܇#S�(�C��'�y�>� nێ9����(�߂����jzB	s�`}�޿�whb�C����%*n�j�.T54#��d�����⽅_�+χ-�;�KOܡI�H��5��vaJ�-�S@�
�r���S.֧_|�;n�6o���&���ٚ����ڰ���5���Я�9�9�ݙ���/�-7^�6ِ��F��gh�!�];Pu� z9Tn݅�� /ϧ�(��۴}��т�q4�݅��E;�r!\� ����ml������-Ԛd���	��`ɏ8m�d>A���E�\z�X�CUUh��Caa	���3x�}����J��_�5n��*�?j.�h:::�uHR@�ž�k4���?S�ce/��에o�"*�,/���``nfb`�5,p�v�6�b�hŮ��Zf;}�d4�9=f| �p�������l�i��Cy��� ��؄`WD�=_~��v�ڝf�=3�W�ۊ�.����[�bL�B�8v��v�]���H7_|Y�66e��6��/��7��+�@ՖM(���!���e�V��f���ㆵ�Ō�鉨�c�j.�o�y3�T1���C�GQ.�.�T�]ɽ�`�3>����"�Ca��a�ԕ[��_�/����$!�ێS����r�V��K��ҫ����H�l�?0���4����j���~��{J79�Z���IA��Y�]��rƜ�!�
�ɴe��Ҿ��}�r�r�^AÜqg���x���h�0[U���j~��TY� ʣ��Io&�s^�8�}�Jw0x��A��e�aK��I��jس���/���F��
���Y�%뒛�Q
o����[v����$a4�ߔP��۟�)���imB2��%�Н[�w����w�{qP.)��@	�Σt���ˊ�/�P��M�)M��.��⍷����CCM5�myh��]x
����<A;.j9:�٦	�3��ڛ��;Q'��+�.�0�m�~	��6'�ܾ́�x�"C}�%�d�R��9��������{�Ś�%���dC��:�oa�Ҡi�MI���"k�!Frɲ_q�%s�+�}�\Rf̙(#I������o� Y#il���UIV���/��&�^��a�;��k���g,�A8��FP^��>�&�>N�H1a^�=��bT=Y��Y�a�JM�q�;k�܌m5�q���9��P�x{�>_�{�3�H���<�%�<�V�ؿ�Z�\��l޲�Y��3�_ޚ�Οq��+3z-�A�p�&7���]M�r����`�!��O���W�`�IF4�i�4���Rr��h>A[o\�Tu8�gcu�md��,�a9�̚�<�9��<��w����X����j�r��$��7Ӝ���*�������q�՗"G>;I��)@^V�8����S��vl����z��l��.�a	�=�l�1�F^Gޟ���z��"Y��:�F>���lr
q���S��³(��Q�ܺ�&	��b��W�~��"B��Xv�d�g1�.�/k��g���<sܮ|��X����Q�p�=�skhՁjoE��5��B?��;�ڼ��9�0���ь�C��Hֆ��Y�F�]62&��f�6����(�?m4'��&���eC���a��0x����sK�/q�\�/���e}��T:��m�C��@���X�շ�� ��P\\(�	�Vn��VH�\�{��r%�+[ ��w�ǀU6��Ï={���xcGZ����tкQ^�	�&����;9P�&M2���G"��CgoS�o�_~�f�m�b�����ń��Ũ�w�����k�_K��ތ�69���j��,�L��~�v�ʃ�0��x�}4�y�z��{�$Lh�J��6Y/NqO"���,=;�����.b�ckwU�����BC!�Ib��L���1��-�������L�w�H�Q�쌡��	������ټ��^���>_ԧ�Y�\��!�v3��"�`��b0ު�hʒy��Ye)��hc�dJ��
��8�މ�fhL=7Z�� Pׄ��KQ�Ӱ*�;5�e�q��"�Q;92Tz��M#?F�$��'��B�y�L�=؆ϻ��3���?icb�ޅ��S�rW���a�o�cɏ��U��,�����$>2O���E��[.�����ID�!��bU���$
�˵���#�{��#�O������b��TM�f�������%J�׳��5�T��8�QV��9H��~�i�����M�����^Y��ۣ��v�*_QҜd2<�&CK�d�f��̶��'e��n�>��������q9��r��2RgЊƑ&`n8[sٕj�C�)�wՆm�v��d+c?�8��Hs��U %�_��`�UM������0��:��Km�xW�"m.2)�V}��`)�R�����NV���	�ϧ�ߦCaR�q� �h��(i邾���{q�!/3�\3c�������]
�Ii�dq�>PO��|cNiZ�(����D����_��%F�Y}9�i;K�,�:�+AR�����I�FG:K��V���ˈ����V��T��"�^A3ނ<�Dĵ�7�迊z��Z8B�5������%����l����m�skW'�6n&�����=�� $�I����n�G�S�f��4֑U��8���iJ��H[T}�茸"Ƌ"N�E�Ҿ^u�RX���q=-rC��r�]�>���[�ҿ���#���,i�1$�]���J�K�L(�����xu��TF{�XCá���Y����1��&�9��:u���cڔBm6D�tV�դw�B��l���q�U����0�2Nj��ș���V��^�1�<i8!���6���3f"Tg���������5,�f���r)��ߥj�-ˢӤt Gβ,��qU���օ�ڥНЖ0O��ʔӢ�x;�,�'?Ŷ��qIRF]<e1�6w����6���8��3��Z�4�ݘr�,)�+Lɸ{�P�Y���v��βPlǪ�_^�%�!`hb2�q^��2��1k�fNۑ����I��l�cC����E��qP�Cv&/�YHu�dw���IչL��a��au��)��H��H�vyj�$ӆZ9)�K0i�Θ�r�a�:g�j3J�)��(7���7�fB�#���j��f��A&�!N(��H6PZ4�Lk��smL��7ВI����g;�܋,%h�U�5���Z�MƺY�I�]�2ĝx�ȯ��#K�ӓ��.�hoDϋ����lj�pƬF���3Y`�>=�2*c&C%uD��b6�y��Oj�v�ku͙u��JF�Bs1&�i�5�HJ�c���pD�^b��1�U����!p�t���i6d����c)H;`I���)h�J�O�ʈ?)����gR���(���Ø-�!B2o��@�dKT<�˪#�b�s��RQJ�u^"�wS�yB�9��j�LbQ9��&l�)�W���3)����DۙQ\�qq�G8D�]���T���X��0%���"਀l�S��|G�%�S�O;�C�z:څ��T�d�17;W� )�c�b�����eߩ?ˋ�CJc�Km
Bf^^�hD��E��Jf����h���HM��*��l��J��$�N;�0�)ei�e���q<�����.�
{$$J�u���ݘeA(�Z�N��l�G�F�q5l�4��A1hZ2��P��K�z�[jй��+Ǣ1�H�&K2�����\�DL5I(���f�I�
�5�Iy�u�&��f\��x�ШS����j:a�sR��F��Y3I���HR��-;�MV��H����9�R�E���pqZ���O4K%
C�cķ\\��?�N��&z�()�Z�Pv#ë�>�*q�����tv�%kPZX؏#������Z`��ް��ٲ`�c�ފ|߮��p���u#;'[�.�I�׭�<^��4��)���6��7�G�����1�d�����������ψ�I��0�j5:l���y����5�<V���0^�����J�ܷ����8E:}�\)5<ié��M��D�h���fLpSyICS��>B@��z�9ӕs�h�����<T]���y9#Ie�D�^NV6����y"r����k�����d��Z����'�\!<գ$psر,иQG��d�U)ZŘ��K�iy�LP^C.>��&U���QwgΙu&J}�
�ک.$߻c�^l۵��5bQuk�f��Wz��,ДI�P^Vj���
��!�b�f-w�g0�M&SRb̬����H�q��+��8d3C�X�8t�_��@�R��[��	C~��O��(�:c��˓���rZ0��5���iȘN����'��H*�Ձϝ��A����Ci�lM�ͷ��/�mȈ��H���#z��tP1��l�
]�،�;w�KPLҤ�w��VeJ��)�L>>ˣw�|�"�ӄ��Չ%���oT�Ui�d�/��QB��e�w���5���Y�
�����o��&AqJ�rvj�*rѩX4�R����B�Rj�t�
Y�:+G.��_z]ŝ,6�����)C@�7"��\��Ga������Pj�p*W��f��/���Q�ޱ��HMe�}RФ�b7� �Z�::ku�1�	��w��Y3q��[���OT�تП�;�n��O?����ac&���q�O=� 6l؊�����mS6�Jҍ�X�CZ9�0j���S���^V�=f���������`1�j�2�,��t:_���Ǟ�7z�ک�Ԋ�U;�o��V|��;X�]̀�"*_�� ��iS�ƛ�?�oS�uʮ�f�;\9�B���7��E^^�\�0���^w��V�8ih��{�`���<v�s�I��z�W�����lyn��T,��Ե����7��XfJ�gw��.�Gb�vH=y��Z�f��8k~�n������jm�1	d�.�y����@q�c�G��^\=�|��B-�Fn�@�I�A�^C��a�����6��r
20X�7]>G���k�aQԚS#��G����������ФY6'f���rT
`��M*J{DRE�T�2��w�uW�Z8�64�V)���#��5���>_��~l�"�� �I��]pŅ��aaɼ�_�����,��6�����=��T�U<�Ȃ*X
Nɺ?�h�7k:Z���5��5YW���\�;o��|i�󋔵kM�ɂ!�т���U�vJ,�Ӥq8�ՃʶF\p�T,[�j���diCV�ڲ�!9�so�NBA���J�d���~E#m͵x����_����N*�[��I��2}�dw�ъ�hB��.N�D��	�y*~�m5��?,̣��st���sJlt��W�/��w�G��hI���NY�����K����#�2��I����片Uq+�&ٳ�D�Z!��~�;z��Z��r��h�p�0��2��x<�M���71F2Z�v�]bd�4��w݂��{U���ҘΆ�hw'~���R+�!��#�d�>��:�lC?*$�atC��H=A?�w4"b�׬� ��@y�IU(
���V��&�D��r�$�%��Y."3�A����}�	���ט�ލj�̲�̼���hm�x��.�)i��d��L���_'�j�U�^�SNJ��JY��`e錽,�(��ZwwE>V3�h�9��o����ӣZ��a�
`�y�^M����C=*��i�Q�I:��k���+)7����h�)a�aLC+J�-��6���T�l`P�'�j�i'NBᾃؾ�F�"S��*1tB��-�p�9g��۶}�r���n��z��ϱ���q��r�6�Z:74��c�����h�� ���ĳ�Q��V��'n��J�{�m����i��f�:>�S;pM�,d��5�qeI�Ѹ_z�+�Du]������[䙇��1����V�$ߙ<�l⌧%\k�-�%ݗ^�'N�4� ��s��=w*����@����4l}�1���������������`��"N:?T��>p��F�=q8<��$!BcS�f�O9i�sk*���=�4���P)��A1��;j�Vj*�aQ�ՍX�����N�����J��l�jE�D�D	1�/��v��8d~Y����R�)Vu�Y���qp%��<��+H�<����<�ȃbI9��ObL�r �{N�r��㨡�$�:	��ܨ�[.1
f	ǈT��>h�K�������W����rnN�x����?�w=�B�6Q�P�CH�g�K���Rp��N¶�[����ϚqJ���0����Ŋ+��-/+Q�}oO+�u�X�v�ޯ�> ��G@ݡ=��V�_��'>�x:~徟v�{�0�\a�U���ގ�?Z(�%Kk��腹Y8���t�yB�Iw�6nU�Vާ��J� a�m�ȥ����
���GBx��G�� Q�'^��]�-N04~��{���Q$�v�x��׋�4�E9�g�r�z��íqL~�U��ԓ�b��x�A�9O<� �}�xr��3�2_�`ʄ�Ps�
%��1��ߵ'dd�bL�2Y�!DCL��#{���K=i�ݯb*���B�;���!	�"=~��}q����M<f�B��E8x/霋�%޺��k$�K��zFe���F��,EK̏{�}�H�)��O����R_��cW.Z�Q���w�w�4�4i� �4PB�(Α��P z�sL-c�� ��g�*�FPM�z��,ÎC59t(��ف����!�t�b��z�n<�ڇ�ER!	��{�A5��b,�e֭ߤ�\9\z�/+q-�p^L��]8���_�(���3�x�e�*�Er��q�Mw!E�9y���G`�k���+/Vuu��z�A���|U1c,�ުIǍ�ȷ�b^���Zk��3r(~��\"!� 9��з@PE�XG�b7��V��Z0`�0<�����p{�:�u�r����rQ���h�Kg�ܼS{����O?U��qT���p�w�q���ǎÇTD9bh��!̜9�7�?Q�eJR�-��$H̝_��������%pz�*o����x���^Y��<�y�eU�����g!�եM����9���<�	����n<���q,�O�����a�D]��U ��bwg3bu��0Q)�l�q�pԈ!�qXu�e���O��L�I[�;�����`���rh��Tt���6t��y5<P�Gc0����4�՛q��>�o�����G�4�,��;.��\|��@�W��#�a����G_���a�4��4r�s�)�g�b`?�X�J_����m�Ǣ��������c�@�xʨ�7�t�+�n��lm�޶iN�z"V�߬2t��S<��{�ۋw�(n����������_w�dI(��؈&N�W���`WX�2a1()�xl�~y���k��&0�$Fz��c��\�R>��n�v5�L��a�l[[����E:��,�=�x}
��_�\P"$�h"������B@�x8;�T�`ѷ?i��s�Y{�<��.3Ђf���eOWn�!�١�)�[!s�-�&h����F��i,_�^	��ܸ������!�R,뻩�"H�!����%�X��
���R%76+�()����n�QB�$�����#���W����a�X}��7�w^�v�2��r/�=z�������
ʑ��,��>�?IJ��y�&l޾K��|Esd����-[��O9YpD.}�x�*��"�
y��:ك������]ҜCRUS����˯c����t���d�R"*(��y&T���o�J�Mq�
oپC���~��^{VA���Mr�,���S�m� +�6:�Iy�o䳊���
	�����ko���n���_M\K�d�2ط�&��¹��Ő!�����Q��1CG(�g��5�#p=�Oc��Ԏ=UX�v��P�.j��d�1��ⳅ��-עGb�o���NA��ٹ����ݒ��U�1����a�4�M16/F��K��I[�ؓ?\��O�tH��8/i�Ͽ��J:?ϫ�:��9��T�X����>I<�\#^��Ҥ������K~��7\�ڡ왡ږ�cUO^����,¶z:p�J/y��������Z1t�J�)).Tfk��ĕCɶ�n�����Y�*Ct^�����f�Q��0W���`�j�-�Z��loC�_����(^ NjyPE�I�>xHø�����1T����̨gk�fL<#����he$�Ԥ2+6{%,rH(1��@�2O� d(f��uu�Q�s)�����סb��ګ�v�p<r�'3ݲ�~��q��ȳ�g��A�O^NVף��E�}���N�L0I�#gc�/�qŅ�$�
�ޥN�GuT's ����	��Z� gQLZ��GH�w�� ��z��u-���܄b	�����R�1C�W�}�5u ���r��n���o��'r�9��]��}��s���ei�0�22�;\]'!�`�D$�MYux���Q5L�i!�A�l�/��r�!��J�՜������AZ����eG�Nj��M�j���l	I�:�4��Z=n�}Y79�5r���p�C֦u����.,)�7?-UiL4�8L��d�����9�B�$�;2
��5��V1�#�<R�͙[,H�K�&c�zdk<e��6���v���)�0�*�j��7��"��F�鉥����	��t���0�9Q�^d��[[Q�-�\ⶔ�&!Y<�x�DO�Z��~C�Ӫ5�VLJ[O�5Ǻ���k����1s�X�8F��N��^��08c"��3���I�IVq^j�=��n�6v`dE씍OIH�c�"I�#���};��¸Řx4y�KFoߓ��[ۆ�����$�P�.t��7�ԲVAY6�OY�J�aa�������i4�r�9�&�d-��8%0���r9,��R�\��\��L\Uߨ��P�U�j�-f�+
0s���}D>��u��|S�'R�m�9L��.F6(�Gg���tE:$���O���^B���]s+�,ִ�'C�f7�s}�-��9�*�э�-�F�P�H���oKѧ$m݂p���lOwhHۛ�քZ��G.W\�8�G�l�NY��cby��R���tK���9*ۋ�r�j�&��v����	ՙ�T������7�P�$��.�L��/��Q�]��$����+���7+@�Q�"9�r��,�CaAQF^�3$gJT��[9�,�[�y��FL�Ix�+	��j�+�O��O��C��I9C.�G���~d�I,n��Y�(+/�Q,g������dZ�361$F���3��,˴�DR�f� /&˗��1YX����S ?Ò9U�<���^�_���t�r��W]�i��-r��i��Ծ�A�ٖ9�iٸ�\xՒ !Fb� �><e7�ZF�9)2�e䩳���MXgN۵��\x�,7�
�n*t>e0R4�jsj�Ϡ�~��ߣ���խ$3&��)B��x�b464����i~�P��iِ# a
�͎l�
��DM"Lήln�+���Qr������{d��r@��{]�S���
�	��J�q�]�	���)�ʥ:�����x�J�%D~�m0s
r�Ag��ѓYV�9���P��B�\Ҹ��`�9iH���5�ݿម�ys�:S%�aR���W�\'��nS}�ʲ��8KWP.�]�}�:��Ì�s�h��Z*���U��b�Y�z�t�*0Q����t�����[�l�����}-{�@��,�� �dmxn8R�)6!F�i3��9c��/�!_�5�+^�LYG���*��e��Ǹ�&N¶�0sz�x�6ٻ�#��zz$M#��j^^~|Vc��������Nr��8O[����P'����Wtj��+(q�� 'M��F9�џ���A^a�l���]ݸ�;������Pr|�b Â���3�����Zu܀�!N�#���$��R	�Jrd�����nS��<��֜J� 0�ɩ�L$f�m!b�?���F���۪�(+��\�#&�ݭ9Ȗ=	�w�Yd����ȧ�>���[^�a�e���������X�Zc��`���`���"Z���Ĥ�1j�:�5%��ԧe.u�byi�G��PT�@-��D,�x�%��8�E���9C������e�Ś]�䒉WJb��-(a���1N���0AC�̘T��.�6���W�!�ć=��6L,�xF���
���R)��9~�'G;
+��@A^�x��\�|-��΍?�h-��MrU�ٻ�8�R���c���m�UȞr��v�Db�G=\.B�&�(��d{"Sg�ODޡ�������M����Nx����'*�LA��N|�d�W˭d�Q0�[�&�ҒbDĻ3e�>�÷�q�0v,��'�/���,�:���G�x�����8�y!J��Ng�Ҩ�[�q[y��F��X�Ғ��3V�B�%��+�j�#��5;��Rc�@qSg�~*���7ݺ���8/�X"�����k��WK�X;���2����&J�JvcBB@6lZ"HT�@���D9���V\r�y�n�o�PGZQ�'�p������ {`B[0��#;��˨�P-�M��U���۟|#!�Wٴ�xH�P!�C�H,�� [2����օ������Ę1������s����Ӌ�瞍�\1X�Z�m�W�:�ɨ�qT��ǏG宭���K����w�˧�tXbx趛��@k@��%rv9�:Gg(�GSGA,�%���[*��	��KB'���X����P\X�]�M�uhD����w���C��������O�UAed�-�������n�@4�\v���\��8m�N�g�g2m(�LW��$Ba�'�AX�N��	�H6����6�ڕ+T4�����n%&i��\���N�u��_P �1k6���R�A���"�:�t��������CoN	5Ə�C�v(/;��ضc;,���Yv�G�b�s�5�	�7��Fc[J��CT�Kw&����w�|#^{��V��"ݸ|΅rPC�RO����rւDrK�9|�p4�a���9�d�*�K�̘�_�}&EI奎���ă�/E%�v����lD6�s�EMm#=Dyi�y�K�p����{��@���W�C�-��\��-E�<:��<v?�Ǔ(�q(A�.�~�)���0[[�yȪj�PZ1Pcl�޷���L?m�x���?�^�S؃�N�8S�S+��=��z!�R�k���8m�	
���Y�{�^�~��-[��N��/=�P���ʺu��)eeI�4�a�6;|�V���V|��|t��c���J�#�p7p`��R�ݘ�G�	M>��<r�mؽ��%e���͢o�B0Q.���q`��[T�ş~���R���UU׌�ݕ8q�͛������Y`��Y�y�Z����bÎ���Ǆ8sXNAx���{'*��������'a��5zV'L<NP��ފP8�������-�3<X]�%K�c����m�����O�/C[{L�Й5�(�ܭ��BAo��kNm0%�:����3�=�8ڛ�p��S���^�v+z��(N�!����H����j�6A�6i马<��6c��#1j� ��/?�!9G}����ET��~�����ހ����x%���BbQP��|���'�;��%�F���c�r�U�?|�&���Oæm���;0��)h:���ƞ<|��smb���ixA!�?׬��6E[�Ǐ᠜�x��7tVŬs���I�i�JM��A�Wu@�B�5Kcw������x����9�tIH��oh��]�@{��{�}���b0�uq�8���Ko���.��{=]5x�����UJ��/�N�3F�����/T�*�٨���
n޺%�$'����t:]T�GEa>v�ڎP(��bźM8P߄��C�W"��<�׋�5�^��}p�UנCP��:9\+Q���2?M��e�n�g�s/)�r�o0��倷c�o?�_O<(��Y�4(9�w�VY��b���z1����g��#<��~Y�%�}�6�i�0�(T��p��q`�A�'��KQ�S�e��I��W�~��~+B54T�U9�a9+��.���e����E���/!R��{����y�\4�9�K
a�pۥ�Q�*s��� :V���v��n�6�9�"O�2gÍ{�x>t��gY�@.:e�8���T���^�G��`?��U��#�)�H��f��@9
�!R{7^4CB�b	C�8XY���=��~\�R�b�N T}O�)�	z��s/��{n��d/{#A��_y]�50��g�����'�EQq-9�c���R
��0�̩wTㄣ�� ,jX�ki�Q�A*w[(l��e2����0-*�-���)�޺�G��o�Xm#�	v��j���nډ���樀�93T�:9��,E��t�Eb��q�9S%��iu5�4�8�� ֪m�0��)b����=��߮r���?�O4H��)��E6�Kb���45F�^9�����w�[#nV�ą_+.S,��א.�:4�LL��/�0k���g~%=~����ك�6jB&(���?��x�Yz�0�r6�����p�M�kY�I�f�!p*���������ͧ_遰X���J�).��?-�ygL�IS��lT]���J�vR���e�`sy�3Igx���ظ�N>Q��U�L�֨ү;�S�E�}��m��oU	?�6v�a�ت����C�N��=��-{�X���gê���o���6�ҙNO	
�r���3ȓ����7���J������_�+k�}%��l��x�b���i	N�<[7lPM����5ʜ��ѯKR�M&n٠�Q宄檼�Ͼ�n��*�����u4�aANEepe�$�ۢ� vO�,���:�C���${�T`�ϋCRvg#�a��%e��.�ҟ?Ei����jژ ���A#�W�č�9,��g#�r�ٚ`G��^S1c~��h��=f�X��q��3�#h�8߇=mZ'b�m� �%˖���Ię�e�p�'A����ǟ�7��>%��zMr�zUP)�0��t��^BQ�
c�.K�6Cݞ���l��D��0�;�	+l�j��`v*y1���A�LV�`Z�	#���Ur�}}�≗���[�*׆�I)tBu�5k6a��oT�3��	k�7�z�	�?Y�%�rnG�R�m��_����(��X�6L�d�WvL�Q���/�D��a�0d����o<�1�$�|���8o�ɚ�hj +ǭ�.7����<Ur+(>�>}ɔUgp�V��ⴓ�G�>�����w��T֛��A6�XKZzaa�^P�5B���?��k/��Π>_��)q�M�����ԼTћ��	ɶ|� L�zrm�Ab7N@�q��Y�ה#F��y�w?�E6�,�ɪ����z8)��{�L�;3�+�# ����(�����g�DcIԘ��Kb�1j�wĂ *E����e{ߙ����>�$��K>FEv�y���s�Q��1{�D>nټ���bhe&IXG
��x(G(��?H�)���Z<��砐jb������y�0턩ڹ!ݟ5g��?�p(����˺*�SyI,V���q���hK�^�c$"yu�2����)��$B*�$�2%���;��˂��+܅�۶I>��)=?�Ȫ�}�p敇@;p46����HC@Ⴒ
���b8 j�X�H��;ҰCR�0��^U��m���֞8?ae�صo?��Q#�rm�~kg���'��Y�b��QCH����$8�V�gJɺ�7>�T�X��Pt�;OK��%�(�8���Y:�E�p��(Ē��WR��?^�	c�k��׈�\�ۏ�uߡ5,鬜c�Xa\�YRd�4��R�����(-*�HϪlw��p�\hjkG�D,ܲu�b<As��'�y�7��ś��.)��ƙM��+b����:�Lb,v�A�͆ 5`x�I9�6�����)uXV��EJ�����g�u�I)����%w�믽-iP��&mJD�p�_�2X\
뫟|�GIn�R�A�gaI������ȧA~�1�2������0a#�@���e���0t�e�m����d.�����Eda�2fS�R�Ei!���J���ޒ5
t�8m7�1�~�}��8#CH,i������4�3|تd(F������'�[���;p3i����5��|��~N�j����N��D�\�/���h�C���u#H�"�i��c�86ٷ�
ʲI��VVZ~�#����VÁ�1!�&X�Q]6�+�`F�"^R(PI.�OR�Z��v��?c��B�)h�/��cю)gV��f-�Z�,'�P{4u共��~\<!��<��P�����=�r`��Պ'f֞��P��Q�F<�:��ˏ��j���,ϰ��{�Z��&�
#\��$�h��� ㈉�4��d��"��yq{�$�g�2Y6.6#��xy'��|o�M�89�4��ܮ|/��h��S����v��,t�T.]W�l5��5k�A5C�٤wq�*��GbJ-�͢�C�Wt�=���Z=��r
Y`��L��A9�Ë��D��a|�[e;�֤!Ea,5 ��ְU�M��A 1YBo���;3���v?%6t�����s�
�1��T�D	�H��ʪ�K&%N�T>m�(�R��j�~�!���0p��*�k0o���z`�r�|i��l>����7 �?�d��ť/EB/^���0�N%洝ʶ-�M�-i-ܙ]�����u�?��횖8��c�p��~��N7���e9���<;���p����s�tW|=�棪��Q�V�%��x%gM+�� 9�~]Jgt�&}���u�����oqO�bєˏ�A�;tnМ��g�s�-Ns��Ý��Z�������J����0�bU���V�^Ze�f��)�gp���m��bh],����K�\?	�I��2y�<H�xG�!FmQv.?�1|��/9�o��zES^�&g�G��)i�І���if�Q>���A����� ��#�+B>�!A1-��9�r�d6�pv?� g|e:=�Ԇ�?�r9T�Qq��l���͏��`��հ�4��0����p"� ERW(����[��9�w�ԝ�<l-'��.�괰@n�e�"Z��G<�"���6e��K%� L��1��nȮ^��)Q��$?���0����":|8�U�KsK��4�z�p3х�g���L��#Z=76��Hq�M:J��G&YeF���o��3�ꆖ�~�<5Y�� [a���@�	%B���d�!�GRɆ�%�rY��lGR��8�qis�Wg6��ğd�\#�5Iw��D�<%1,D��1�4y��3~�bJ+�C�b��gTT'����4]G�Q��\��N|�X(�����%X����%�卶^BF9�</�2+�/;y))(��N܋� ��s�F �sYܖZ�#�DY�jvD�J�H$1��g�Y�L�j~��^@:r_�����LkK��8"�ߔg��%�s��_~�4P��,����#aQ"F���p�B�g�l���<y�I3y#�`�����@^F�<_T�+��.��x#e��OvK7R��J�|�M'L�q↘VJ��##X���4�u㺛�d:&��ӱ����ҘBu;�g�vZ4��y1pc/���N#&�j�GaQ�|�sn��4lb'-��dD4:��Ϊa�ԧ۬Lf�nx��$�m�T�ZSjXN�2'&��B̜q`h�KMf佳E�C\g�h8��`�W����E	��*��^6#�sy�'�>���_������<=�,t��C6��?��?��"J]g�g#����T���|VI0�P��;Hxb���[�,Ť�L"���zr��-�RT�!br��#Z�Oe�yDL���E��.T3ĺTVT"�Պ�#�bˮݰ{|*@:9F>z��)\6G_��3ZE�|Z�`ջ�H���
��慟uh�I�(��-�|���#�y�¤��u+�_�`Ii���HM��Q
���AIc�J*����H�F�yv��W�3	�y����ސ\+f#`a5�Ӆ9�f�N/ɪbm�m��P�HO ޟ@B����1R�~D#!�}Ʃ�rJ6c�|��K���%���+ɳ����H6S%$�)\���sϻ��!�iα oǚu�v�f��J%�i��d�<+cj�aN;d�8��DTŴut��_��7 D��;ЬZ﬊��vuコ����#�􄵍�p/<�s�6�ǒ�_�:�jtC��%�.F!�w7�ر�p��KQD�pv�x�39��湣�x��UqQi�����ɳ�}�(�蝳'�Ҵ�!w�V�ӅK�Le霣���;1դ�����Y�щu�j����������i��+�5��KԱ�w?�P!�<��������X�2%z��r�U�����J*�ɪ����f|��{�"��M��<�w=͸�+�[��),R���^{SuM3��d���[y2%�9f�0�<m*���i=�jU��%K�B}C���ޣ�'��zwzX��̚9ՠ̦�c�7V���p
|�)Jĺj�9U���=ND.�M�_��X����4c���'��!����VN��P�Ks�_�M{K.��l�=�u�������S����׬����4�>p΀�ɢ`�mM8q�$TH�O&nb�zCY��c~��x����	����~���7�I����O?��P���˪2L>a^y��t$Q�ѡ�ˤ�Z5ec�l=�;o]���Úy�ȹ-Zg�4f$�e?7nۭN�j7M��tw���e�\��M'��#������p�-���?�&ܒS3�P�ʜA�K��].J��2̙9]�tXH�85�b��{:0}��(`�{�:�]�RFUޜ�������֛oD��K���*�Z���n;~���Ϣb�@�Ө�I�x��=c�n��&�14Kd˖?V*�fL7�A7���B
�Ęyt
ZSl��X$�I#�q�)�U�,���"I)��+�����=���1�@�4�%E{������t���~q��HX��D�N9f������:�kv����:r���܀A先�7�-�8��[ֲ��]�G�t�m�N�xX���Ţ��,�m��������*�[l�[y�����J�[���C(�����&T1k�T1+a�CC�yN[�%7�a��萿�Mn#�&؊� Sy�[n�
/��>rv�x��*�HƜ�˪J�p��c�jFW(�"��EE��%�����U8��&ʕB�$�q*�P�g��Z�jզYסāU<�֞>�����g���2�(G$����ܐ민L	P�}r �-���������.<����/�Ԩ��|6+�ڲh�;������ B��Ȓ�|�}�]������R���Vƪ^R��k��8e�q�./U�ޖ�.TTU���R�������Z����*4b�FSr��B:��M@T�(���a+����MM��[p�=��cƫ�m���!t�6�r��m�*�αhl��}�B�m$��C?v���ҮXI���O�~����w߾ �p�N���~JK�-�Z���A������QU�"�tbx9�9�Љ�ϝ�D��m=(��Ҵ�,��#����!U�Ȟ0�ފ��.��(��%���ooґ�L�Ee��vt隧$�h��|����މ�F�8��Dd�>o�lI�%��,�X�/Qb���]��#�{�ܫ7��Nq���dĜ����0�٧��s��X��klܸA�x�5עB���z�G���O5�-�u�ii��݋��N����>^�]�(+
���g��:�R��Yx��O�4 �@Wg+�r�8����9�%ؾ�6lP�̈���;�;l��6�$i��.FV.N\"�_^->����R��5K?g��P�ؠ�U�%bP��\RV�V�}N/4 �w����|�E<������و�z8�	�����-,�q��
İ��w�uW��o}$^�%���1�)ǙB�6DuE�zqx�N�n}Ƥ�G���o[�E��,�v�ԂC��/���\B�؇�����8=Y�8n񢭸�����K5̴��ڨx����B.�A:DftB|l�E��Ue��8px�!�{�]x��t����v���`ώm4�Z��@~�q�\�V��8m�<����U�S�h��x���Q�"	��z������+t�Q�2q�>D�p�����e�'�H#��\"�1�G��7K���NO����DEu�kCk�<��#��������Ñnd�=�����R��(X,c�����r�
%��*b��SQV����
L#)[]��"P^����J�Ԫ�����hlm�{/�&1�4L�9[kGMG��{~����2�>�^�z�ǎ��IJ؉��X��J���{0p�v�.�3U;&�5�I���umF�^.B[k��t���� �F����{-�yCV�%9�������"�ٵ/��I<�ؓ�i�����3���cG�����ո�����C�I�8d;N<�X�;{�¾+lN�2�D�ݲGg�L�����Ηu�(��7���h����~�_��Sq��}{ϝ�ş�xZ������}�4�ߎ!#����k��?n5ā���ʹ�˥'w��S�b�n� ��a�5g|b�̲�k�m�S��K��a����?j����נ��֮P}��;�J�2y�0�=�$��i��w�yx�����N�K�7_4�\db����[��F��a�Di]Ī� ��w�,�B�
xq�lD}K��(I8�����vk'k-�Ko/A}}�Z�>���#�YS�U���S��x���(.��|�3���X�Ғj,�v~ؼQ1&*�l5��3fa�ȡr�{qͅ3���_���L���r�/kk�FU������e۳�Q"�x�N9u�J�	c��\��� '���9g�	�X��F>|�n��b͚��1b�hL�r<J�vq�m�������ZM��N<����5��/���
�M��=M�㲹硾�g�2[6?�D+T�?h�F%��j<�қ��A���W����=c���]�z1����9(��x��e:�%Q�~���"��x ����{�~���i����뷉�q"jM!�t(c�\������6m�-�Ƙ�8Ңo���+.�����b�w�=��)9�Nj����h�cgc����e,���9q�п1��+;c:L�����.dű����qvbin���b��%]q�n��$�|�/p�g�H	1�f�����2�~��^ɥ�$�vW��.�Q�E9\i�oQ>������%�;�W.R%�F�˨؞���UC��/�]�Bq@�A�:�>q���R�񣪕d���a����G��A��(OG՘��G�����>�u6��-�s�,Ƹ�O�{�z������E�nGV"&��������FŠrXb!޵�5e�}��iŠ�BP���/Vn��%'��;n��c9�"~����T*����H ���~\�sfO�����*�*�����c�W�AI'Μ!�R�C=��_���9W:gtY�lކի�ko��d�!IرH����^��p�z/���D�2/��*.��_
�����>C]"
�Z���W�U2��$/S]��ZB�t&�m���NlܺS�jH;��`Nr�e߬�qcFk��)!';©<K)��<
m���<\'ZG�D()�<�X��j��E�z�$���'dU�h��Q�h��3"�w���u��������޺]#�sN�f��;\N�l[;����忽�٧h�l�ص�Di�HȄ͛6c��!����Zb�f�J�"ؼe��}}�Fo,6�4���J}��L35E��I����K�w�ۓ:[�)��vP�˰R"R�9R6xX��ẙ9 )G��%��whv�ާ^���]hn鄣����bDM�:��匶)ź�ZC���c������R����M����ч�ӝ�Bg�y X�M'�R����pL	�n?��5�%�������W����ԡ��R(H$�Ө�,�>���;z��Y�9ؿ����S��O:Q��I�LZ>�y!��[��?��=I�%ُXo�hr8.PZ����x�b���ڍ�R�3�_^|%CP����rz{B�1RU��")�QC$up�0�O93��$�8[^xK) 9���a"mC{wX�k6o�c.8_"�>Y?�ѹR�ʸܩ
�6�c�dD���MĪ�ѽ�$���1r�@X�&�6(�b�y�d�J	���QxF[��������mª5�����)��^d�޵���*&�1�(��ϋL�u���r�LN	��q�n%�~ĒI�-��/^�<�ȟ5g%���"0��Ĕ��T��ڲ�	�].�Y.����Ah;w��J�@�hD�G�P٥	J��n�0�<��DYA�l���K�a����NPp��mW[N�R��nI+X��f�P�jb6X�'e+?k�\��权H�CgT'����')yW�4)���v�2(�Pk4gEo�����)k�/ta�#b XP�P�1z�n�Bt2��b���{8r��&�%a���`;4�W#sT%�kj���@��إl�}��ǩJ���P��gt��
�ab��Z��p�,�F6I��r�6oف�F�6[{�� y���j�
uh����¦�>�w��IQ(^��c���<�H��r�ڝv%�ټk���Xe�ZU�f�)> �R�I��)Q&�I�#3j,H��(�i^4e�	hZ��f���[��Tٯ5�5M�Rz(�p�HҦ�!Ma�+>���^y.㙞8�]±%d�:�U��@ޗ-]�K�C5�4֚�l%L�g��>uB|_�ɘ�n�;�s2dC#	8�/ȑ#F�d�?寜�g%�8�V��ДG	�����!���/�/���d�,gr�����@E5�9�9�5)اCe�ތ��]�v�<�@�����Ѫ1��v3
%l���TpGǴ-�H�t�"	+�$���fٌ\�K��jC��J�GȖ�c���q���S�$�����x�K1$Y	�X �3
�?���)���4���Y�X��F7�j�?ȸDak��#�Щki��_����T���mf�*��>�ţ�65 !�!�A�6��H^������N��a1��l�ҁ>��h2�$�;)����&!i�~~2O.d��a�M[�*|��$�����#I��x�2�E$.�cʐ�c�.��Fr{�x$�X��7�^��!0#{$B�[�)9\.��]����ĳ�$��m:���'�=r�rP9����;��[��1�[֜vf�����#fS^F(�#tL-������I�%Qe�,����N��[e?�:L��gדHMӔF�����#�'�3�
�nubH�5P�YF�tfiv3Z@&R�Y�B���d������c����!8;��X`m�:(Shu)]���&`�DW=���������%e%*}��ݭ]8���u�I�BKr��b��J�3�d�Lr���DsN��݋�SO�w�V	�.б ���yd����1c`n�3hRa�e�J�րyW͓��P��x,g�uPiNֶ��G�x���P׷�>
�%�Ѱ:jF�'�4M�-E��S�ј!��޽[¼��8d�����l
��u��{����a��i�u)K��b���hi�'�� =�=�'�OJ����5TWWjxkYZR�d�*�l3�#��D24ZY�"�R�ٱk�^�<i�oXD�w�]r�s����s��O,�������IQ�,|��V�Pr�Q��-�Ɣ�'�˯�꡴X$�K, �=�HIh�S~�"2�3m�Js���芡D�1!���aÑ�k��H+��#ZB��m����s�~UD�G��(��R����㤘V�-�{0l�0��'�=��j�[��QVY����̝�g_~[ۥė������C�*��
g��90ж���ET%Gp1
\^�\4�L+9^?hP�NsN%�2p����[�P�E�uu���݈�|f��%�qț�S^������=uRh�m&C'�3�!0�9j�v��}���u�|�`1���K��\А�e\��D�H���1n�$�/G@�9a�L"	쯾�"Uw��f)U1�{�2d1��ݳ�^2���Pѵt�,�Ǧ@����"�R�(�_�v��o���O�W�� �H��6<����_s���Й�P��!�Hy)&%)�عfn�헸����-*�@�_w�!�w�o�A?����.���)�38��Q$F���.8���c��Ȋ�I3&OFP�3��$eN&2z�h�؆^��g-��0�D|��Z�$����Kl��hcq�ǌ�T��ɋɏ�5T�lb}S�1T�T���}(�M�F%/T�I��G���-��Ͼ���T3#�_y�֨	X�z�Hd)1hVY�T�Os��\�H��'M����d1%4�t�I·�<���w�&�=��.�7�=qz}jn0�0��0$�G��.QBZ��(�C��9瞡Pr�U&����~I���0qĜ�z�L8��ǎ��C-��dM���͖�����HO7�%e���(*R$�a����O,�M����]�?��im�hok����~��[6�hP[wL7��&��ݏy�ߛ$}H���s��¯Vja��B�3�W��;���S`Z��$am�W"���V1�.�:�X�ݴIR1���$l��]����]*)I�#�ˈ�\�a�d�e�{&�}�
?1-~%��ȅ;���qx�nY//vl߮��J��zv�{����X�)�ʪM[e=p��rM��样�SAUeg-�߯�vrߺ{��<��S��曮�{o���K!���z�(��ԓ&���|b$�Ӻ���3�y�N�z�8�k'�^�x��Oi�o�t�Z|�߀P�Drr	�*�;�G�abH���w6�Yp�-z�������!)E�8�J���u�����b&�J8E���K$���8m�����O������X��F^���ąg]�<�-,��g��#�� ��K>ۻ�"�X��=;��wbѲ�ؽ;���G��S���F+����+q��jm��������1��<�{,�r���X+�3s=]	��g�W�����\�Z84_,[�l��{�ᑇ�ƒϿ�7_.U�9M��9�#*�!�u��"lؼ����T'a�N<��ho8�Z!k��T��g�����p�3� ���o��}�SkS�L���OŖ�?H�W.���J�\�I0��I$�z��X9x!L�q"�N:�>���U�>^|�)l[�zN�z��lD���d�Pb�$���e8k�Ltv��_݀�[b��KH=��_�H��Mk�k��7������x5������Xp��ȈQ������ɋm��k�ͷ\�hc�b$���k�>8K44���65@>Ijw����xo|�	֯ۀ1�5/>�8�wƌ���$K��7O8��	?7lچ�ۊ22��<x�/��_@�v�<e����p� 
%�{��W���+�%&�Ǟx��q�J9L7W̿�v�Q������g�	�_R�/���k'H���o����?�k�aȠ!�ͯ��K���<'����?c6�/zWR�F5��KB�^\.�_LK/��OD��`ǎ��/�kkw�"�a����5+�3`��7�BQU)���#݁�������w�D��3�狖�Q;}�t�۶A��v*�⥗^R'�e��K��=x����d����܈��}���q�r�>m�/�r9��v�)�O|_4cBa�0����x���	�i���#�j�*XT"�s�b�|���x��Q5p�F_������.I���2~B��;k2n��j=;��N4<dP��g��9����Z�(.+�#�>��=�4��h��NR�cΐԍq,�XX5a�eX�a3l�4I�C	O����o���|�,�]�cj��8�Ș��xPk�F���b,��V�WT�;��B:J���]���M�0yT.=�qI�b8T[���נj� T�/fNƼ�OEw����S�E��!�X��`��($% ��T}ۂ��,\�����a�<�ۛ����k�6���	o�
i[������(�YZY�g��&������|��߮�˭X��K��A���X��ke���/�S��O���߮ڂ����ڄBIM�x��o��[\Wy��_��hJU�
K*ݝG���.�o���v�øp�#����������J��.�a����(E��ԑ���ɻ}�~y-�=�ض�;SZ�y�ގ��Q�k��34u%�ޢe(/���ǚRԜم-���8���F!%޸���q����OS̎��PX5O>�2�%5�hM��� � �W>\��f�*���XӇnI�w�U��v��q3"��y�Or�0�sJ����ʹ�b��oQ]^��dOXK"��o>׶𪍵����v����%���'n�w[w�A�%�_�Ʈ��Uw�qLR��?�Eb�r���Cgt\�,�7����v�`Ň  ��h��Ok4��z�Ӆ��%:w⠠�)i�2�",Y�	�D1���z�RI#z$�������s�v�Y�A��΂u~l�fb���#��Ko��Ii�j7oR�a��-:��_��[���oP>h�1�Is�19<�,��m;��������\�O,;��q1r�1�NXt��57���T�Ϣd�0�q���(Ö��e$��D<N��n��K�ǞTF�F]�c����P?&��N����c���E�H
l�(�!w��GGP�R<�Û�HB�X�'Ń�⁇���O?���Мݭq�-|H��G����=�M
lٴy+
��%�M`{�^�ܵ����>ߪ���rk�hŢ/�Ĝ3f��F8��Ӧ��$?	K�������׍a#�'�`i-�T�ں��Q��
����y�x罏To��Ѧ�x���V6��������u���qV���je�ZZ�ڎU��y�G���_yW_}%�H���S�mZ$�(--��"���0�uv
���)y剪�+����B�*r&��ؿ���3�#�����#Ym��M��Y��ߩẺ:����p�'����ۻt�"΢��O?�/-
�O��?8�.,r����ӧ!�(���Ĝ��(lرF;�'ԁ�|M$�Ӿ�S��K�����չ��GZ�~��Յ�b?ꚱw�A�#�#k~�'4�ۋ�ڜ|�D���+�� ݟx��?o���w����P�7|+<
좰nUYS��/�9��ɔ�B�������>��>:)�?���+�c�.E��v�)!���H*{_"�����-;d�0�^F����U 9�˯���.8��=�}�v��.445b鲕(���r]$�&=�%���=Y�Ï�t�xL;a�*���]{���{�X���56�����?|��F0d0^z�u\w�E��
����������ŗ��Ҋ
�W�XW�����$][��f�I�z�P�D6��u!�܊ϗ|���O��o���с7e�!ՁD����^\v�\��[Q"�I'h_݆߭���c�o�K�Uyk/V��Il���%3F���"a�޺zԿ)!�����>��T��]�mI�Ɨ⌙����&�(Ʌ->,��[����EkniĖ�_ig���T� NQ��1䴏o���k�x:��d�[r�A,4Q�]=a���oT���v��?�����#�KW�R�mm߫����Ҕ,��<��x٪�3<�	>[�-܄}�汚�K)1�$�a��u�âB&EW�n:�J^�?ˡ���O�C@� �U�0�����_����(��d���d���㳲mi��0���1mL�%�<Ex�aqM���T#���P"3��&����R˖ED��t�E�D�l����u	�����W�v.�S���eF;Q��tH����UZ��lM@�vm��������o4�eZ�y��m��PFwNeӣ�$|�I(�3Jew-��T�����3k�ʽ�H����}}��N��_>�-��AJ֬<^��P�g�kh�ԏƊ�[����R�f���4G�]�F�_:�=A}1�o��j��y-&k�#Ƈ@I����(�0m���4C��doZ:�x��OĪ5��ma�>s6H-sIՂU��\F�ſ�QIu>S�|�Ӥ��ΏW��[�^1�7ʋ���JGaeQ8�e�X��`�e�ֱh�c�����tjW���U�K��`N�mSZ�z���O7�� xLذ��I��083l�B�8Vᕞ.?�3�%�e�,V&��`����e7)B������^�߲Ӑp#㲩��R�TA��,�+��X	IHA�qq�N�z��
ꐵ�U7%R)��&8��A��@�a lY�>��w�]�d��@rZ�����#�S��ޤ\(c����D^0Xq��LfN�6AI���6��PK���!AF��*ؔ1Ɯ-]_�C8;CT�+��`d$�N&�����sd�F1��hReRVyIB�$���Y�Y�� �2f) DHS��g'�b]�8��p���� pɿs��'.�%uO2��:���hҎZ:k�2bNzR*aɝ�^ïW�d���pjN//Q"O�䔴�F�4X��J	}m��=�;A�u�(1�A����$ɗr&�7 N(XZ�sD�]B���u&�P�@?�C?��Q#H�8Y?�U�̥�)�H{ҢR�^��( ��󯐐J�G��0ރ�`�S/�R;���G.~��/��4��UΓ��4��+̤��j��j��'!���eӃ�Ōʥ�x9�5F����ݔ�E�I��H��j�/�ae�\d��?��v�1՘'���L��F3Ҳ�y!8�OC���'�BeH�M$����	��Y������*3VF;5��5¨Ԟ7|�F�����h8�3X���/Q4�P#�&�ُ2Y��)�1�T�(K��<!�ri�r���`j��"g�!:��qG�?b&��u;�D�O�,K~�m�kY}&�N)�*Ő�4�����f#/��gԘ�w f�DDcK�>��nӴ�5$��ږ�ᯠ��Y�<ˆA$��<��DP�3F��L�����l��!"X�]���(C�rj\-y"���>�X���ESVs
�gtz��1��g�9�ݟ�j��(� ���h���f�l����Y��X�"@������b���A�+��#�����_��fP5�sG�����f��p��<o�_���RDRsHS�!J?���ܨ&��辊1�8�11*���p�+�7ќ�@EI�HL� S2�팴Fɍ��O�<�C�]��vBy�@ �hN�9ְ��.�$3��"�H�O��.��P~�i����%傑Xь9�V�*�K��L)MZqΩ�7x9�A�M*w�b����{�I��մD��:}��S����`�D4���nW�>�&Ǆ�BI����Z��MQ� ǜT*?���cz����S��`/S��W�=GiѱjZ��v��,k�P�V>_�׈�Rj���X4*�G���]��� ��o�vv����$ �hOI�K�G~���� �}�L���Y.`:e\|�~��9-�-���}�(//3�ih�G>���r	��k��5��p�h ?/���A�X5X�)�ŉ��k��t�L��t�u-n���nuX����"w&S2vG�q�+*�2Љ�t���Q�^�,b=��yʅ���(�7އ5k7]#���2���sU͍��q҉�{]z^�%$g�M枽��.)�H'N�i$McA�Etkwgj*+p�g��ڴej�R �m��h��o����(.9��O���#��a����� %�՚Ndr��90�G�&~��sf��cǎ�5�:�zH �ҫ��1"Y4�WRZ���s
�Ů��E��.,�v�"'�D��:"q��	�-Y�W�C�0�C�f���$���_�g(8z�����BJ�����3g`��pZ���G��%�Vb�m�4X>;k�W�ܜ0i�{�ܱCbډ���T+k1;T�8"���-TY: �!��آ�!=�����m7!KꅏDz��gQU= Ͽ��d��_D�ߴXO+���r��'y�]),�QVQ��?�Î=��#g�v=Hq)t��@[s~5�
��
���"#פ��v٨7(/W��e�y��C��/�������Uo��7�D.�c��~9(�d&�j:�xq�8!��̙s�g�N��>|���*+�j�F�۹_9-�+ק�����Aq��gjg�������f�4Ͽ���x�,Y0X��#���9����REp��6u"$�!�ū�(iG!z%}����U"��)�bG��)ǩ�!��E��ҦK/<O���������?��w߁���(�0VJ���#�Ř2�8��A���r&�h� �!AOW;��Vy�B�r'X�L�Ӕ�b�~���E�NT�F�F�$���c1�iH���t#�P3��Ϟ#��+�EQ�!����蝿��G�����|
��zymqy5<J�o�<����Gծ������:�Gn*�xͥ7|��47�f���vܹ����c��Y���ڔ�O��Q�#7��n����L�[�h7���_�m�8�I�8@����!��-�4���D:ԍ眊���LG�sy�;�~�4�M��qռ�őO��N;@b[��&����@sG��^�Uq����%EuY 'O���z�e苳6��ה�t��o���>�
)
y*�ln��d�����u7�G��I��ٔ\L��]�j>�k����B�|�ߋ��Q�� \GK��
�u����J����&�Zq�)P#�>�ƦV-8�R�<@M�!{)Y�s��P��H�G�'7��
��:��������3��pl_���Z�b`��衃�p2���6]#�<�ʦ?���q��CA�R�,�d�"ϣ�)��
�iL�4R��>�K�ǎ���mM�;x �%^�}b��Y���Y�]x�H��{~�`QY��(a�̈́���z<�� i10A�(��`�}�x֢I�$��<90x%Y+E�7]u9�x�5���R�gvGV5O�r�%"�4a�[�%=���?����eC��0������{�z� �?k3R�\2�������l��u�����)C���D{G;~u�\���W%���:�vd�ψ����q��qDAsCF�U����u��*�3�4�+瞍�߭����S���ttBN�\�̙y��m2.��z��JUԙ�g�4	��~"�x�E��S$nNj��Cmu���?A��	>�C�	�p��
u�*�e8��g��ڋ����D�=�	%*�JJ4�p�_|:�N�ֆ�g+�����[� �Do�]H��x��?�;�E�Y���1~�=�řyā�����@��'{�	܄R�:0v�h�W'ʊ�� JR�E>�ah�xN�u½}��ګ��[��f�d�ȃJO��U�l^�����>��[�+J�.��SNR����N� �#�b�K��y睇��Ò~��m��#�"&�%y uZ/<�l,����Sǁ>���	��[o�Ӥ[��L.NRޥG�IR��B�͸p�,]�Va���2jHK�G�ނ_]+���/X��pTCsrK����	f��0m�d�۰	{7+�=#��!�݉Y'M�p�R������(����*T�����
/��F`�DZӄ��9��Sz�7���@g?v�܍B���%����;��~{'^{�cĨ�(Ǝ\L勉r�E砷�.O��?ٵ�ho��VeB����N1~��þ�f�� ��B��=CL����rH��Kp��^[���2
���w���>R�Z%�>s:J��-�L������p�:}6��եA����.�F�����bEŘ1s��~�7��o��;�*�$*�����;1�)X�~���^�5�$E���v]V+�n�n�وG�8a��P�����}���E�٥@��Օ�.�.~���hlm���TY��ǌ����O��5�,2���bPu!.:�j�<�㏟�[��(�Z���D�g̚�ӦMA��x�޻��g���Pg��t��J������%g�+Fɋ9���b4N>i�v�
$]�����ُ�?�
i�I����fa�1��+)�܅?��)�n8�eʀ~�%���C���s���ܪ�"cH���v<�����f(v6����_�l�aQ"^G���k����ݻ�e�b�1l��"�2a��&\v���z台�ܕ���:n�NrXk��}ظi���ղPg�q��KiY�93N��Uk��REx��.�W_y9�[��Vaђ�X�a�Vo��:i�w��T�1���ر{�
�	���x^<^֨��ڿߑH�[������䒳$zr�s�1�����?�I�C1���%��wie�ϰw�A�{�%R�w���#`���c'(��'��;;/�?	��K�cY��������h�T�+¤qc1t@��&��p�E೥�4������n�ıƳ%�|�*���x�Z�'���K/�a�����g��w>��@�ȳ��]|�9�joG1�$%�۾s'�n�YאNF�ƀ�
�/����%)1&Mf�Q7)m\F\c[>z�u%��K��B!�6��QIE���r���"8�E*�<q�1(,p!NR�a�1���P�@������=�rL�ȁ��)���3�7�  � ��^�w��mYÊKN�qם�k�u���"lٵ��bT�6Z::��Ã���I�<~2:��$���P���<,�+���3���K�������w�q~{��rK��/?h`���%2��?+*-(,���
�aُ�#��]Bw�i��>��,DK�"��AP���u&f�y�bl)�~��["�,��;�o�W�`���N��_� ��@�e��a����I�R:r,n��v4�6���`��W��E�,U3�(���F�ݏj�{��Z��W<�#���K"���O�y�5�
w�\"�W��>n��;�������x��ϴ�H��n�]��.2~�o|�
,�0^X��GK����c$��>��[�MN�����U���p��p��$�2H�LZ�7ˇ#9SGK�����o~���k&q����]�x��$7l��;�1b�/�Q,�[ÿi���g9�U���l�O�w��7������l�
�=Bg@H?8y�x�[�A�p��2_ˉ�b��_X����otuF$�*|��%����*���pP����C��7�����#��)�u�G���42��U����_|��~1M65!��'�8�.\�-@��e�r(�Z��h�X�u�v��l���ҶW\x��@B椄��zP6�!=g��n��i�o�-FN��"��w��$�y��(%,�F�����O�A*|�B���^3?\���=*��+ٰ��"�{����1��?jσ��a��,Ƨ�7���r<���
�&j�b�)1�K����93�I8��Yg�8��Q��v���������6s&�����^�ߴǎ�X����<�	ͽn�|N�qfξ5r���9(��K΢�+o���.�Dg~���;��f����ͧ���*&�k��c����+�?S��rLsS�8�Lv��,���JTkd�)٠C��Z��^���ZS&ߙ�񆞖�vve���+�ߞ~�R�,y��\D�x��>�\��>�g�:C=^m<P��H	5��{���G��ze��(��f���D@ӎ?V	�(�X����$(�j6&�I;���'?[.w��nI��o����b ~޾SO����V�;9qR*I�1�V:o>�b���BNI����w����K���)ah�d�n�A��'���;n�V'CgN!���v+��K)r�S�Psr6��Sf���C}��5�4�F.���P/��&X(��$�I6�+)���{�09�>e�{3��;�����4�u�s���"�v�jFKW��27�ġ$l*�S���뼈���T\W}���]���nڻWR�$RV����l�������I��j��Ix�z?����Ȕ;��iu����
t��L��������d,
�ӑҮ����2�$N��Z/�5(y�E??%�3�H��ӱx��)���Nr[��ȿ�S�������/CT��i�K`ፇz��J5~�T?
Ѭk�5�z�+��1�� H�b�Z�����[G���rD��8
�/�@!χ�m_�5p$u�I�oB��0� �.��V�2jc��mGiI!�2��ϔ�K��8`��R��r^02"�?;o>��=�z�����I.�ϐ)��N�������S��tiݎ�	y{%z��`㘽�)�X�]֗�$��zJd_,
p�h��mQO,���&i%�����E4���w�5q����.F���$�r�܈��K0�������W�eO�^�
�Ew�C��
��C��A�z�r�7}�>�9_��:��N�u�h;�xr�D��(+�#�ȪS���h���h�h_D��\��5��'$㒍��E��/�R:J��p�]��t��{v핵�a.%K���G��$�著��차�HD�8�gI���>PT�����A�f�k"��8�m��:y,BbtT#�d�+z�mb'"�)U�"3����O��p����T�$G~		�9#��h�Ϝ�	@���jN*?�b5x�8e�'a=gH��)�a�(w(� }�x倄� ����3$)��Lڝ��2��Q&�y�����i���{i=�fE�vIT`u��JT
��&�].3���xY�j�����"��i��,^�j��w�)a�䠘�@�_G�i 8R��+���x��X�ek��5����TF���J�	�^t��S�4�Jҙ<@��
���gT.Be�H������9k��@I�)(�¦�}w"_Y���W�1�A1Py�>�O���`�BR$�0(I�A���5D�;��s�����R���?�O�i��(�;98�"N6�d[7*�A��RR�N%nN25ыm0��a�W�\{v�ȈO<�<�'��86P k�Y�ci�=`$����CUR\����������i�#�bUUJ�M���TtoP�M��$�a��F��p<��gP���=.9{bgu�L�y.FT��¼�r��v���#�����և�2��t�ǎĮ�n�%���H6A��Q����Qph�-l:+)���Q]�aÇ��@B���w��bD�R���!�")�ʊ�6�X�W��^V^Y b�F/��8��h���5%T� ��M�$�<�_,nB6�zc@ʬ�1����J���� TR�!���9�*vU�äv���U=h6�� L��&%EE���zIb�>��P5�(u7<�,��!�P1S��B�MP�'�X�	ͻzbp;�NV٘���(zoEE%�%v����� V���Q�٧R���̹���ޖ�Ht�L�Dm)ńD��R�4¡����,�@�7O	��Z+!wFP"�P�x��< � р3����� �G�MR�¿90F(;�����^|��r��ʼ��34?�:|$����5b�`kR�x@<�a���y�*y�!��%!���rY����\{�E�4;/��R�I�#���t��PqK�5VF�o�wb��J��BT�,�8���d��ನ\ �0��W��]=�8�HW����PD���Yl���j�G�L���J��$�Niq��ӧ��U[j�UO�)�`i�+)��� �F�����,Y�D�&��b��i����ߞ�s7X�%��q	���_3�*${��Qs�@<���fg�au*�zĘ�h����J
��(F���&w�FP^U����H�F<���@��.�0q"v�Iz!Q'{㱾�8��zx7λ�
8d]ñ���!�AԳ�`KF{PYV�{�%ަ7�T�O~&)�QR㾬F�V�l��H+"�ML�x\�,TO,� .Z�U�H%�G�Dr�1j�j�fTI��O�s�ϧ��0��S�&���"I�D�����x5r-mU^"!X�!��l��~-�������|��R��b����T�$i�b��iX��{��!�4�]6�Z䰌�\�v�v�Ũ)�P_�,q�����&�1�|��TTC(e ��v�
��CT�7+����[��p��_5G�ĸQv���K�C�T^T�ו���)��5m�<?�,E䅴k;9.�B�D5��=�4���k((��%k��n��
t5�S��Z������<$6.��'�9�I�-��0�gB۱sN>��-N � ׄ�_fe?[:�ʡ�����K���o��DD�L�N�vg0f� 5�lc6����`��|��1q�xt4��ߎn���)�素���1:���q'GiD�/�N�H!'%����ͫq��s�l�*E'Ÿ���<�p�aJRcw��G��LEe��ΊG��:0qd��b�d'i�$��q����ȁ��=K>_�L`V�mp@�;N��n]z�4lݼR.s���UP�g.��j�75!P���������p�2PQ�D��7����|w��'��{$5u�����=;�� .�t����$��mܾ��q:�n���s��/!@U7J@�z1�܇��f�#����c���t�����hG�zP(���+~��?��8�IB�4��O�u������������8�=����/�E�9��/���� �%��B�.�ط}={���ٙ�!/	#�Ɯ���_pBb08Av'�JV4��*���������ڹx��$*�ߢa����@YY1���$��y�
�A����e߭���W��%s��G_|�D�C1�^&�㶢�;���˿_-�|���Se�l�cb��������W��6.�jG��u�߂�b0�rK겫��`�F
�>Y�W^6��6<��?�ٗ�c/�A1�s�?[�!9�-Ln޲U����ɥ��/p��W�S����W��b��� ��4��%\�B�"��b~�b�v>�"��I���sIX\��Y�=�W���ghkk��֋��]��6���%��h�"�H�F��ޖm;0e�@����r?~��c(*(c${'����n�.�n%q&|��H����˿U� ��]͸���������H*�S��ÐA�5˾.�z�v 8�C���TkE|��b����`Ӷ�J���s���b��mJ�����V��4�Y��,X��W�Tֺ�� �V���/���+��b�	p̈��'��	c��J�3F�K�ev��q*,b�.�d.~�������JK���_c��`quI4���-p������G"� ^y�-\q��i�*<��8����y#�B<|іg��z�Q~˘�:
l��"�p�Q�r�y�F<��=*���Ԩ��A4��C��.m-��y
�V.<�n���w��7���K�G���{+���#:؈r���f�� Q�|i X�[�����c�XTZ�[�/��1��Ĉ����3��ʤ��ķ�aEe���"���شk�N��УDaq����Z��YZ"��,�'�iܘSQB�q8�j��t�<��V.[��)�O��MZG �և�~$yV�!�K�My��?���fM�`�]R�8�����PҐ�T^�X���	���HJG�2q���
<��s���ף���?��;I[x�)��&�'��Hk�\����Ȥ4�u��䋯U��R�SsC=���ɝ��v�ܰv���&���.�����2:��@���x���}��p�BmY�=rhB-��N@C�����e�//�,���7��u�^���L�<�5CB{��w�Ҽ����-�����3�c;3���C��'H��]���ҖR7��B��n)\��8�ͺ������y�	��~ZJ�3��_y���9Uux�ϡ�H��PHs96���`���Q�8�Z�}k�`��������aunehP�a"��y軇�쀫9�m�+`�h����c>V~�.~}��JJ���I�]��y��6ハ>eÐ�𿲐e� �x�9�=�'�vac���-T���߼�z<�O>�j�5�#��j��{�7q��G#Gõm�J4�����ø���4��\�Zܻo[  ��IDATo4t�j�.8��jSN*<���8��30�}�{Ϙʵ/�r�͛��z���XE8�K�Y�|�#��a
�~��~�I������*,���F"��[�����b>v�#qb6�`c"���������#_�o���x9�S�=��ی_��!�?n��e���S#�榪�k����7�@Cߋ������ƷÝ�VIJ�|��݁Ǟ~�x1�r<Ŭ텸kz��q�?�yg/Bǆ/p��oƍ��~�tS-��U���[��P��:g�GL$�6s&n���tݵ�R�ټ�f�z{{�:��砚aH�>�V��ȳXN���!�Y�p�cIW��~ȁ(O`���D�eδ+��z���̼�۾B/�½f��X�:��W�t�#O����ģ�0}�ģ��۟�s 0��	˗��[g��a�q�Q����U3�H}��:9ũ�������W_���nz�V�Q����Hk6m����WBF#׺����y�X��;�`�G5���D��i��UUր�����0*ZL�I3	�'(�$��q"��x��v*&���6^R��|Yw��nk��۴�3�#O�)��_w?�+/�c�C��܌�V�_n2�j|���ǐ�hJ��iі������
���;�k�y��$�*�u��4�\�:�IV�QK�5��ʈ��ց��	���X��+�亪�a��k����}�9�(�F�'èw�Z�pϽ�*�u�a6�՗Ǩ�A��0�hj���y���ܖ�v��/��?��\u����_c��6	��E�/������e՜Ďie4./&�x�|�%�R�[Ôbm�H�P�t|��7n6�?�Az5hiP�@��i�˯��c�<��'B���~W \�x�������6ËZ��r��P��o렲�(����>b(s��+W�!���lP둧�ex6�\)i]v˫��*i|~�����o���)�Ps�GE����g��X����٪S^1�g�ƛZл�x%5_�$.��4L}�Sc��Κ��ͯ���hT;W(~3��B�X�*�Z��;pم�a����&,f|���f�Ê��14�i/��0�J���J����@��#y��|�[��|�]<������ahh���5�v�y���ɾtǀ�ʥ�J/���a{���f�2k��8O7ֹ���0�+j�I�pm��x"au�v������p��gr��j���/k�}�6�w��T�=����QZt�y��M^|�~������X97���e��y>�b"�j�.� ���T2���Ɖ���d
-^�"���2�����[RTZ�`�M��=SK�U��=kL�J�y��&�F2<LH?����=��6|%�8T	�/�\����b,WIL�$=C;QLE]�S�,M
;s3.G���@t���<�h
�1���wo���u��[�`� 4vp����V�x�m|]�eM�Vƫ�����>�?Tikfr�&���Urt���[��<���=�����7>\e$�6;$��uw�@��.��G4��^�&��<(=[��V�����
���a�Z%Ao�0����ܞ!���&B������rL��ȕ���v��3��sW���I�򧿙����+'U���ٗ�O��P��#RQ��|���7����L�l�J��h�#E!!p8JN9��@'�1L���o�����P!觃"��YT�L$S�Ұ���mZ�^?�.~�?��H�t�Gok0��D2 �8tp���/J�+��j�&\|�?�<�Y���x屸5"z����?��̶J8�P7�(���Y���o#���6��҉D�lycrc�qq���[���/����SD��EB<��s�K���K#�$|
I��༔����H�XѹH���S,�xO{��g3p�l�2(ٺ��yvL�:����;�7!qbn���om��Ha�]61j���4ol܈�h��'��%d�[�H{�9�P���Q�ӟ;��x|�d#����Mq�>�=�0O\���{��h�N�Xz/�@%�<D&�b�>�4`b����N��a��|[�1pi"Y�|�*w�U�1��p ��M�yJy�Ck��S�1���������`bҙ���1[o���=E��|Œ�S�*vU��>��|�$��t��s��KѦ��A�����L�h��&3>n�T+�ڔ+�
��$ڤө!^����Dee�2�	�Z��N!��$�&)8=!����g�tf�G*��X�5$�	� 66���/��,��GT����2Ӫ&E�'���%'�%�_�?k����5��+TY�?�D����m��G�b�7�e��c/��a�q�L���j��1�%K��2�x�"�Vǘ����歆Yg�;>�"(�lԁ�����y�1���a�*d�)��}�+�)]W�3
��m���e�f��#g5�X���5g��:�bw�YZ�f�s�W���@�62o�^&j�����]��D���
�����0�!�i�� �3�J<;.�-|���m��.K��3*3�(��o˩�}��-]X��j���A_��򞌤����44S�[��P��蠫���
�_pf������k�	��h6k�b*��p�����z��������o�>��r^�hF{nnE�唝��b����e��ٜgk�ҽc��劎�)!V�֠d5N�+�s��e��WnG�D�~o���|n_i/�f�w""Q'�JP[�XzӼ/`��O��(pJƅo8)
	������e�֚0��)�{��2��͍/1��N�J��Û����A�|�W#W��p�]�����\�\�cgQ�Y�G�9�Ncϊތ�����T�<VQC���\��+�.��+�n��z�����(}i	[��>O#:u����c��91w�n�D*�(k�ì��F�Kd6�cPW�ؘ�:4�NBcM(jT<��!��˩�Z���SH���(��l6e)P�I�������h�@<<))���V�z��+����=���b�1|nCS;8�ocJ�#1�o}	A�,y�/�	ǌ�C��\ֺ�.�I4(&9� 'æ�)S����,D<���rV���	��RF�Wfk��7�,�P`"�p<e�����G��P�{W�CB���*܃q�1Ѩ����;E����X�'U�//�/��8���_q�V���-֩t�aɘ�d�t&�VSnF�ߘ��f�oOco���f*2��t ",Hs-襃��)cCw���34~!͂C�ˠIOu�Jy=9>��B�k2�>�� F�,��}���ʱ��n�H�DX䥁�,C����I�*�Yck�v�659����j�smb6�Q;�����x�x�	�C&Q캺��P�KbC�.�H�GÎY�va�y3콪��0:܇a�(}cCD�5f��Bˌm+o�yӄ�w�eFP����zI����jԑ�1һĴ'=��" ҟ��J���C8x�=��	�!��Q|���k��li OsU���Uj�W�³8�ݎ�w��g���5k�Wf|r��wr���C���{�.�k��]�{}b��!>���BY7b�da�V	(����;[����u)�������Ӳ[t�~��ʋ &Ņ��������ys�X�A�yjo}��O�������Ƶ�!c��An+��[���QG��3f������5$=����e'/�Ƣ��8V�E�یCݏ}"��k�y���w���-p�Ė�#lq��\:���Z}�1�}���K��F���OP��`�[4����>$�.�(TKN����3%��R���z�����=/��Q{�����Dl�bt��y�!% 3�V��D�=��is�󎚝�Ŵ�Z�:���q�I�BCu�%y�?kh��g
���-7aa� �u�:����R]E9�;�랜L'PWӈA)2���_���)s��l����f45i����چ����X�|5�kkQU��E�����>>]��1}��^Y�s�������V9b߽p�)'����ɑ�x��4|?�ůP����͖������7��P�2T����w��B�gXե��~L�1=�8��0i�a�3����:5E� )���}���ʺR<��gZ��y�\�u��6g'���ʟv�5�h-?1�3O\�yӧ�C$\f|�������9Ǳ��8wRy6I���G��_�lI�]�����L�N�6n��QYY�2˧8khIq	W������3Q���q&l㕈V�����cݟe��(A�����J����7�����P#k�ǢA(Z��� �>�DvoG����C�?�c��ⷷ�ͨ�E�j��Wˌ0�Oc���}���C�F��� ��ik���ko�O�M�-���k!�,ƇFp�����0ֹ�1��q)BkΠ�+.�=<��yΜM�kv&g�W�!,<`?L�a����2�=Ui\���u2x�1z~�/hp�	�VF�p�v�;;�jEr��FzҌ��pA���������ko�ظH���3�[�T�.<�t#"��NZ/�O�H�z��o�_��-�&m��߯C�8�q����K��;1�u�Oe\�lD`�C�����W�b`d�D�e4��0B���A,:�zd^�QzwAX��-��Q�PQ��>
������z�R�����k]c�SZ����10��K�$q����+L�W?����?��~*�=o��%W�FW="���~f�j+12:�u����1�C�7��Ϗ��TI˗����-�ч�i��ؼ�g����\�G�����w.�{�Q��Z�Wٺ�.(���0�6�d����2J�	�1����}�8�c���8%�sBX��h�
|���==[PYc��i�4 ݈��Y�������FD+�fҲjټ��4zߦ��c�����@�?�G��=@c�y����+��/��W�\����y`��e����Z�{�噬�Q�*0"�m:����W��-��|b��c�Ia��{i����ߡ�����Ƭ9����Ai�����\	�J�+V~@�����sf�����׫�J)�-�,ߔ�(����M��q;3뵸)Lo�ӾߥA������rq���h����f�믽�۶Y�Z��B#U����6>^S�	��g_zۚR�~!�yxu��~�ш�H��&����l�OS|��iz<��e��՝�X��8�@�n��ي|�m��B(g���$p!�cϼ@x�Ё���)r��ښ����*�d�r,1���Fl�괖������K�!X	#A��J�����F�m[�)ƭZ{]z���p�7|�
�~�=(����]|��H7����S�h��Eg�F�B�՛�Jz����E�p���#�����To�֙TG�*�g�R�����	c(���&ėR��G�x��e�U~����&��N��4"ܣxM��E���RX71؇���}�q�C� �9L3�ռp߽�Bto�d�R��9O =�|'��M9=�^��g|�1I�P��rJ�e�8��0{f+�{��ܶ3���m��3Dke#*cQ'x���{ �
��-m ��0���qã�����4�k6Ha� ����O�so,���>㤵��C�g骋�g�R0�Θ��߇>>GUC�U�*h|�oހ�o�!~����#��A��&�p���i��m�u�nD�c��x�]X��D�.�N��1�|�9|��k���k��.~�u\�槸�u܇ז��Ь�f�a��;����}����o�`��0�+!<����[�gIX�_�؂�V.Ƕ-��F�%�p8d���`��(�vt�T��jWW�%�h1�;f!^z�MD*j,?�l�4~ɢ� ����E?]�ܤ���!NH��-8c��xc�'�����K��������^D�M�>��[��+]�p�Q�In.PFk]E/r>�d�����N*E8~
��Q1�Xދ�>X�Q��Y\��u�p�ֲ}��O�CO,F��M�F��3o'��� '�Y�$/���܍�-u8����ف9��o��/b<����)��?�}kG������[b۶�6/3o�N�c��x����#8��xo�*��Y%&��N:��:�Lm��K��;|��j�sfN��Y������5��O����Pg�,�w�����H�_z����2$3.S*��p���Kh9��v��G`�ko�x�R��^���hk��x�i�,�ǽwab2�X����pʜ��Z��S[���b庯��~匉��o�=��3RU���1�����LE(��NӦ�Eǚq�؆� z	/}�1��h8O�wO� �\\3k|����;�Z�Ǯ�|��T�Jo������8�{�y��Ӕ�(�� f��]y�|�� ]l5��o~�3B����8����xi�Ȧ�:7�#O=�HxUiZ���x�wp��Z[yp��&Vn���9 �<�#�b�����D�5UH�x�̘��~r6�[M��A=Cי4J���-D�#$��sq���3t��Z�a�>��ghЋ�����s/3;���,_��9Gz�M�^s�%�����a�U�:{�ȝw`����B�����ۿo�����U_�F�a�����w��B�=�����h`@�ڗ_t��=*���3/��	s� w�;�:�zÏ��g_^F���ћ)N���p��nDO�V�Kli�1���D��V�1,<�#9j1�`"����6ɪ̷����u�;�$�o6��ӧ�w>D����c�=�Pz�^��3h�o�՟��+ɧi�_�����?���QkK=^y������#A��Qy�
�v��>m1�dbV:��Cq$7X2LV[G�p.�,��N8�p����;�?���j�$/�|�j~���;'��DS}Vl��
y��8r��i�ǡDrus3~����;�0����y��=���P�D�����`E��c�Д'!���u;��g�no�j-ڛ;Fq罏��x���,%��	X�Cs��*cF��=4�%K��f���-�dL+�~�E�.Z`�7�C,�ҏ���0��OC�B���x����:���܍چF�	��&�����(�.ŜiMF&4�,,_�A���	Q��OL�����F�!4�L1�	z�M��xt��E��c?��}p,e��A:����Q���}��|=��
D�q��ٗ��6S�Z-��e�&4�v�Y'��T_e�P�v�?��w�T�1L��`�ˍb~�T��{p�a�̟��j���\�(�`�tq:��|ϼ���N�l����Z<��K��͹�vL����^G6���B�:�����~2��t�y����A�7���4�Zo?�\�&X�%�J��dHR�����N�},��*֛��~�틙u�����λ�.�R0Le�`oà�i���_��XD.�}%�?�Dk�t��{��~�J��~0>\��}Ą�<��"�i�^�`�w����ڭ��1���������j�v��F�mm���8����V����n�M_N�O��cO<�
=�^��>Y�]Y[¼�	4V�M��:)���L#J��/�➇�˰#�4��4W�،?��o��.�����1k&�aQ.@��	Ɯ���w=�<B���x�B���?�v�7q��r���0f��&��+�@y3~�?7�;bz��������꯱��fZ�=Vnl7���:	yн��Y=�~�St�Z���A>;���b� �� �;�͈�.��LmiÝ��#<�r�����y���������@-S2U�%����=�'S���R��1�R0:zM����5�*�� ECP0z]j���g���к�in��/PY��hӨV�������c�}v��W���?�:�wU������+�u��4aR�zI�{�'&ѩ.Ȍ���^z��6Yxy�2��I���
�59�����AT�+�����W^x&b�r~~ԪV:�yz�4�W�qF�h$����?YT�N�w8m�jv����@�P�f��)LZ�:g#4ȯ���rx��8'+��M`ZsV�ـ���Ѩu�7����bѰ5�}��*T7�J�1nK�Yzo� �1�˗�;5�Y.�	�+5n��sУ�;fJ��g!^|�k-D���"�j�[MzB�c�J��R��/���5�3�v��,���I�/H��0�7�D0_m�d×*��a�6
c#D�v���Stf�$�4�s�3Ѝ��qxS�%CD��Z9m0���e�X"�:��P/��9/l2K#RcI��	�&2��#UW�^���OW�����b�����-r�J���ћ��|�z�5(f� �<�w��002؋7[�U+19�AJ�)A��Mc@��J��ЊfU���s��l�y�47��?a9u��j�������i��%�p����K��/m,;��3�1^5�i�[c�"�!�-'RYş)a��٠�����7F�H4���>kHRk�ˊ>�'Y�k�6��	����R]����T�\F �)���sY�hC��k>@@�3�-�v��U���n*�L}6��1pU��E#��3��wT�T �	�85��D����I�+jsn�:�*���Q�BZ^S��d�5H��I�?e������Pv^�#��<��{�O�jb�٪�vAD�7ݕ�u���Y����:4��(��1�Q"�H���$�XE�5j�J������%I$������c;��a���-×����c�0{�㸊���&�B!�K$����J�$��%��?c����p��O��W�T�N��B��rX�g�f�C4��ҁH���X��DfQ"���)%{c�$͛�S�r(J�M�5��g(�����p_�����B�����#SV���� B�������"^U�}J%��]=#6�ю`�܊���BU_��(�Be�-y�|.�U#�Ǜ3^���:��LN�p�}&�����d�;D�rU:#��z{��Tی�|�*�aJR�n��I|�ܴV�H���\��CɨӖ�H*�m�:NE�&-�Dr̔�4}��C�r�7���[b*�$����ցR�nH�6?��f����(AOXVY�"=�ȃ$J����(����\�	�pe�s@,��h��IC�5�$�b�A��q�F�G�$V��;|!�=[Q�<��C�F��G��X<j�T��O�6W�(�ГG�+4���2g�D}Z�,�8� �66`0ىHM5�z{��h�Rb�
0��Fj2e�o�ݝNd>Sb}r�J�m�b^<��q����Y��$Z�Oq�j����G���!=��Mk�3�)���p�*ߎM������e%oV��������)���ށ�3���7?4���1|����A�./���s�|�6C>��`�\7hڱeD�.^ZQ�k������_"�1�,�/��M�g#�g!/i
��4}J�K۝H'Ƭ�����>���F�G�ӑ����RD[��;{:G����0�д�gHZ>�1��yD+�Hd��4�!#�VZ�!�VL2$�=���Ћ��!"�����؇�v�7�B��is�y�f����zv���4�V��vD��|�B�a|�C[e�);�As�rĒ�4�":�ysfcʗ[�)OH8�P��#��r�!Kx��w���#g��������S��1���[h১���{8������+����2��>¥C	iz�C�������F��$#��?��5(��.��VT�x���uv�5���W{ϣ��ʣ��"/�!�e���8�ŨU]�|� ������_�������:Ӯ�R�5U�]=�
$)�P���~
��/g
#��ц��� :=��Dm|���X��p���z�	��A�1�N�[���{L$b�4a���w���D����dFQ��x7��B��k����&I�����k�\/��8pl��<�U�b= ��p͕a�v����(�iz)j�������[�F�f�"2�J�ea5�y��Ito�QxWnJ�*�mz���X�mzk/�rA-Օ��k�4/Ġ1�:���pi�N�H�T���1��Z�@��uD�A�y�"���bتy�Xp;F�P<=ч�3-��N�y-��{�D?�8�tIF��'��?�4�Y+�jE��n|����'��qz�L�go��u��x�[��K�������D�*�ws�Ax��e�m�!:	y3ԇ� ֮E�(!~�w�h�VC��w��e��}:n�ۿP�Pia`U�}\�k/;�DbA����	Ջ#4*��X��7bN[����t���}�?�:�q��WXJ�%�E���N�٦��0���w�Q/�^�����?:����&>�7�K��Y� ��`?�?�$�?�����_�W�M<�W���;���h��5����K 'kts��0v�?��iEW���w����WЍի�`�E�5��g���]L(�LL��2\���9����!��$w���K�x	%u0��S�*�U_��v��i�ԭ��4Uct��Jo�ކpe�5�(�x��q�A�"L�př��Χ�E���'j"��ւ}1cj��9z���Ɍ�����}�c�s��4�	�fO���c�H�g|��˜p���r�2�|��Ʈ<�e���hk5��iյ��zg�FL�`N�Z�}w�g���@�e���	={�n����~�v�ϚI���uW_�G�}��(�Ì�z�o#���D��/�J�����{��Gp%/���.=�<���<��9�UG�Z[�쇔�5���Ͽbk��PL��G��l#��>�(T0������x��;�l�٢��&���_��.Z�Kd�pc�m|ם6��k.�[o�����3�D�8f�� �!������54�W��'�W`��Ga��+q�qG`��v�z���Ģ'`�gXapE]-z��Ot�<6ئ��.�o�&����:<������p4�{̞�ٺL�1�/�Q]�y+|4F��gx��p��`헫�_���I��1"Y1aUb�]vB[s=*ba�O�ɧ���)Q����^��(���ڋ��;o�%��N���Y�0���1ޱ�V|jc9� ��S���?�����p���a�⧟Ay4�i��8�ګ��Ո��yν�R#�R�%�X������N��t���}�%�ʘ)$.:��:{�) x���B���غ���яS�85匛z������AIg򓀅��埣����
��f����?B�q���&s�"tm��:��l\o��$4>�t
��w.<tz�7��O@�f{Wji��A_������Q���!�4�Y[��)�T��s/���Ɩ-[q���SO7��;-n�y�PS��mAcc#y� G;��l����c~C5��F�����3�p,mHG�I�����q��K|�����ϼ�
�dG�;N9�=��s��tۿ^ge�/x�7v����d�O|���,}��|"=�j)�>w�AB���v��c�M���,^�t����D��j��Ye��g��@'�lۼ���6`h"�G�����\��>����=���q�������6x��&��8���^0*Q
(���|�x��-�b��q�׶?5-('��l�c���-|�OV�%�[���4�%�����Oq�ӱ`�9f�G	�3�ǵ�J�ܸ����"��\)'��Ž��Gq������إ!�sEV3=���!ZU����OcKG���	m��F��;665Xxx�Imv&=A䙒�R��w���#�s_����#�H�q�C�q�O~��5_��E����e�����ޯ&�GF���Ĥi|e��{���"L�E0�i��m�m!`f��梊|�OW��{D�B�>�����be�w�\y�y�^�
�\~.�o��/A�Q:�a���A���cʗ�e+�j���܁�������f��DL4j��Q�/�V�Y�ѭ�p��{����ٴv�Y�T����G� �����#�������P�O���9�e]vR�����5	�c`/���X�$4��9��d��,^~�-q�A�n�Lrn�/7ԁ�H�2�#��3v�8�a�)�Q䳄	K�^�*N^t"��V�0f�M�%2ʃ�u�:45OųO�`�_�����KS���]��G�,�s���}�r4��S���I�����<�V��k�,CC˴���2���xd1~r��бm��:j���!��n��[;:�����D/�K>�*i���F���S�ޕ�c������#d�%�T��ɉ�8����%��gJj��l��o����aƳ:�p'�4���0���{�i�xQ&K3C���Q����>�����c�q�[���1�I������dY�H#��B+���r���̋����܈�[7 ��#�u�,�:�}��U_��/6X�0�CS����7m��C���J�C��:���J)���yF�-��p͝s&;5�X�<ú�{�5����5uȊg����e[�������ϐ+)ʀ��!Lᙗ^��#Ɣ�Z���T����uJB4`+׬�Ko��He��i�OQ�-�3��P�ﭷ�'��;1�i�Z~i����ʚF�鯷a#�Qo�f���A�|u5|��p�5W`jU%�x/��N���vgx����+���e�<�jqs�Gh�dH~����?�!6oڄ�͛Q�CH���ǒ�ǽ�ǆ���GJ���E�q���[p�?�J�C/GO_��t�������ޠy�m�ۑD����O���I��.��mڸ%���W_Ǣ�dl�1���eΆ��=���<�6E����b�.{����/:�[�Gjjn�g���|r4���}	Q.��C�7(8����S�2TU��|���:�V�`@�O����{�y����~������$ʫ��²����ZS�DB]�!�CN��g����PY��L�jP��L�
��|$�_�}N>A�y�n����I�7����F�g�R�V�R?K��
E�>�{�3�"<R^c�J���ϗ�Qڴ��	�U[<n+]Fy9��5u�!46Eģ�������{�m0�Ҭ�.�w����C�إ�r_�f�i?_�%G08<�{�Ym�Jf
>����Eq���e�Go�@�?�0=x�
"��6n�qs%ȥ!�	`g�Ec�e�
l����c���F	�5 �8�ƻ�*�YCS�35j	Ȝ3�)��iЂ���ށK/��9��Pچ�4.��6a6�Y<n$>�J�= V���I7$y��~�mvЁ�M��˭�j���Ƭ�f�z�j���㷰�V����byˤ�;������S�Ik�R������C��1>��k�(����sp�#O`��sM�3�2N����?�W�j[��x5�p��c��/��_��_ร�v��чv:.͎}��稡�Q"w��Y<#F�\p&��D?5-S��7b��w��T����p}6Շh@�<��M�i�.�*I>��k���[�^j��3ʬa*e�@�E"��_��1k��"Ԋ�_�z��Z����p���T�7�O�?:��B=ieHyoq8�͍rZ6��������lh�Z�sVI��}?��'�Y�'gm\Y�Ƒ�*d��6hQ�l�Ў��g�0���e	Ǽ�&G4�Z&V�|�L"��qdW���h�r6����L���K�%X5jit�}�he=r.��t����hs#�c	�¥X�f���}ҥA1m�x��^oiH��Ryک�m�7�����!S�4��[iW����j�+3�%�h��3E��D%�@8ND��'_np4Ex�z�sz���(��Mu@*Y�)+�nT�� �t�x��O�"�w��wATq���LE欐���Tmܦ���ҷ�^ǲ^|�b��_�-s��cƨ���
�Ç��)����x}+�~�%+W�{ӝN����5�o- ��ڤs�IJ���T�6a�-V�v�(��7w���4Mj#�>��Z,:�&Y��fq4L��]��r>;�;��ct<6IZ�X�\��b���O��J��	��.�vts��lC��]��)c�jp&�]�ФIK��ä��c+"P��[aL$���(	�U�9BT�Ҵ�#�Q�wuwB�MjQʈ�Ϲ��A�c(7���0�ִ�(���)%.���N&H9 �JW���`�ʂk-���l��]�YŨ7Dׯ�¦B�]8}�����ao
���˰�F�%9����t�e|p9���"Ѽ�_UI�3�l�P�(��9q#�����Vl�*:�y���������9jz�A,��0Sb�b{���z8��]熈Jh|�eQ����LIXJ���LD�0�@z^M�\f,=A�{�`�v!��<`&�L֊��F�������Lp�w�����Z O�#����SSޡ�w�A�Uu�Sxq4�2�:����%9!*��@��-�hs+�)L:�:h2R����|��]f9	��Ș���%7�f����yh��o��6�rHs�G���]��3��2c�ޙ|�!�Q�S��-����j��r�~���|�b���.��򥭱���^��Ƙ��bє���T	�=�DkJ��2+���<��E	x�|�,q�'�z-� ��cTe�{O�y&�0I�2��Ah5P��QLO��|�����7�;b�%�������~����,�-	�����GK���(��z��_3���S	��k�������׸�Fҕ�zq�Ċ����[°Dbc���$S��Hg��=F�+�A������T�� )�ē�)k�Y���'�%Q�,R�o�_t�
�] ���[W�%C�J0�r�E��D�k*-��U�E2t���p�!��
�����+XK�2�`�&Z�K[OV�6A�/ϋY��LL�6Rfy	��J��D�G�	��-��1ck�@f���x\颪[�<:�[���F�Ρp.�}�t�����y����^����Z����J� E[#�|�X�`W�m�@��P���q�-w�Ky�!@RBzǡu8B<%���M�ʜ��*x���)�o���9/;�4���rIhJ'�GF����|0�,� %��b�2*��rc@ݖ��dx�3�~!�4�Xh�D�*}v��v&z�� |�}�YØ��D*���fkF�����nk-��r�����ُvY2<99n(A�/�6!��3Cu��_��khӻ����5>>��	a̘=�Ш�(e;���q=^g�J���xr����8��C;)�+��@����v��$f�������c����s�Xb<*:���ݒ�
O��2O�K�P=��.�8-sҜ��<��W�rTS�z7�$V�T���
��ܬ��:�B��M{E���qx�#��~��	�'�#�-�w)�XQUm�o��9�y��ө������NC2�2f#ux��b�s��� g�{���Kи�K!G1o�,�ҫ�<2<���-X�v#=g��B5\�1n��4.	��$�T1�yAA�4gk6������m%�%y0큦[j��8��hX���'J�j�Fc㶓jC^�$�c8d�ːO�"���o/d�@,Va+���+��`��+�e�޹���rȌ�c�=wA\}0By��Q9vv�`��mWT;�s�%� &1��1;c4�͝���.��U6�r?��T1�.�`)���%�5��$�M�a��w��=��c����)X���X�q��_��\�RW�;p���?��G($��������w��7��a,������7�WE�o�`f[�]�@A$�lݶ���?�(ע�Ǩ���(+.�[PH]H����7��ܯr����J�嗿AyM�!�΂5H<F�$����v�8a�F�%*ǉT��J����`Ū5(/��*[6��1�Kbf*�'8t��8���_����ƭ������_�bQ���I�Wx�ŗ�3�0֞B	K��Zq	��wv�ګ/�g(Z�]���*�Sl��ųϿl:�@QJf*�adż����Lᅕ�nr��?�	��HO=���#�T�� �J�Z����X]��Gj����Y%���	�|�)���˼����Q*6͎�����G�VPL�ҼL2T���٧���{��ube�J��*Kr�2<�W]|6���MM
uDf5����'�g_z͆�R<�2��O��Q��ƧG��p�A�`���4��B>���3h���/�Xޠ��DFUc�N�T0������`^X��&��ϞaݛBe��>w>�8*jj�S���wrJ�ȉ�-Jt�?I*F�2�gh�6��S}���b����D��`��Yd�.�)j��Sm<;����bL�j1�����s��gA9.3v;��A�*����؅�V�-Io'�����n����=�__���41m��t"���8��et�-S�1<2������Q��mlj�Z�c]�j����όS��E���W^���������ӡ��ԏ_����ֿ!Z�d�:B�K8�^���}v��4�����M�r�{��ù'��_�Ϸ��3�M�`���H�Ao��r�O1>�ϻ�5B���qG��{�??��q��	�7Vx5h���Fn����sNüY��$oi�$���<�1:��6���k��K�%�$}Ǯ��b�}�E�8r��e�2�mo7��":����	��[*�(��JS����%o��������`�ޤ�m���{߱�6�F>�Z9a]��_�ҋ�����5����:�p\t�2}�A��P�2���n�C����$�� .;����SM������A;y�#�B8�CxaG	>$��ϫsO�>�����J*�v��T�3���?Y^�q��e��PFU<������ğo�-�g�V�����ɱ!�w�"�PoN�yj�͖�q��t��xu��Mn��;�=�po�=� L��Hc�v�#��\EW�VLm�72XM��l���o��<�9h�=m��/M�^Bl=c������4�w�s*��
P�PbW+�kz�q��K�6�E?Q�V(�<��$���_�AGO�u�*W$�\�%%zx�.��Es�5u�Ñr#C��R_�sN;�>�$Qd���ғ2Q��CDsC�%+*ch�2����<%	wm�w.8���^�9�B&q�j@�����Y��*S.��jz2��p%�+
8t�}��g+����K�5��@�w�Y�!�S�p�i�TTVb��½q��k�����Oh����F��s�=v3�5��gWQ���шir\�؇�?�N'��<,�X4��\f�{ݎ;��K:�Zg̴�'IB(���,d.�A���s�����hE2E�.�C�:�Ӆk.� 3h0�Z�0���&��UR^#���=
�D_��ڐ��vy%����y�;�4��}����Cg{���XtҷQWCX??28dJeZh]hMt�&�h����0|A����+L�U�I�����^AX;n���ռ��<-��",�$H���]����7-�T39).�*u��{��eԋ��k�P�4^���a�.:v!{�EK�8$�+C���|���5S0���4���}�V�?w:���OV��;�,�-]�Br��J�1,���ɍ��͝غn5*bDx���F4{Ӎ�����h�-�.dr��|���*�po߶.>qX	L�>_����l�!�%�����
"s���O��1h��^Ǫ�����_FMu�et�~H${��N�iHư���:�H�i���[4J"6
��w��d�F����;����2G��k�����S�ϥr�U��<�#1��_�?_��6�y����Q�{�]w����"�9b^x�-Od��n|��9=Acp�CBKcӺӮ�ӭ�a����#r�1�0MV"��NX����zAT>r�o��1�m*$�;m�p��Wa��.47U���
��j|��ST��k.�oo���mtp)~"c��?�����u;á�ڦ���P����{�9��yҪ���tɗ.����z'�$�?��R46�4���ϸ�g2�g�c�R�]p��h���ӯq�M� ^�bNT%�9Dv�Ѩ./���oeN<�4n�RT����KcRƋ9Æ;?X�5+��1����������^�}x踍�=��[�ƅ4�;ͣd(��;��K.��Q2�u�����������҆�ν
]�yLk*��O��#�##��ƕ�]��5u�=����\��y����0��7ނ`�Q����?�n�ޕ�}�,����'�����M��B5=ɘDx��k�<=�(��W\nM\����}�5,�j&Mȍ�v��ӿ}�'o~0t�ʵ��]_����j�)B��D�?�c�A�C�"�?�Lz!�|
�~*~���LG�]0��ӛn��CX��>r�SX�n�����x�Bn����c'���B��B9.z��:�q�C�ܝq�O��l���3mS������9&��K�����)K��sښ�RW������T���I�2�����jZ�Tc��9<�AOĒ�B�z2F�(���;0�_�l��v���02>��	w�܇��;7���N�0�߅��|�۷���G7��@i_��5�7�_nMoW�M�b��:oτU5R\'	��vb��V�������_!^�0�qm�@K��м���mV��_��(+�0ԧ�8�K�*q`~���Q�<�V�pm_�`%��q��ǃ�ӌ�U�JIX���ٳ쟱�z|ĉhh�E��v@�1[���܊�;De[142�{�5��i�^u�ظ�K�:�p����{�j��D�+�|���n�^�33dr8C���y��T��+476r[�n#n�����"J+��՛��ܙ���;q��k��܉�˥���ꅆ�{O��t��eϽp�.DuC=Қ��gh�~w�?������/�������.C0VmF#�˙��4�l��7��h��ɜ	��C5�0�;�t�bA�oXk#Ci'�׸�ԩ�H�uY��9]�B�ͳ�Ƴ�Z,���k���zB�8~ᡸ��K��>{�fDǱ���U?D���)|ӱ���D]x��ǰ��~�K�V�Ï>�:6q������.�����ܿb�9��R��AWWf�0�S�&T��S�n��o(j��J����f��j�}=���5���UV�QL&����vz�?��� #��s�'����� �d�HZ$�+����_'�6l2~�$=���yk��F����%�r���o!�gjm�a4����,w��Q�H5�2n0���G��q����`C�$�o�.;ME.A4�܎圔�ʘ�:��?���!��:h� �@���3/����9��i�xT)Q;n�-��,7S���h�6�$PE�4J�۰O�悦��q��bR��X��t���?G�RS���MsD��!z�ql�C�*��qV[�?�����C���1�C,V�?��!E���&
��1��;�3R��J�Cw�*�D�U��i����݊�i-\�2D�*y&���ci�Z�	m�d�n��C�p��Q��������(��W�"4��o���i�B\�|n�N���\��6YV�| ��n�-��ȮV�H��xᕥ���Si|'i$��O(oIx"�\%�ip��o"��-��p���$<���<hm4d��^��*i2gG�T�	C�t6�W�[�*������S�����`�+�c��Z%��w��נ�A��(�`*WDR���b�;i�;�����5�����;�GM\a�&�'x?�y�]���R�Dܔ�)Ի��~��k�k��������_(,��b5y�ar�:�3$Vj��%1��Ǜ�;M8f���(&n���
�������U.�`D9;zà�gCJÄ��=��Kkä�$�R�#�?�������r�6��+#�2�M������{��fJ0�����)�	0֢�S~���ohȈYrf���|�-"��'B�GE�АJ"3>�?�j�zL�~
���N2�l�F�e�,�1��5�/����&}��#�X��f�۩��r>˲�$9�M�٤��i3��ދ��z�2�s��>#��Tm";b*[j��ԯ����#��M[�'�˥����E$�K��Ƨ��W�&jHS��c���E����ҀÛ�䬚�4d�.x���.�=2l�X�]H�<�[�(���T�s7l|(�#QeA�Mi]�#�4�8�7܎l��#��1��a��-�j������v<��*d��|"�������rb��嫪�`Ú���@�z%�w�Tռ�
5�/I��X"U���9�!q��|Y��7"�s;c�.��\U ��F�	42d�T�$�=����ڽu���RbzxR�1��4�[�'/�zz��]�Z?MCKVl볼�ZBܟ��>T�+�HƬMD�2�s2Κ�3��zjl�Q�Z��\T�t�ӛQ)�xW�{\f91P�A��U����� �_���dD%G"�l:1%��h��I�h�3�㙗r��oi����v�i>�[����e�_�LR�C���hBҧv{5�9�/��@�%��颗0�
�ɤ5�H�:���aU�B�tE�VU��-�=�)������8?n��&? �S%�mĪQ�H����s��c�v�I���0����8Ms�����51�렃�E�66:b�$�#�� �u�y^�Q������h�\`U�<�0��2�.�	#��p��:{5+e�i��(���] \+XG��?8:$i^�hM5�C�ڬ���u��O%���Y49Ǣi�����J]|�9��V��Њ�`��2OYQ5%��gh������v\l�y�G��������Y;�_��Dр��9�$�v�rG��-%.�]�`��21a��L��	�#	z�V5�@�T�!%7����z�����@X뷐��s�$!�H}�D��P�%I��I۬�@�r��YmX?�!�{���/-�2���[ّ~��9Mbn���4��8y� ��*Pr.���d-RR���F��9 Zΰ�x�ˉB*c��b�(X���ԅI$G��PG��D��Ms�,�����7�"�C4��{���x���Ռ����0��X�&]vf��w�g�P����2:��J��D��[2<�U�aoZ���,2}݊�
3���1[�i��$1BƧ�m8c=)�7����P Y���A�JɈ���QfdCELi�7���*�X5�Hv��{Z��[YS���68Z�<�>56DX�c9b�@�F�˷��F���:�4���/6"��R5�tP�^��i�&
�O��x�� ���K1 @O�C���؈��^;�������h�:¿r���&a�|�$�1ҩS�`��t�Ob<��8ӧ�N�YW[i$&��d]�JX�ˠX҄m"b��aJxx���o ��C��Xk� ��t����.^��A��q��\+7�''MQ�mѳhTk�I�q�J)�dbq4f�E:���ۺ������ϼ�D:lg!iRp$(n�DO������b=*�cIc'�p�0��9s[��������w��bT|M1D���i^ bykv+:s8B����թ��;VX_<��U�P[^f�z3��%��(�Ć4<'#�i�z���x|�b�C��2Kt�&EN}�~{���ncsFڪb����矉���	c���D��sjC���q�)'r�S��Q��XÓ��pA�|D/�]�Ua�8�9�U�D�3�h��q|?��c*'
UÞ�������6o݆��0|
�!+a��f�@���x��J�L���vTڲv��hni���Ɠ�8�k��ҷ�ilj�(�W��iT<D	NEID8�Rá�9^%*�����ǞG1$�6i)Q}����L<:� ��11n}�j�JRɴ��w�K?b��4��4|�0��P�V\�5��\&��Ն5�	��d��D�#04=��}���_�9Ry�,���1G�XE9��#=��Pm�q�aF�-����02�㌴�Ʃ�ѩ��Dy5��1�>�e�c�Y����ϢSO�4.��m�v�z�{MAʤ�h��r�/V��P/��5#�ƣ�N!�8�0�~��sC*���R�seB9
���#� Mv�2F�Vr$�G�������|�����t&z��聢v�5-����$$"s-觫7�X�'4��c��9�7m".���z8���}���1�C7�����������k��bw`���-+"�b�����0��0L���?��\����c_�3w>�w��zl�o�M��j������@KK�wy�-��n-�&d�\r�O<�(�nj�x����,��(��ȃ�նuj�3u_|��/��^�oi)�;K�p�&{}:'���!��H/>9!�m܂��
1�g�x>������%H��K�F��u���9ϼ��xb�Q����op��S��ю{�݊g�{]	�iP}��;Nx�!��ذqk^�X��zy��9���G(޲k�G2�}'��A�Fi�xP����ft*u�Gۛ;z��BV�w�g�z>��s�ɜeQ�{�E�K,�%kk�Ƭ�6k�֛r�]�n����݂�/9/��H���Z�I�
�'��h�ve���rqAS�1м���6�`7�s�қ�"��/9�`���d��<aY{�2��۰����8� ֵ�7b��q*��{4*pز�^B�,���>v̒�o����e�٘Ǣ��WU�z;p��gc��ߡ��%�x�?�Jě�K�U�X"�6�\�!���|��釋?���BP���x�w�g�5�W^V�k�\/azD�y��%x{�3������ �?� /��4�[v`�*�0���z%���V[��H��[g�t$>Z�	�eI ��eN;�H���*׷����ܬ������%�࣯p�?�`gc#N8�P|��Oؙ���AEY�|��HE��k���㫏�Q>�y�X��6o�Y.pyN�۾�i՟H��ls�1�blU	:�B�K��Wނ�bh��˪C9w�� n��z��ڀ3�;߯]�M[��W��%:�F{����_V*��I��C���y�;�L�d!'�.�.z�*�A?F�{�4
$��h���	���d�0�va��Kqꉇ�i�F\=k>���6}rxp��b��O�vh����;�ŋ��\	E\��G��+.AOC#j�>r�MvE�A�.=�Ӯ��c�ee��G� ��/���NC��#ų�q�1�&��9����_�S��ƃş}��)C(��+aC(â��'��ߗ����7��G�[uv�]m��ų��ր5�����q���o��_\x�����*L^�C��WɊ�GKֲ��6�+H����_u8�Q��C ����2#F��oq��[�E��!ho�K�<�����XQ���|�����r=�������K�,��̓�����$��dW�"N����ÏTB!g6��K+�����E����ƉG,��VC�h"��g��vm����K＋A�,���IB�f���>�
�O=�M(
�ڰ�ʋ�
������K��v�f|�l��QP��1	�z�<|�u��#�݌��>HP��(�Y�m�^��1	�<� ���;ZεM���$Բa��	:�C7_+h$���}���m�C�b��Qx�g%�wK���P��1_�7�p;�M�A�۟±��g1�cAi*�*�g�w��b�t�,��5��[nĖ5�jo�/��G�����J��<rB�no!�w7n��D��p�!����d�/�����a�Ckj0����)�V�:��r��㯾�g'p���}�D���ؾ�O47v��������!n\b�� 
��'��\��+��ā{�9'/gي]�uR	��Ak���C�r)r��E�$9��5��Y�ē�����'j�Ӡ��]�5�8 ���}��a�u�ưB�O�T���?�'"�n�Ǳ�qcF����M�Q��aԈQ��gQ(��	-ͽЎ0{%�>��`ޝ�޴��\�%N��Aڝ�����?���G����r�(��x��/�����[��>1X��~}bx�G'2K+���M[�ܺj�Ⱥ�r���ݳI���[���y6v���A�(+��Ukj�DO8!F�W��ԁl&1m�� �`���G�~�ߔ�/)��OP��-0��t��_E�l�R�b��l��~Y�
յ尦��cï�A+�*+%N�PO<Ƈ�(�ژgUîj|l���u��7��E3NEF�_�W�h726�����K�0�j"�Р͉�g���o��k�>[��d)�Yʆ�hD� ��=�l�r16C�T;��:���_}��MVժ�{ɸNm]ve��a��F|��G��:F��Vc��_X,��	7�����|�n�G�=�p�b<�+�P����
���"�#2}`��o�UJ��rֺv�iz@P�S��#��}x��'f���e�!	ռbR�ٮ�yw܏瞸��DI�(x�� �89v��sO?�itZv��ڈBs�|��XQ�8/��Pu�5q$�\�b����o���������7	ds*�dG'�g{�}�+G�`�U����{l��[�T����.Y;v��!F�O��K�I>��[���$)Q��Ɉ�V$L�3��V��O�R��Q���Jr����X��U.p����!l���'$��8���[q���5KMn^lG���lmڈ�+���jҜ�͏�g�{���2h����_q����$d-��`9Q v8���yI.K���2�"�Ψ�vN+��cp�3/��CDͰ*AaA�2t��+�%_-U��l�=�/pj�F�U��a~�]L�oFa�T~�iOF/�u��uK�@m2�KHe7�M�,~1�	�$���?����S�6��#�ղ!M�}#0���\���\��)cP���fg���{�y�qp���A�\DI�9Y���/�.����� �1?�lP�ɻ~�ӏ: ��K��p�<�]B�n�����2����QɌ	b~?�a-a۱x�2Y�CQ�sk�CB.밚�X���|��$�QU5h�|vc�@<��/�a���v�l�p%�DcZ������@�\vBE*�4	��$x*�Ưl�@8�����]�����c�z�Z���7��^�P98���
s��U5n
���.�<wJ
��z���B�k���'PP5T��%>����\��U����G�J9��5��棉�2�'�n�����%�**R���c��Ysymf��Ko��n�F9m�4�$��$����;�[`��a��*1eb���T
4���״�f�4�Ʋ�^��{�Df�/��U��T�)q�\�M[�+�*��,{��-Q�@c���ӯ�Gmu����6��]�dVX������fP�ÀU,7���#�r��&��;���mbH����0e��a<gr��k�Al�Ig��tN��CBƯz�r���t��B�"���rP}��@�2a�BQ9�m��O�r���9k�����Ͼ_!��3��`R� rxT�ڢ#�����Nt��Qy��8|A�Z_������eJ`T�_�W��Ps��F�r0��r:������V�[CH�g��>g6KJ��ln�Q&���JNH�!�O���ԁ��V>J:Co�����:��P�*&@��X�/~�C'K�?�Q�
�^\�TCj:�W+�V�6U��k���|�H�W����B�p�)��1S���8�&�[�iI�ϼ���s���}f"�ȍT�"e	�k�5{�D�Nj�y�а��z�y�[6?r�lb������o�;?���=��L���_]��V�[s�:ImI���RY���A0�:;Dy��px�����f��x-7&}�8���"��8�d�y�(���@q!�}�e��rd��	���8/�XW��͠�7Y��Ӂ.�ļ��ص	����.�*��݅����T��j����H�f���1	��{@#ń��]�!e1��ߢ�z��@�X����:lf�� 7�W��42y��ϰ8��S�!c�d�r��D��ŞM�d����\Rf�Ĩ�X�Q���;5d`��b���f�1�'�!7��9wa��yd�͜�NYhos.&�1mkS�#�P{*�Y1�Μ&Ȓ�b�w� Iai�ѣ��J5gџ�ӫ+{!�95�Ғ���i_����~2�sT���=D
&��0K�h��U`6�,q����h;s�0���I��������tyI@�KǴ����6�貆d�j�A�ï�90x[��/�L��~������F3V�0PʦN; o����,�=X�,%g������٘���ye�"8����&-�;�~�d?u��a�Ϧ]����`1)��`��$D� �P������v�C��y)��9��s������l�w`; �-\%���Y=�9&pM4����*F�j8��aLStrH0;���xs��|V�ct4?o@�2����>��f-)�����SAJw��qCI�Bh�n�t�/dapRd>��"9}.�j��ش��XՓ��{F��)6%�k��)�(�0��i������񈼞,����'#�G^�ڙh�Lг�"����o��l�6
y�=�ѕ��lMv��ǵm�ӵ��rl�&�1�f���w`U��}:�FC(�Mn�İ��~UNc�M.4{Xj���g ��h�%�����1�b���A��ԉ0.�fQ�x$/ۺ��A��T\�K�����S� �-�;��|�_	�������sK���i��g�D��L\S6%e)j}^NCK�U!�٘B�[:�F~mw&?�ٖ=D0�1t���!g�/:��#/i@|�ׄ{�c�D��A೦��<�Qƨ��b*OɮˤŬܶ&������AR��U9P�5ʨ\���ukY5k�+�:®9�T�����h�A8%T�a%�"�_ָ��R�����tH7�w�3�����1�|�]�4x�u��˳�2��Y�Qq�j2�r�6=��B�uJ$d�4f��4����)z��2&%|2�SF�U�Ť%��uT��4%��'�&*�j����R�{q2�A��=q��3�P�O�p�@<:Ɉ��9=PVeqb�Xl ���$+l��d�����s�z���?�2#!��IQ2i�-n]ؤv)҈d��`;��#mǡyX�k�'Y#UyaTP�d���F�K��a�s?��b9�Fb�Cy�@	��>�Lg��P6*z����6/�1��������(��2�,�&������1k��m�b�AY/�6z�(����z���.�� {��'����ϷK����#13zj�(���զ�!��A2;e�":m��R���vT����$�3cxU��Is�F(�VFC3��A�h����j�ߗ�Q]]-�a7Z[��,��ؑ�!��a��@	�Fl�Ps��S���TS&
a@ �Q#̡{��TS><3��3*�I���ELIs$�E�����6��`@����Ǎ����5ZZ��
EEt&�$�K}SL)�'&ap.iL}��)C��V��{�q��gj(��%>+?/[f��1����O^�L����6�c�8ÇԢ��A6�ɻ��rX�b܁��X�!E� T��iYّK�Pۅ3/�S~�Ҳr���ڛ�RU(L�J#Dcd�# �CA�^p��ړ�إ�ͅW�ƶ��a=��i��^ҩsQ�4�,?\�),�)��x#-����ѪE��q�!�c�葈r�@�K rJ<\SK���J��Phy�^4cxxznr�Y�ʋ�c ��!fˎ�-xlט�}�E��A�pw.�x����"�Ooc�.�R�،忮�XΑW�N�?q$��f�6|b�V��-3�-�Z}��Z����!��z�wb�8l�ڞ���	<Do)q>G���ᔋI$�r��4`1w����#��P�_/�数G5n��:#�|{95�~�{@~V����g��!�P��lV��ؗ����D�R��z��K��t�8�CQ�s�;�˾�WVb��ߩ'��w?�^�*�Y�IӲ -��1���N��쥥���lǈ�F�u�,��wljhV�o�_�������ܣ��)G���vMx�3���<�`?�`<�������Wn��J�m��g���+Ʀ]s$QAi��9`߉X����h����Dfq�<P�k���G��3i�x�Jt{�̑S1��/�]R�Ҥ6�)�1HT��Ӟ�U�_-���}%�roo�V���r1�y�m��2B�����Q��ű6̜~2F֖)2-V���A۵�>���/�H�����-"{�����R�aݟk1~���q1���}���c���y��4�c���LY�������;�r�ل��:%�m�yga�GK`�wR`֖����.�v�Uxp���-i�WO�﯈X�3O=��#p��$�7���C+�p��S����p�}
�5���|$�"���3N/�)��G�Do8�d(��
���ş/Մk��%󞜂٠��w������Ҧ�nUbI;�k�aP<e��1�\�$^��WNC�>9�D�:P� *
+u���S���x�d�Y�c�s�j�O9�A��L6t��8��CQ�kCY*A,$�_�*�g	�p��}PWߠ��+���Z�P�̲3Ԅ���ۅ���QS(���KB����H��\�S�������m�yW^v�;Z���5u�ˁ��2l޼YT�/������K+��yyY=��ٽ���7�T.3������ء�藽����p�cO���D���a+"�zz�#=#jʐK��'�B���
Ƈ%i����A���v�Ԧ�wrF�Ŧ�L
'�z���!M�8:$d���3 �<,@	���þ��s9�Ճ3�?N����-(- �s�1�.X͛~����+�;�A0�"�*Q�p��8{�ihoځ�G.�[�� 99��.`���W]�{Y�����$�\�::2n�v�\x�e��}�s'd~������;ճh͓E�h�lQ]:s�����������F:�wH���^$F�Cx>#?�j����Y��暹ʖ����GF����̺��.���<�p�(-�F.n�5��{�;���w#-g�v�h���hmlBUq�:�l	]�q�ɰ���J���-��ա���p;.�y.��=�5eB��Aq����:|�(�;��')1SEE��ƃ�A�wu"&a���z���m�����0"�醫/EH�C>�5#zU�;�M�r�&�8}x������QU(��γ��jn�՗^(зC��@3�_��.���$c�l��DOo�RէT�У*Q	A��x�l��(�$PVT*�+��[�ḓO�򟿂��u�\���>�5{Ū�w�orā�1���dX�׊�D�!�)��4��^�u�a�p�wH�
�����pMi!��۵[ �C׏*��v6a���PW�eY���P.�w�nA@�8���+��p��P�N�{Q5�h��a�	){�P�����C0������/�+-�^��b�P.�q,��>�,�������-�#(,(D����f<t�\<���0�;$�ؓ��ô�GcRu������)V��Jˍ���D��0~$�Z�Y�6��)��)g���9	&	��ሲ|��B�mm��Qcм}+���ܷ�_x�Z��6�����w��]�ހ~���b�'N�_}�-���B��L�1���~�9�b<��kpx�$�J�/�^��R8r�\�>�k�~��=����M��/��7��R���Ͻ��E�r�̚��7�vANy&�Gx���.�P�)�&"��� ��o��LֱZ�JFèL4��� �S�x	�p֬�Ѿ�WB&�;�Ϛ	�)�}'���}^x���yb��3�Wq內�Uَ�.�Ǖ�t���[�^�����u�H���O⒫�TV"km7�][���<��f61���3�שq�_:�a|��ny�9*'���uw/V�X&]<DefL?UD�t�y8~\�R��2r1X�>|���ز���/xO,YT+%Gy�j�R�0X��������be�U��^�1(ErJ��⭅�����p�?.��1m�͎�%�z�z�:�@��뮜�3qY��{�{�~;�ש�,$�!�2	�%�ӎ;���@� B�8\�p�7Y���)�M .��#�>�X���f��p)n�{�2���v���������0��e�Ϩar��0 0���
�����!�s�Qb48���z��gM�+���iS�����h���z�r��P/��0�3NBI֊��bT����MM�P��y+g^4C�L�x?F�3ϻEb��$��a쇣�O=R� �aÇi��:��c��,)@gG/ʇ����~�V��a<�?y�;�Mv��a��s�p�7�%p�ZL�K�̠�jn��	4�`R�5��~�$A�P������VAL�3an��s/���-��������7����"{]6z��8m�Q����ų�8~<61���(���CO�\|����Ϝ�b�*le�D]K�L���	��ss���0��w��/ԲvW[���/��B\qͽ�u	Em�̵������M�\����ܩ���0���4����4��.�n1^s�:E%>}����b����ܥm�}=������s���k����}��$k���t8N={�|Jj�*����U7އ�3_{J&H8\^Z���]&���?�j؜Y�?��~���
m�g|@RdV��|�y<��honĝ��Ͼ���������gIH�-c"μ�
���:X�0�tؓ�=�^x�qX�on���V�����j]G#�nx��v\���6[v
f�F����L8FNǪ�7৕k�by �����i��c1moA-a�=i<V�� �ܣ#Յ��hllqy��G�b��p����DD��s�y�n�F΢�)�(� �@�z�x�<��N����At%�{ʦ�I+.�i	)n��2�dQ��J��yg���ʋ,?�-�+�FaE�y��?1�a��DV��7��;oF���j�ur���.Ñ�vv�'2a���!��A$-N����o	ܜ�"/�&=�oKh�%���Ws4=�-,����y���0�$����}�G�I��[�Q?~/BQcr�y� e�f��_v�m�"��Șȭ��k6o���W�DW�����.�;�3�YC�U�U9d^|g�lo�]K�$,�mk3�޵8�詚��HB�G�yxɭB�g��蕵���49l��,g���aʾ�/и��P�~|�L{L���s7z��q��W�Q���1	�T�ε[v`��Q(�Y�)�w��MbX���TUh9��	��_���Lb{��v&~ch�0����䙉ʥe%&g��K�[�D/�b��w`0%�΄4A3� ��;��+\t�����y�f=G)	���Ə��9'����R�c09�p��������G�����}L�NOR��d�j�T���;�\��fN�0|��8|��E��ǣ$X���rl��2��h����ar�Tyo0M*A��p�I��+2K(���#Q���Ҧ�*��v������b�J�{�Espʺ�X�`��'�	�[�6��ڒf�����/��0/�!���YZ�ړ��O*W���x���j���� ����5��'�n��|f	��Р��<���~��.;b���PW�@;�셴}����X�t}�}ho놫ʯ9*��.t����މ�ؠ</�Y�>Yw
�i[#�2�X�&���4S��?��^r|��r�2���N���eXދ�Nf�c���e3����-�d�>��қ�OkVy������W�ʋ�4f������$�h�b+J��G_�%O�b��߄|UΊ��v�;u��,��-}����l��F�o�KH����%�I9��Z�w�B���j���g2�[8�C����/��}$#5[c/Z�:�p1,J,N�/�נd���29d?��y����)q6QMDS��_\.c&��|�JS��"gp�����;�\NQ�Og>X�d��j7�>��A���)��8�v��$&%�)$�����"�)e�r[sRc�ߖ-[1m���,GU�2����P�SU��o���"�K��9�N�V�!��[!F}��iY-pZ�j$B��o��
Oa@Bd�ʙ���,��M�f,�a3�@R6j���9�h�lt^�CU�8��镐4������%غ�N�©�Dو�aZ2O������r�����ήe%KP�M��'�LW�f�g�T���/pO�J��\�Gj����G�D<�_ɚy<V�
��>�I"���r��;Ki���j�����]IwRTM��N4<.��4>���Zy��3Zڳ�mJ��r=_Mu���7�~��}r0�������.m&�ƍ�-v���u�y�kU��EUm�Lr ��o�֭�K�lK�yt1d��t]gg�!f�5��3*C@c�g�*�u
�h��(��tŪ��A=��py�JDd9M*d��䴏c�IEYBU*��dn�M���O.zX������$Y�R���<�n�j����I�A���Ŗ���b�P�����l��w j��٪�"� $���� }1�3�$J�d"f����s����٥�����M���,�m�!ve�&+�C� �~A)C�ʴ;����1������1�I2g�y}C H�1��5��=]�2 B�4��X�56`w�.(�D�l(�S�Hޱ�Ч3|�~YOδ�Q\1�䠟��uii	�bEIHÄ'�;��:�RAa,�aM���ƼM�[�ϊ�|v��Pƃ��u�n(�y�N��Զ�j���l��S��F��!Țƨ�$�w�Tf��MY%�����B^|�$+�QEb�<!�F%b	�<AE�oQ(��%���{k��W���.��)(0��'$���]�].��}O��~�c&}����>�
�75k%*Mb�TV��$q9l4R��v�HH	�j�!�%�TT��1���bw�@69 	�d��Pk#eBL.=����R�9ZAfs=.�da(Y��H��Z6ͦ���"��e$����$�M*0ZV��V"���WoH��Cڬ6��T���!K��ݗ�9ɼ].�S����5M]��ȑ��pZKF�x�hƁ1N�x�m�vC�N�?�)^�"�p����4����/S,��K�Z���'r��>Y،6�T	\��y��y�W��UQ��`!�ڣ����j��l�4��)1�	�>�e���v>�P�+��ÑվJ6�5� �0�Fޚ�`J%4���nMi˸�	�(�ވ�d�ݫ��ɥh���
�X��*�#��A�ṔSI{K��ѩ$�b���s;��#��`Sv\�tw����ֆ�Z)�ͭ�q���0z��MS���r���\'Q�G�a��{����!��eAEM�6��׃(�)F�*���Հ8�,n��W�DlknC(�Vb�w�`hm�s�8B�?���I� R&D#I�XI�{�Yx�W�+���a��dc;x�(1�vt���
i/R��'r�Y����$���)h�Y�?��}f9�>1_�8���NA����L��dM[ZZ��T����8l��h��	}m��i��N�I��qԌ��;u��w@����IcƬ��mJ⌓�ۋ�j�0�Ug��7_=G�[J�W%��P��I:���ug�|��va��6	C�ؽ�7]�r�Zww���}�eS�cd,ʖ|��G*����d��b6�`Y��w%�s�}Zڪ�MmnnV�.�@���:A�W�dS<^B���2{qо�R�5�6�@��q�	A
���Wc̘1���)1���Q<b�\t�6K)#�\�!U��j�������69�Lk6�Ȉ!m�e �Dca����>q�4ly��4�ɡ06���KϞ��8�n�6��?�������Ȓ�bX���{�ݒ��N�0#GEww�r\x}�0�<2�1,��"TW>ٌ߮�ɯ�ڌ�����V``�v		|*� W�h�a#�<)�)?pܑa�?�)�S��	bʱϘ�r9�Z�]�~�:��
Y��Є)C
���U�1�,|��/�ZI��p��=�ʲ�>+ߝ�jt���KTj�����Ι��Y��#a^nK
eA7&���D ��xa�V;墧S�O�����ϲ�($Z�IPVǜ.	!�C������(�ʁ��Ҭݭ��a�<���#�',�^ySBM��v�L1G�qάt=	�)����+P��Sj��ˡ�r0֏SN���֩�� �bQ%T�8�Z��ذ��R7��9+u<��Ԡ�nΝ~:�X�^���I!u��.:�L	3�e-���u/�����P"ݽ�|Fݟ��S�_|�R�Wi�WD�>�<;�*�ʌn	�@��MN����H8[ļ�n�7_|�>i�6T���5�M���"l��O�_D�9�l��wLs�$�1t8��s>��3�
"9���p���"��H蚂��c�â%�	/�� ĵ���15˃����s8�zɩðq�Fz$v5l��3���?Be����nڅ��ESm�	D�e�r�,��S�a�V��.�c������'b]�%%��jW3�:o:�v5�����_b*1l��AlK��G_|s��u�p��#���k�YmZ����?�FK���BY�\,n0<�}�f�A�01%��K/������%%����a�X^L#�*�{,Q�0ޒ�˖�~lh�Kč����xfO��J�B�P[\�c������X(����iYzo"�>�GM=��.̻�,,\��w6��'r�q��{�F9P���E�
GƦ^%���g���w݊��`dM�n���[�L2i�8L;L��.��,������pzj���32a��E����L<�Գ�J���<v�~��8���/�P.,g!��8��\�_�m�~{���W��kgc���&m�!bt�aBŷ��Z,Z�&�O�a�D������Λ�O��~�������{L֪C&��r���;���_�]P������؍1#��u��?qǜ����QAL 21���O7�9�w�{�@����Y%���E̐}�2���NmM��ƌ�AW{�:��������!iM�?�W_:�r���W��k���%:�PS6D��,��._^z�u8|�L�1MX��G���#�FF�>�8���wz�ikz�C��#����{�<MbH��.:p�����?/��ٯ�oS� .h!H
��AD��2���-���/�a�͐N��f+�y4i,��b\l8�Ô3����%�qȹ��2�4�Rl�\��@���ƠH Pc���G�zF&���b6Ƕ��X���R�Do�;�٠ V%��lASS
�ʱ��:t�	�qs ��O,a�������L�.�l,���>>�bR`)v���v��|��P�Ru7��ۼX���8b�A�65��:��g����U_/�#��X~֋(���|�}�y
y��.��v��^Ay���34��8����QQ=���v�1��9�r��_0㔓䢬�-7\��ͻ��ݏ��S���Uo�<g�h�NX$��F,{9[;�] �ı#���	2�䂳Ѳ�]����!�߷4���jxR[�M��n���{����GR���_��g��x=5{��Jx��bL�ej0��4��8���0����։�ؖy���3#��y�6���d֎_~[���	O�K2�!�l��6A y�!�퐟+v��}�ku�y+���\>|��4��r�ٿ,�V���O����\�?W~�QeV�x��:�W�m����v8�i-x��TV#���%�2�i.��kL?�48d]w�# 0i4�B������T���}O%:)R�R?�"�q/�cu����P�c���bX��Uڸ�^� <w�~ߤ<0�����j�^iy�������J�t�o�p�c�/����ڌH�Y9d8���.]CFq:,�@<Gw�^�#�M;.	�v�ߤ9�E�RiQ(d�zï�g�����fY�ܲ#�N�����ӏ��`<
� a/��G��cxM�����X�ɗ��fՇg����R,Y��;
�nx0�mo�1�FC	H�����rr@�1�2��m}���E�K�,��*�,���L�P�ᇕ���;0a�P��>Է6�C��4;W��l����k*Pg4��.���K�ƕ_(�m7�w5`��Y�%��b�����o�<U��H�\�,i�x1�DA���&�iݱ%�2��~�F����b�~�2u���H=�}<m��/~�駝�
X=m��¿gc���_�f�IX���Y�)�>H�苯1���Q��	STB=D���iǠ�5�6��"G�>z�R��4;X�N/~^󧎰��x12�hشI{;�����X؎ϗ��K#U���f�4��P���"�t�M"��Z���4��b�����j�����5?��(�]P����s.<O�i?����
�%�H�����^Aa��0UZVW8�'����[�<^��0�w*/+9D}�
�]���:`w4L��bvĲ�B���j(��:��:l�s��Vtut�{(U]�/��9&&��͞�lL.�G�Ӓ/����ӮI&�9�Y������㯿AL���:jVFw�PVR=���%�\t�R:�Li����C[Y��=~��}0�b;=��ل�j	^x�m�s�튮�b��97ӟB@P�U���O<�����#dSʨ�f��&���)���*\|޹���g�fU6!"����+�i[�^x�萤*��4_VR3�z�I̻�J�sFC#VT�1�:A�-�X��<�^̳��)'�9�]��� /�dj�K�����t��jX��>�s�}d��D�r1^��;�}ExK��Y���FDf��B7���9߭�]% ǎ�կ�%PRld�W��;V��>��,G�uJ5���^(�#�><��[8��㕍�P,~�c�n���c��-���F���ҋb( 묬l��6nCg� &O#��@ii� �^��>���7�$4����Y��#��*�fu����0rXJ���<*|�д;ۺ�#D)�3��bM�f��"��HA��A��7�Ҡ�]mjLȚ�ھݡ���d�ݩc�9EeL���Sh�n�L�8YB�]����5���G,�OP�!8��p&�t���N��4��=�.W61����R��<�:���thД���ޤL�6��y_|�}A��ɥ#C���D������Z y<�*�����πA���a��N��)A�}��ա�[&[#�����&E�����(�rWR����{����B5V�eZ�$�[���i:[�������� M���Ձ�o�Ζv��M�Z�͂�
�i�6�i(��|v^8M�C�::)�-~�o˥O�{2��s�ή���耗�ј�Q4)׶��
����0f$�nى{�Ę��u�4,�F	U�8�opT�t���%JW�l���O.��e�ِ/�Θ�|�ɍWps�S$�
 1��3��w>��^a�����ɺp�������6���]�e� �E�\6��,�Ig�6Mr�X�����33�Nf(6�Xăy���Ƅ�)O�<�,M���	�^�u�VH�QjΈ���W(���	O��!/��Ub�z��>��dR�X�O�2�TȈS�V2�f�(Λ���g)�&���7��~�Sbθ��F�K���i�?� �ӱv��s
X�*[�ug��?��D:�]tv�_If���?�����*SV�~�5�W6.���!��ap�BgoLF�:�'p���I��I��65��$�
���<~�a��NX�7��e�F�O��D}G�1��
K��G��*Y۔��`6�E1�˯�rt����a	���u���iרu��r@����0��)��"3�,��J�s`����g<�6���&.��j]	^@Y�����1�?uu۵D2���[�m-{9�.�F�(P�2�|�Ϡ7�dq�lq�Mj�uh�b7�JM�"p.�b��2�fS��jѸ9�"Ҭ�<K������l~ RY�Ām�s�e�6exr�0<geʤt�T}~xR�JY�wB���_ɚ���*��O��6;�e�z�ւ=�DU&kJ�Ǭz9Vx�lA�A�,���y
U�K�]��g5?��0T�u]�{@�������S"��euU3���Ua�,ZRW�9yQ��*;���:�1^�����M�P#hOJ&������iTttژ1>C��9��z�����@�-׶��bX��Y�h���ZG�"��l���t�un�����})�y/��|^ :>�Ʋ�ckS��"��Ăi�����a�k�R:k1������	�rd����d����Ã��&s�r��|)��ANs�06��tkӆu�!4.�C�L���$��r8,��a�?���4P�g]Wn�/�Xs��=�y@�v��YeG�4��ޕ�9S&ox2z����I�7�,��RD���1��|&�C�c���r�26�1���"T3��h�܃�����j�j�e�_F#F�Y~�1̸X)�y�JC<��쬱��*����_�2�G�� ��=c�s�A��ܞ�ϓ�!5R�wq���Q�c�Yi$���M�u��)tU2zw4B�wR��<���[شڴ���?25̃���eK��y��I�����VZ�٠d�2����E6����9.�)���e)\{�l�Ġ��R�9�+���J�xdY"���sa� �³��!�㸰,�6Bq�I�1�:��l��zMLJ��^>�BH�V�ȀzY�p�m:	�SBc=�$��ò���8AƈyN9-���R���A�?��D�;���J�U��j��ƢZp�Sʂ'��(yI��(���SȲg� b�Avn�"������\l���9�3<_T6�n��SNH�U��LQvyV��|�Kk6ɴ�����B�_D.N"��q�Tʸ0d<#τ��Z��l ]�sյj�d���1��nUf6v�:��aR�hU���9�΀+�I�gp�IE���^^�Bi�*u:�DL�&�T��t�+��ߣLW�r�8�ap�R>��� 9c��˦�:1bp
��]���JF�s�cqA{�x���3yHo�'0i4H(�~U���I%��Y����C_�&�)���3ر�΄�_{�S~������Ĺ�ք�{��¦,m���gY�A͹���abѐ�����4�\�,�+I��?:�����p�r_)t�P���Z{�|nC����KE�<���mNG������s߄#��%t�z�J0M�`�woljV�Ik�-���CeV`jL6?~�m+J*���!� �M�R��V+U�B;�P/&O��hz(f�m����/��֦|�H��xrQsf�z��M�0�F5��b,��a�+T]�<�:����Ye��9ډ1#k0e�aH��H�B�z";�nS3I��nv�of���v�0Y�� �q���kq�I���^�h*��W�Ǻ�;�s�T��I)��$ĉ�g�&"1�8���P"��q'Ə���xmx��P6lR<�T�d�(6)���ܹ��:W.LVG�y�yfAN/����J��;90��+����l̠sw'�8����T�"�=��\��͛�ê_�,�CD��DD�Ia�1�p7?GO=�~m����#"F�Ͽ�5Xh��ё͉;��Cc��,��I�[������k�#%1�Gb�/���1�J��RH�Qa������W_|��(%�l�@������Y\��ě����j1��� j�+12mq1�r�����u�t��w�ܠ��4r� ��<��eH�yjb�&;)�9�&ӱ~\z���T4I�^���>A��X��W�)�L�I%�������ц�>�#���鳣/���\6�{�|T���,�D��l\�R�$�2m���-^��g�t����j��{��a���b�>�_&˳��;��L��1���e������i�����z�aT�-�lL��;K4jhnގg<[�C�uJ�+��E�+�����uƙ' L\��� ��~����Y��R6\�'�Z�<�g9�l�ӏ>�]��*��Y�>��������GD%cC��+�n$v�ŕ�g���dS�l�9����#'��'����F�/��ٔ�x�Y_�p�;	���H��,��Ρ�̫�����p�W�hG�E����FZ�ɣ���`���@P�0�OA�QÆ�@c[��"G�0jN1�l�noż�"�E'V���?Ы�F�r�n��Z<��T�WrW:4�� ��x������y� 3@�+�;�0q�x�ni�ŵW]��x��
#T"�$�$�|e>�x�4T�ɻ��*[TH��#�(��������u�qK�NN�)��c)A�Ua�>{+K�sڻ�Q)�*,��=�q�iZ��2�H\�;�j�IJ�d�-�����P�n����nt��[<{mn��Y����u9��A7�;p��1����u�1����ކʪ}��5e��Q�c�ʵ�\��s�S0�Y%�� �C�?=�ʳ�<���bA��p߼[q�-��|�0�)�ZʤeWΒ�b��GyI)ښ���staTH��Y�����{Q.�U���(�!��.�ɲq�/���ݝ`krh &�݆�|�o�#GO��vk��,V����޳̻Q�?j�3^�ĺ;;�I��.�C^V���i�Y�IQ�j���ĳ��/Ϟ@Uu��,mxP[Q��������a����+��ip���F���V<p��(��i������p1IG�ԃ�kD�kww?*)&lgw��MQ��S��G��H�U�pi��rica� ���PY��Q�l>�ݓ�6ӏ?�}�����V�+�e���[1�3��8�J���P;��� *V������2J��!錨���){c�xj�1S	eS�݁�N��t幘�����8|D��Ҝ�)��X����*�C��Q!_Q��6KD�p��S���_�vs\��������!�khk�*�����J�X�+�.9Dnq�-�q����yA��*�z���v�ۯ��إ��e5���zWG�V�\L�nۈ��Q��Y��!T�)�����#�ʥ���M��q���
�3�	$-)���C��~��Z��3F�.�T$��N����� %Ϊ8	�$�I���K�@5���ϼ����i[�8�l�����
yF+��%�rص����׹W�>_�}av�RĘ�{��=����wf4�%&|� ����UlUq&�����u�AȂ�zz:1�� ��8;(�Eqi�\��yy���DdOi��y��j��n�a��C��sf]��1
�c�����pU�����I�{�uW��Ǟ�͉���k�ZE�zq�	�Ț;��N>o<�:Z[wc��!�k�H	���(��3�����!�ذ+5:У���<rv	�2f�?>��հ��ç��C_o��F<��h��FA��s��u�V�}�M�h�ia̎~D��*)1e:�JH�ϹW������JEkj�����K�N������ڕ+�i�f	���᐀e1�99Pŕl�҈���2YImM�Q#�r�����U�<���P�]��嗜/�e�&����C�(����q#�j�����9/��И�u2��T�8Zn�èQ�2}���\�_��T�a�ӔFnxE1��r��~�@C�,vd
�?z�<IմYt�����U��؄�`�w,(���֦t��yQB��8-��A:��c�!�(���/�`��M�$��c��� ^�c�Rf��a��$b��5��d����.xE�ry9`
�o/��!ͷ�8�$|��r��^-o�����@�x���j��;z
-�mʆ>^µ�O>Ve:[�q�E�♗��RFs"����K
��Q6dz�y��yei���L����X��!�N�KQ�k�0��tp.�+f]�m;1j��x��f�z����~��f`w�V1�\|��X�ŷ�s�6�0%g���O[��;����"�����\8�hX�?�4��p�Α�#�,��S$�H��5{���/���M���.�s�v&�:���{7�wk���R<��*?Q3l4�{�}1,[�B[����7�J�Ǒ�p��{7n��AK�5�L��d�.���e�~�m,_�Zg<��c�Źg�}'�A��{�w=����(���cGa�{����v�LmcNk��:X���>{��qWΞ��>� g�J�q��C*2���8e�%(��D2�F[_����~߈��}r�^2w>��n�NӦ�q\z�lx�(�Lj����s���8肀5�<vϭ��{����]�ş}kd�dhǍ�PBB�@	f�>]Ѡ�9�lo��n��
\��ٲ��z_�@�%_��3N>�0^{C�J���z�$>����){	��lp��_�����B�y�*^�������m8���x��9�
8�(�=U.Uss���X���;v��(��.�H{�<�����*��.�ЮD�x�DdPE���rr�J��`��m�R�7����O��;o� ?MP����/�U�?&��b�J���K����� �d�H�d�r�yX>���^�C���Pb4���Uvr2aO�� �1����
�s�9|��2��4�)	�UU�q("�:f�M����x�ꑸ����x
�+(݆҄�6�}�D.�Y,�k;��;K���uH

�)� ҹ�CG��=�8IwMD㲆���_.���Xir�j���])Fm�SY���f�`!n�����WYn$YŨ��рO�~�c�GsV�&��\�J�`2�MŘ�Z���/���
.q8����Q��_2S|ݠ��tG�6�X��>1�#5�2q�4�b�<Z���<��Ë�p���R�Q`����SϽ�*��`�VRY�;z�:
��Ꞅ!�Zzp��O��/78"�I� Zb20.�9tH5:�}��;ll�wQP��=�����_��1r$
��vu`��4v��OLP���Ir�5q"N<�R��t���������FJ�F� yA���v��۱�8��W݁*1~)�ʙg����[���o`�1C%�6�g{oX�3&Nc��F����ĉ��A�b��=��������O�F9>�C����X�u�T²��h5c'b֌Yr���;/�V&�⩧^�/-���u[�a{5�*�&u>�b)N>�D��$�����^i[e�+x��>ĳQ����O���W.��D�ž����݃H�V}�I�mŚ].	z�+p��/���ި!E@Ά+6�����������3l�ׁ�@�ZY���'��waG[��0��
�/�����⺹�a�$�����V���D-��)q��o?oi��cx8�e3�b��z�v(�n�=��7c�	�z[6]y���WT�f:� ��p��#9����T�>U�2Y�4�X(���/9*-���.G��*,����@FJ��A���Td��{ =���d�����Y	ƶ�li�D���-u8hl�zbo�O�،��ˀ��Q�)�aW\�eZz��a#��͹��JJp�#��9U�g�8k��'J9q�lT�ġ�e���dBf444��,�n���2��;5W�Ib��3I�򷍂f�Z%�>�?�ܰs�������DS�N5��*y��迉��[%������`Bg[��"%{�\�H�\�Z��B��ʜ��D%L���H�l�f��p'������b����^(y�Q����QYH��{<�r�]LcP.5sѬ�(Y�na͟��ߘ��w6M�;䰐*"(���z�w��2�O������dJ���>�Ee�[�/G����TJ�fc.�cۼq��v���lm��癏1��(OIX�4g���)�p�I���[���jUM�s*��S+�LԋQ�*E����+qm.�����	���@8�/m��I�s�!4�cȨ�X��2���,��ಲ?@�&�T��i�2/r��uWW�z3j�6nܡ�d�x�a�RF�w��v�V�F�Iֈ|>=}hpP-�K�]�� :�-)�5��He!YOD���>�?�J�$�O�b��wuvcԨQr�Z�f����Ґ
��I���d�ʋ���Bb�XM�`U��N��q��{z�9|	i,�s)8�m�d��Ȧ�ذ�O��V%���T}������^w���,]AA,(6� ��P{�h4&&�4K��]�"����{W�^��f����s��7��vw�y���s�9f��g3"��a������;��:�/�|��úq�V{,T�b�<��mC�@F$ek~@�߬�C�>��>����!�۾�ɕ�{���q=*|�$�/{?�ȲY��[t���OP}��`*Tx�u���;7��bdB��5U}L�˗?�a�����ҵe[ɔYfL�e*�G@1Q�8]�ƣ
Y�j��Q��S�$���i�+\��L����ڱ��
cN�߰#�A.�
Ի�H�"���!��ţ��5>� �&E�XB��&��k��NO��jm�:1tO��]b�]r3=��ym��*J��P-��r��P�Ԁ��ł\p�<;ud�HD�.!�ve��q~�7�D�XXyc���S	59œ���,�H�@zH�x<���V	s�W�Ԧ�K����N���k�Ѝ��+�w&cU1��>#����B�F*�^L�x0&Q�f,���6�h��^V�\Jo��c��uyU�����l������.�h���/��e�R7����bm�l�rRʎ�uT�&y���<�:���8h�s�&'��'�6�o��$�*���<D�0�S��B��,BR��L��%꺐�$����Q�"�x��,���E>�@Ie�Q��,�iC�H�J	?R�(Zk��X6.�%{�r�v	��v�n�=��X� �E����FC�!�	���!m���uS!�-�U^T8r��9l�4�k�O��;"7UX���j�!�1X*��aϣf�r2�$$���A���^�yuj�\6Mv���H��T&�c5�T�ON�8��f�i���jW<.^w�L�2�RP���BFW�3+k�FY���ߘ�6� ��LY�^�;�#�4bC�4"�!�g��^[/�!���n�0�E�2|S��!����"�r)�>D��-��9�g���`���̋ѰY�(����6{X͒0e�h%��ϰ�G2$9��\��c�Ah^�TV4#�UŘҲ�il��^B3_����eZ�	>����~�E{�8!�hC� ��*�k]����'����A�S��Ì �beM&����MC,�?=bH X����AS���~�xӠ��XI$��	�)�!���Ԭ �e���C��s5���;���K��f�Q�MpHT�6�񭭰66����N�&���<�>;"�1�>ʃ�hZ2��Y�d�-)G�G�90�`y���$�"��I�Ԃu�dJf�.�K�x�TF���3f:zYJ�J��1<�x@�ܯ�� 1ث�5~z��j����Q��/��zAF�9�
� �'6ech�P-Gw.?a�1sb)H����,�O?U ���~���0��-�1e�xɤf�	�!��B}�p@.#��ASF��ݙ1deJ���ߓ�,>�IwhSZA����C8`��ᔰ�����g��Q��J�@���2Q�6n��s@�wU�5HǇ��|���=Hp���1��3c��IJ�FX�R*{3��y�vw!�T����������r�B<��Mh�f5��*	�D��"'�ס#�;vv���ǿ{UU�r��Ġ�Q'���"բy�r�ĨrQP�F�:ƌ{�ՏV��v�r���N�%a��M&4����
^6����Cik�AO8����$��(&#8p�}��2/�n��W=T��E�|E%E�0a8��/�_v=�������f6��3��1x�k`�gDU��YR�3"aPd����M�şn�G�W��[G*�:wb��'iSc8��;TRA0�rmyx�H�9�\lz�)��r�$#�<l���>���)�����5"����b\c����>���n04؅��*�F�V�PGW��#�:7�ә1y��.�8��C�b�*Ğ"q�یP�0���<�������Qc%dR2�t1�}��K<%��V�s��ڈC��OҪ��2�"�jkC�����KM6"�]^��}�a�&�6n���2P��	@~�1y���=)|���hji� ���aw�Ac���K�lh6��l��͛%>� N�q:�^��l"	R)@lGeU%?t��&À[b��]���ve��_�m��L�ߜ��{��#A/q�feGl��6Llo�I�~�}��7:N��K��'�8��k���B���3r�rڗ�&nԩ��P�f�<��Asi��Z�^�X���P�p�9X��U�|�	t�a9��9r@JZ�f�m�m�nl��|[�o��&�8����1g�=�͆Ny�j+kaI�q��h��K�!��/{|)|���İx����:KKi�G��Y��寽�aC��'�tdD�����s�:�P�r�q��7^#+��	5����8VyO$�E��c����z�b<�l���*%��r�YX��s��v�찉A>��1~T��N�X�����i��3����G;C�(N;n>>��l��)HƮ��3�����b��WB8>��'��3:r+��2zV��.?h�~�O��'�����$ޞ9��9M���Ј2|9<��p�֑�Wη?�n^|�&�S�~��/7��GGG�N���g�yU���1YۊV�J_����XR���W��+�e5a������'�H���y���r���\���֌���q�5�ۉ�O���|�����Z_���@��U���e����x�8Ʊ�Ïq��}P,h�O7^��]���^��c�=�d��
��~Xo��l|��h�l���NL�6͜����vlݎ�XwWE������p�Q���G���L�7��$`Ӗ�Y{ϖ�������,}a[Fk=�ȏ��/���!��bRK{����[w 0c��du����&�}�#��5�b�n��Ͽ�&�2[<@;��q��C�es���Xf/��lHo��pS�Тz�m���bNg�(�s���ՋR��R##�ʏ��@u`��.�j��Ֆ�8��{�}���_}�!�=v.���UIܟ�V�X���x�"�rP�\��|V�����ys�*��{&�7	���m7\��m�%,��A��1���#F��Ecs+"y��O�֨�Ǟ^��9m5��k�T|�z80k���Q �nI.ȫ���rwj�@wR�=�̋8aޡ���S�m�.R=�HV�b� �������P��6-l����8�ȹ(
"�Ѽ�Ke��m���h�|%ܨlh���ޏJ�G�05/@�В�0��y��q�����f>���H��L)1����Ns^Hūő�7��O��'�_����9�s���HL�!;7!!爪�lچ��}������wf�i]G/,�oq�{a��/�,���(����v�%��jq���W��}:Hhs���	,y
��wul�C����'c�8���3��,�����C�ى�vQ�����>���7��U�����lP�,!��$!��'�TтG�zN"�jAc̷y�1-_��'����;���c���],!ZF�!sJ������ ȬQ��x�pcM}3�|������ǳ,����Q�6����ڶ1��;0w�ݍ�`L�x{��iy�^9,�_}��Z�����9��Ͽ�&����T_�x����us�ǋ^�FqY$�;�}
~�R�]s̏�%JȆ���G�)�<�z'�
��%�1ƃ|�cϾ�,9ΒX��x�_p����o$l����VLm���	�Hȥپm��/>��k���W�!���;�fgRV|��je��g��G�Zg�x�≣Ȅ���U��~RN�ۧ��&����1I����C��G>A���1�����,��nY��WU-�B�
e\k��ʺ|*����n�lz��CQ�gC�VT�:�Ef��(Xc�Ӫ�!�Gbc'v�w>�Qs���?`��Zͨ����t}��Va�>�ucw��g�Uo���_��tAmm�c��9�yC$~�$�Ǫ���O΁1�QT�AOi���so��N9VA_��!&��v;�DJq�P"�>�jZG����B��d����z���۸���i�je�WA�d@gY�۟֊S�C�Cc&�ԗ���	x�����Y�m����WTˊ9JV~��A�c1d1mY5�P�ǎ���
���E2S�R&����0�F�t�mry��e�]2��9�V,#�%O.Ņ瞩y�A>;;{$D�"g��Z9��+o���%�6�.��c�C���z��;���S0it3:�yZ�[�d''!��K"���_ߤ�L��I���	�]}�oɓ���Eb��12�k�%��Aj�����*$��U�Ң�	�ʺ6�p�q���֎�ȉs�8��!�<���Í7���"�����l��U~�۫>F@��x��d�\BNm�����O�S���$�MFB�ATV7`�x��^~Y<S� k�w9�u(�a]�$�{m%.�x����8p%1<c�A�1�|�}��^��9Pę����uj�^�y眉��.nm�Wsͣ����#MjV�N�N�ř5t�
�ߴU.���5:tg��`sK�5�k��"Ƈ��%�.iw�E�k��1�>�����Mk--m���<P����_���5r�
�1�,bJ#�R���_��A�ԣ��J�;�����˂�XF��Rrc����9�nD����fb$-�v�(��*|O�����7b395qX�~(�!U=τ�,Y*��|mGN��`��)��e�x�JCĚc��(��hv}�(<��+�Ѐ�g�<�k~٬�%d�Z�F<g}cy���+W+��mer	,yz9��w�:�H$�S���ୂ�v��q��v�����:�5��q�\A�ry��B/��~+���[��!s�z�5xVz�~�
^��Ѓx�3L�6-���Y�H�����x���+9/0���Ug���<z*���Ǟ¾��JAqԒ�ڒJ��?�r��Y�d��0:��J��T���8~�rm4б�id�0���BU�B�|��>��nS�	�w^%���ʺn�nl�ۣ=k7n����PU�UxC}���M�gq�^~-��>���~/�g>��Kե����g:�dc��l֡��׬Q�vo�R!QZ˄cړ4�lN��᭬�s�_�r�]K�F��D�a����V����U�[NGB	I(����?���%�m^�Д��p��-�C�C��C��X*$s�Lf��?*�H���n�k��%��&$���2�IKX<�� .��n�KX��nBT�T�I��!�K6m�'K�V���)�v@
�L��T׌����.~:�'!����a��"Q��e������^��>\/W�k��ЉW=��*e0�y�k��h�U�ni�"p��r�x��P,[.h�#>���	�̂N2T�w�1ݠ7(蘾9T�֎�z���W��v�W���g�(O�jH@>���+e6��E�̠�nIY��}
O���N�K�\�Iy@�v�B&m�*�&d c�(c�bś��$���#S�rJ�*4��K4ٰ��nI�_�'߭V�ʹ�7@V��!�Y�
�D�y��]l*�G�W��㥕(�3�̚�!�s{*�ϔ�y}�ɧt=8��$w\�S�Vk~Z�U��Aɬ�8��#F��+�Uk�i6tm5EO��;��[�~�a2�V���)㕐V�[j����P��j/����cE,!���߯� �FP�ɦS�*y!k�1�����ez��ΠQ���B(uSvti;>]2��>."kWx;�CeY��6������1d�HƖ���Y�^3�b��;���K"����ێ	��SH�\�K�&���g������X}�c@��t���Nɒj���.O͖�OC�Vl��q�(2]Yg=9�5��l��S�r>�U���rA,.��5��3Z��A�����fu�\�����0��P4�����|Jag�0���[�������W���%̈姺���f�Jm'�e,�08M�.�M,�Ϛ�0�0S���t
���}��EU�3�����9d��Y�`[�hJ�g�
)�2�5��'�?�P�
�*���2m!�FPPg�S����3��IKyU�=���U�B)���L�gƙ����y�͟�0�#𤕷)����:XL�����Ī/����0a^�Dj�\� �*��f%�!͝\&�C�����*������y����&�1n3���Az�I�Kj6�Y��ʕ'�+e�x�~9��͔�(.�l�6����|y�J�Đ8�8ɩ�/Y�"��L�NPn�N1��W�� rE�����\�
�J8�WA�2s��cS� U�ƛ%-#�1������	U����c[��Ŭ_�r���OU����dp8Z�_d)�ڛK�8!�Dkw$I<���d�r8~�bΗ���A�,[|����l�)��-�[H	G&'U��1nY�����,�F�/���烇�݉rQv�*A���~eR�^ЍQ�^���`L����T;Iw�>&��ǐI�i������iɶ���ԝȔ�K3��r ����Z���P�-�M��0����kPi�S�JTD.��l�J�bza��AAK�T�L%Mnq���鄱�e�F�Ɯ���{UR.�R�B	��]�I�K�6��ј���u���Ք+��A:�+Ck���)���˾>��dg��SP3C�uo�c� +���i��B�HIgt�z�sF�?q���.�B�ͮ���8v5r]��؛Li��%����Cl#<�����b~&D��,��P�� ?K>�\��0�g(���R$8����eA��xH���.	����io�F���މ�>!�q
J4�;pP�tH���S��۷BC3�Q�J�2�Y�U��x����
Gb��M�sQ�PMm� 㙵�g.�D0�tV�u����N��:�,~$F6AM&y�@O�! d�*d����`?�n�.O��Cci�Ҷ����cբ�N�Wb�|8*�٤Rp�|�Ms��rV��Z�`l�3Zd��H(�¾vC�p�J���C�0�d�t��#�A�1�DB�t¡UUנ`('��BY��l<�@c��_�(F��޾ACie/]�PU(�%�m�`蓊����A��x�V�,N�n�ءc�N��^]"q�vy	%v KZ<����*d���@�І	-:���Yfn��@W�v=�d�������GU0�G���������%��kO@�l��m������������rEb���ذu��$�{�=7X� �ɰsxL{;�L�{ސq�ڶ�+?�U�Mb�L���Xz��Q���~�	���ߘ�-�_�!Ϸv�:YW9[^�1(��)���M.���>�~�� �~	QA�q������֗��"(e�"j,5228�f������а^���z���ʫAA��(�`*\��9�U�X,��_�F�XL�}_�
��x��TH6���`2rt���#�;w�s��nW�����Z,y�YA����$`��F�	��Tr_{�{p��a�^S$$s#���y]KV��
�~�C��U.t�wJ��M�!�v6��\���p=�� 9<�U*��F��>�}�UX��������K2��e
xj��ڇo�4�LW( �����t�"���-[ᯮG\����^|�T�7+�4�E�wQ�%�b��c�蚕�ӃD2������_}�xT��W��.
�i�s9=��-�s<�Ybj�8&�?�߈/��Yh#�*[g^��6�a���}��ޑ`�����Ӌ��Z<���n\��fV~Β�|��{��{M���{��$��v "���E_��ߴ�K��l�h�?=�Y�6H��#f(��(u�A,���JTK]�^����4Vf���7\)��������ߣ�ާuw���w��y��շ�C���6W;5�48�����S�U�ö�z��(���1�ʵ2���~��r@�ɑ-�t9Z��	G��Wq�P�UUb���Z�Y7-�mw݃��m&�e+����ǣ*�t����ޅ�go�
 )�Ȗ���7��vǧS)�F4_28�����-8y>�4�,�7�򰕻���N�>�폇
�	in�l�k"���s�n�;{?UT��]m����	�p�e��ĳ/��{+ڈ8t&CY���H���]ǎ_։����Ij��!�GT��Y����O���,�j�G���ݲ�s���k4�x���=
T���JV���k�ǿޭ��FU�4�$���PO'�=�4�mk'�m ���w��s�_�揿�Ny����g[�]si�5֊�Y���DH��	*Ā��$��<�Z�a9$�\\�͑ui�q�qs��g߫��d�RE/�� m{L��fN���lԆ�j��`N�����8��Yx���ĺVib���b8r	�5�ȋ�R8�,��v��g��yg���o�����{SdQ�b����v��l\�x�Cqb5r�8����cl�.���k��4q�K�3	�x���\x�n�z&��"��
Jb�;٨��}@�
9Ah r\;�C�8���g����'b+)�b�{G������W7��~�<����Vb�=�(X�����u�IB����V>�O���^���Y&���B&B�|��"w�DzcR�X�iG`:2$kt2~j�D��
#AX���C!5�K�
9e��I;�A;�1��Z��A���OU�N]2�����p�왘�^��l�&���d�Vy�nܼ�J�q��Gu1^&�ٽ��w$���AM]�x�>}��t�c��Xx�IxM�BV3�Ų&�U��)�u����j�����~yNء��fC��*���cO(�9	��r��%k�����Y��`���0q�����n֬#�ݳ�_q)���{௬�2��Ejߊ���z]s�Er��J��ssS�#&�N+�L�(��~��C��H����m�q����p��~4�|5�l���Sε��0������ވ��Z�R]u^�͟���jmpWU�u �*�5�V1.�6C��X���"�2��8�B
�A\�h��������a������a)���AX�hE�;��93y���s8�J�pԡx�ŗ1B�w�vP�T	"8l�:K�X�lk���a�IU5U���є6���Ͽ����Ւc)+�+�����ہ�Sg�����w�!�ƕ��:W��O���x�b�m$�����p�� ����J�2DUe�	��;�=��N8
�=���ե��n����h_�٬e�T���~������[�];q�Y��ѧ�jc��U�	��Hs��*�S��U�x��O�ǰ����s�8o#!��S�
���y\Z$F[]%��;}]�J�S�<��� �Ï׎qm��n��������SY��t��v��7/Ɛ����/��6�\��N~�k�ǉ��<�GŸ�{�)��ޒ8�b�N-�՝}�a��`x�ǨI3�igV��H~�����U���������f�x0�G�{��='��T��2u��x��e����g�QsҰb��y�\�_|]ַR���U��������-g����j����	���BF��������}	�S��aY�����%ԉ�fb��W���/ 2�܃����c��1]x�IX"��S�#��k����W��k��⥷?���O�C-����b���~	����j���'UC��:�$����Po'*}�H��x����Se�����k�؞���`�߯F&E�A1��(���e��vP��_m�Ï�^��E�CVB%7.8�X�׆�|��_�?��_p	j���,��w���}��h=�]}�o�$F�${���8O�3�a�����}��Q�����&�{�E�"�ʢa�nXt�blڶU��� ���e�����h����/��� ��c�����s�T��SO�8�m$
f�1��M��Yb�9a��T��ֻ��q\��&�ׯ���=qL�l� ~ټM�X�0���2tuv`���p���[[+����ܻ�,8V��$��Ib\��A*�D��[�p6oZ���x<5���J:"�ӫc�5r��u�m����8h�>���d�
b��
�ˈ!k+��_����^�두ɁX�u\��D�~��	�|�qX��J���n�@�"VW�&MƂo���Q�~���7O��#��}��ޯ2�vvj_�mN��!���?w���ߡӺٜ��O�0����t���:�����wk�����\|�;�a�����ƻPrP��S>��b�#�p���p�fXI̚9���,.R�QɾZC)��j[�`ѵ��;�DM�O.C���!�}�\y�)rAR8Z~��G��Qr#��L����9�t�{��Ե�%�+?C�����q�
≠�}f썟�3IJ�2y���������_z��F��?���ᖛ�DahA%���CO��3�T�_`��:��m��p����MB�Sи,�]���S�������G���C��J$$�>�سUկQ�a����+@Vt�Sx���q�9'˹n�w�a����kM���b࣡a�\���?�
�x�Œ�_��:q� ���$M?p�}����	2����>�C5m�?�����9�gk����%Oaٓ",�+�����\-���*z�̞�d2��ѣp���2�aFA�T.�wV}�L<��)�'��O8�o��)������BA�QT����N[�}W�M*��e��^�?��v����a]���رc���W%ٶt��o���/Ma�0V��MbuXf�{�I�"QL"#0�e�d\y�M��Pd�S��h
7�v�z�.U�s�d|��/rH}�q?e<�zz�¹q�S��]G��4J�%ӭ���+�b�~�h�K����"�a����\:"q�Ă�j,��H��kl*�L��޾<��k�o���6ԣH��v��d�B�DW�GrX���b �H����W�>�2�>�LjvaP�bD��.����o�n�\�^X
k��|��M~�`�oJh6�9�^}�'bp썲��D�iFC�J�z
��F�������\OVp���6��W�l�^���Xe���.L��'y��դ��[?��OH��S�5�2$rhG����`�>S�dT�6���V�d}rQ]:���۟����&(���1��Paշ_��3`I%����%ŵ ��xF�"w]=�r��	��!.BЌ�$�Ï7�P�0A����0�<����,�;�IU70���xb��+�=R��Y1�}�9<���q�\��)����T���{�H���|��M0{M�\T�aCY_��x���p���ᦼ�v�R����8Z�Nk�r/ɥ-)XȨ�7�P������󶛕�'��i^�D��0��wⵣ^����@US��xo��������{7c
LጠR����8b������v&k���[��^J�H��Q�X�A���?���>Y�~i[R��&9��x�]�!�I�MYT[c�)�+�E��>�g�q�+?::�T�BCU��4�E	a%��	�O�iO˿v�iS)y��p���^��� �4L���o���q�Z{�h:g�N��{L,�-`Q��^~E3�W�㲐2��U��̴j)REk�e�f�I��l7-;�(B�2p�e+yh��n/�� /�BV ��8�[�RX�n�6�V%��%x��!��Z��kל�H-ٱA��`OI~��rhr(k4�0.Vr�Py�g��
�K�,�q�-��oٲY:��Y�\(�Z��:�&����]K�I=(��;A���ς�\��F��lh��ZsHm��dY�cܘ1����͘@ki�pK��+�~/��,V��������VSmVUv�ɥwhY�#�h�K�U��Sو��z6_��_�cϝ�#��O?b��:�Bq{�f�Q,+�5imn��U����]��(��O�X�$޴ifN��9 �S9E˄*+|2���;�d��Q��ۛ�{�2�)1�Nٟ\"���r+	L�U�Ex��g5��Dfn6�1�ϒx__�1�!��Nb��A�/7���p��5����Y�8,v
�qP�e�<B��#Nq֢!��RmB�PJ����5���͋j�	ڢ6����$����j�����V�*n��%�8M_��6r���/��ʝW>���S+�^A!��0��j
�0d+�Gz�eC*�딄�.h�+���x9tӤ3H�Ysbph�hN���
j��%�|(�����8�o*��S&�)~f�3�����|^m���f�6l���ѹ칛X��֫�����Il�ڴl�jl�x��OPFcօ�Ⲹ�H\	�y���5鐏\h%�M�竀�iEMm"��,��\A���FQ7��)R�%�jj�Q���������gsV��^��������CSLdҪj�[>�W���<VA�E��lha+�EB��Mr�,�$����&#2I�t�BM�'Ȗ�%�$����4�Y$�3�(76i7��L�\��Į$�-i�N����U����@K��-�|�ֻ]^l��&F�E�۽]�E%��$�n����tj�G�%Wݍ�x(�͞�D����EM����9A"��Ea�)"�rL�Q���Z��d�?�YАx��(�d�$�C��Ї)�Z��b��_�i�L��Y�
<o�	H��UgS4
�P#Ȥ�fQ�Z
���A����f%�a�z��v��n�P�r΋�˥t��ZJ��G����0Jb U�ۤQ::?��	U?b�r?��cBª��J����Ⱥ?
�q�9�yLHx�t4N9� ��Z���,� �#3�#���j��4j�����g�1(�˻�!A�1H�;2���$�i��UR$&qy��s`����"����Il��V��m�����ٍ�l2�T�=���a3��پ�C�8�xt@�/�h8?�is��p,�c��,���A}V����-hj-W��r8�S̮��yy��@��y\���E2_RY��  �*p��{w�28c3mn���u{�k$�mi�F!�F�p��E��l.Bmu����5cE�Ţ�m45��O6��ʄl�pL���`0l��tt�O�5j9���r,r9���
5�U��ģnGY�Wj��7�D�LD3�L���֠@�=���-��@@y�dVy(LrX�J�B�p�p�#���C�P.���d�����&b�w���g���y�ʴ4�iHH�]�q��Jf�nBDb撬?˽���y�W�`���1����'���n�hP0g�C˙��KT<��ǡ;����݋�����UĄ�v�^�;ת�Yƅ�z��9�WL�m<v�f� 7͞cg/D&�W�ľ��?,{���#��ǏE��s�d�8���8R�5r�95�ѕr����&�!ә+K�C#;�}�g��B�BRp���
�F����1Y�ֶ6tF��l�%���QQ�*H�k���B^)�oP���}���O~|_P;4����y�~�m0���is{!���	���@7B#��l�2���Ѹ��7�p���r�ܪm�&/�T��;p�⿢k�1���a�	zsR$KB��'���O���w
:�j7�N��MMu�y�Ƌ�}�}"�RV97��L�{1�1m�IY1Ғn��-ο��g�R�c�g�������I8UK�2u/��C�ry� ��&��ȖXv��Ήѭ�r�b���(�E� ��%��bb��|���R1��_�7m����G��Y�≗^E}�B�r����;���R��f��^�]��iQv!���9uw��f5|��Z��	t�xR¤�>P��	9�#�Ngr���+o�%_? };��ϔi�a[A�Kl[%�Z���>���r��0)��l����9�����9��ߐ�͂85[\d��c��m���87k��h��U��$�q��#��bnft��Ѽ�&(�)��9s�l���i���]�dҤt(�����}8����������xd��5�4<b z���Ő�ޅa���9�L'3����Y�0:+-�HHV��<$:�����J9	,*�d�s�q׃�k[~��6�]<�d��1�����_d�oO�/PS�šǷ�m�6{�l����:Q��l�,���OJ~?�I��;�l ���aT57cd$���Ξ~��e�"NȒ$�V�X�8�X4����Dǒga�����"���O}��ׯ��w܊=�,���#9e�j	�‽�	j��,��Ϊw�o���b�׮ߢ���_���s����E@��+���|"<�g����Nyw��	8\^E:D��CC>T�Au�\�e1�v���l�<���ߜ�$���ǆIYs���y1�^-����c�i�л}+n��R\w�-�����=���1���$4jP�^��5��"g�Fө����%�?�p�w����SO����>��fSq�:�`L?A?���oK��r��q i�~�ˁMk_{A ���~/�Fk����e�v�3u�r��d�>�Ȳ�l�.Rf^�:��unCP⫷��5��N��Y�D[�z�;���ƙ��Eb�M��K8��̩s�Ձ5"rA�].�Ȓ�K`��Ͼ�lS#��8��#���b(�FC�s9BuC�L5bY_@mc�"
���K�	�X><����ǟIL�R���f���V���C$Kʓ�QB���x[�0��~,:�$��]��:NL��K���_�`��h�}E ,y��{����s�<��y6lآa3�{O���P���}��zl�F'94Jh����ct]=�A��W'n��
|%{�5nՊARdh�H�Ë�X��V��l%��d������#+��K/�7?��j6'Ux��U{����[��}.�,�6*\%���K���E�c���pΉGb��y�\6EU������g��ܬ��!_�XmP�I(��?b̨*��j�&��u��?�\U��45w*{Z��B,��S�-G�}���
�i;�z.9o!:;1k�I�g�)ؼu���
����&�:�����m�N6L�Ǝ*�n���˸���e�޶	�z��bIDcQ��9��e�9�c|��jt���akI{���;q�������7]q֬�Y1�	�#*��"��⾇�E��ފj��/���[n��P������_�S�t:A��HR5��6��~�;���ꐓtś�*7��э��u�_�r�Zd�|�^E#!8�����Ix�<�MK�v�[iq�w�� �}]]8�ع�7W;��T��\36Z��Ѐ���a��-:��>f4,�m�|-�q��GP����^BN��І�}���s�x�jlc��֠��Q�t���(]d�:5R�?�\[��'���0�E6t;�%'����GNb*��k��I���;�	�K�PĮ=f���>����;�nı�A1l�z	kH.렄=�;{���o!X[�q���0�"�����QMC}M5��!9d�nFJb�@�W;-0؊�F<K�291Wu��S�KϽ�"�8d6�	i<f4��F�Pps�ކ_~W�S�ðrЮ�!5	**��U��FW�f�5�	�|ℳ�Ň�P�Ђe�Wb ��u�k�2��N�
<~G`��Y�P%�jg�.�=XT��1��~�\Y�܀��P	zb��Xp�1��EP���d&���%���tK�� ��B��v0��IP������ ~���pb�=u�J����$-XS�WV~�ۻU���b$Cbr�(�����3D����Mn��IR�z�x�ض�?�W�Z�ږQ:���=��T��y�)\tکH�"�\��M��#��0�m,uu�����a㛜s�\����S��?���:1\�+���5�A1���?��K��ޫ-����n�0'\���׫רO09�61�.g�r�i8Kb$��r�_������������^խ�͕竞Lvd@	��¤��K�z���{�a�&w�՝�C����Ko��Mn�gNAZ�K<"��n� ��)9�x���.!�����V.SVO{���?㶛o���?�R%�Й��"�����uH<�G�����q�z�#z8��V,��Ϩ�o�hu���Mò�Z�.�U�c�9'�c�Z$��p�%�Lđ����ʫ+7�}p�Z2�&� �Ay��0�h"�U�����n5q��$f�����2�U�R<�9���\ޅ���1�x��٬3.o)��f��6��?��}TVU�AJ��ąt�r�W}�3���rlټ�7�u�0="P>P���}���JV%na�:�i�%s�N��k|�r`�G��#/^��~�-���}�+�wHJ�g&�lrQ]��jҾ���}W]r>��L�s
c&5��~���-�d�ysQ��<�U�C�R���<�'M��>�
_�V����d��FP�W�>v�-kc�ꖈas���U�ќ�r������P%H�B���J��c :�iN�&*K�/��c��t��|���`�8`�&$<��ų����n_@{x��T�#\��{�p�<g���Y�� �g��Z��t	�����z��*�RńnFP_ڞ�#����e/S�'��
�qHB�\�%�?�� C��I����|�Mbت���0���r�ƣ�lGH¿8��ZF��ǟ@g��'��ԉ1`����|/r	��e�nډ�/>n�K��,^��=;�"Xz�8��4�g�}dx��w��T��ko���/��&kVɣzz�в�t\�hj��1����5Y[�p�߮9�b��}8̱��^0�0�������`�G�ޢ��	�X����iLU���hv�o�c܅���cg
��V��k��G�+�b�l&�ڰ��㺭���r��Q����+&.wMr��/�y��s�컷<�l'���¿����Rzx��T�1n��!�u��>C���f�~Ӄ2>&7���*AlaeDe68d��������{�����W��;�tTxk��2b�����q1Ӊ���Y�&j?�wK%5Y�*C<��m�y�͌�U]�pP��P����Y��KZ���9�Q�4��
x�)�2�E��Z�/K-0�O���cO���7�i�$�H�iծ%�t0��wؘ����x��ux��K�Z�DBQ9G�^߯k�7ƿ3,E���e�\n~��{�
B[�d����T�ۢ���%5G��OO�X�!�NA��f͵�����ie���;c-�ڑ���r�|��f5,&�� {��R��Jy���1ޅS�4�9Y����:��R��f�!IG�g��0��>���b�(�8�A���Gxm�{�$9&�m �H�Y,�e]c#���N0ł�mw�[K��CIb���Tr]�X	OT��<�X2�CI�J����ڊ�/6Ά��^�+��rT��r��9˜�x��/Q����Ǟ}Vs�^q^d�S�@���Y�Ш�S*���f�8f+���ù_��e��R��f1��ʰ�h�~�f|��:]d^LjJ|���e�њ�d�����a�:���J��,�c�2�V
4�D�ףlW�X�W0���L�qd�����H��]�V�����1���u�.DM`l:g`4k�3Ğ������`:�:�YݕA$�:M�w���h�r%�)=D6trd�9�.o�2���H|>�toJ�G~�GC����P<�,a������(�I�#=k�|��e�����px�G"!��kw���N���P+~�8�KWTNƳ,AӀ)��2VY��X4��v�w��ƛة�F$�(B.[PV/�KkM,^#��GR�JsXɐT�~�X\6���D�3�5ȕ��)/��;�숁"��u�J�}(���;��T���F�'��4�_4�R�W3f����:=��O�|�˚Smv��k�r��њ�[���*��QxJS�H�P4�J�.Ƈ0�dH��3Y�TV"j�J�����!�˞p:7��Em`�}3�-�Y95��x��p���la�?�%���4����`U���Ǝ�;��@Em�Q�ZdM�sQ2�v���:���UQՠS��)򑦀{�q��)q�9�o��t�$��Y�@�ДL��y�w��v�$�x�"*�R�mЃ�|%�#�P��4�U���`_�c�,���Ӟ�)Je~s�8ƤV<%�2d-���Khb��Ԭ�i26L�YaLy��GЅ��ס�#V���Sq �FRY�d��$�f2)Ë��g!5�III�1�Za��cX�Ƅ�Cg�%K�Rg._�2�g��t�5=w:�P� mR��������Z�|����k��hz

z`�2�ڽ�?a2�ʇ��+�{�,�RKE�7��u+�U����
�>�rr��qx�lp�h|ϰ��'���D�f��*ɩ�G��,cb�0�W(�3)����'g34R�]�o�I�u'���5s$�\�ϋ��9EM��3[�=/��A�h�qk�h��u����>�fEwyU�3�~�|�LZ"7�0��l���#{���2O��\�𛌰DɕL�+��V<��/bX��$�v5P���<hf8S�I�|9��~6g��e�]��,�u�����2�`_�[(�YȪν��d;�V�ؚ�:}~6/�W,��T���#���w�������2ИP�F~	a��H�\�K�:5�Ŏ>#�f*���f���34�'���ţ����aq�/��Џ�MQJ*�E�_V�����t(
�������C��n~���C�?.�<�9�iUU�24��T��(?�d����Q�6)'o���CCz�8���"$J��ԩ������L����S�<�?�J�����I�#{R_�,�۬���r"W��|@RB��?����_���׵���Waxp���e��`�2��I�bW�46h�E��q�&�< ���E+��d�%[3�oe/�~��@mu���42��ؖN�F��Z��L@���(��l�b�@Jb�l2��Lս-�;�dݚ��m�k�L�dT�k���T��l8���	�I�k8B�u�Ms_N���n���$��e�ض&��"e�i4�6%q<,���re�g)���3���@7v?}����Q�쭐���=jb�<���Ԑ�{�V�4���XDּIU��N��r>�6���DG����yN��HB�P���'�{��#!��Ў!9>�هym��++=���Ѱ:���tB<� 48�G���}�ǥN*/�q�7�%�ce?Řq�c�Q'<�FF�%W#��X�v�%���e��8��p��>]{����Le;p��.����C�P�d�AU�?Y~ҽE�C8bΡj9���'�����_)���sr�y�Ԙ���h-������gy��ӎ��~9)�#�Y���\ AR���>C���Y!Ƙ�Z��{.*�^�䔒��00��˯�!P-���U(ܔFpl669�q�� C2�S9@(�DB�}JMp%ۂW-fCq�?���1q*:N! �ن-;���'�����P9��T<��brDu;��G���"=�Z2��s/�*�J��#��[DQ��c�m�I'�֦�FBhijB����;�=���BK�d��f
9
*�T����W^���h|uu���7H��Y�~�-\>�z��ߔ�;3���p��)F�F�>��e�h$�������g�dJJ[X4�+�uqk%�_���������b�Y-�g�W��|�n�٬Ȋ]��|&1���A���j�UI?�1��Yd����;%�i u�xw�ю_����\q�"�-y������r��x/<��u�=p���*�~�3������Ϝ�y�/B44 ����;��P�{o����3^z�U�ׄ��~T�u
r~8��n�A��s��o��/kY���ߍ�n�UB�DÂ"HYX�{�(�J��ʇ��;Jb�8B`�Vң{��;Z�,��=We��#{F,��h����|���xވ���&�f���_v)R��R��PW�Ñnܨ|��Fe%�{mZQ��p�dpx���pႳB	�kK�ٜA}K5F�47����t1��M��&�K1�Ħ�ӎ?F�$3�x�D0uB�,�&�5�`��yX��U������+����I��S��^SǢ6HZ7�zŢ~/{��|N�u�|<�ߗP3j�[�s,�0�1�����<�tT9$S�A9T	�:e��y����>�!$���l��e�e�F��� !D�3"Ʊ��VTA����w�����O= �3C���a�ƩwB9N��Ʉ�xעx����>
���RK�%s9���Ur\�yTW8q�I�h�)������0�٨��_s���K��e�Ci��ݠ����[���?\����ڽ+V;�rV�aLӦ��o��/Ph]*g	��(t�,1z��:�`"g&��S#�<b:&p�y���ҾR�L��0<v򯜀�P���!�(1}N�#'��������=}�:]��D��TLP�	q�,<K{B"�l� Ҙ �w�� n��b\w�mh3�pe�/���`����F�غN��M�]PRPG��|7,�7��.1B^=��EF�6��N�u�_�1��Ⱦ_�ܤ�LO1�����q���D}c�"D�Е�$�
xp�e��?����u^:���a�)�����6q��~l��L~�Zq8�-�iq�Ew*[H,N��{�4�E�kh$��j�>�ZO�Ňe���V�{�Q�w�4��U��եsԕ�%��a�K��0 ���l����	!�E�/�#��b�t]��.��)�:{q���.���*)��q�����NKR�-d��CO���$ھ�Yy�Ҳ�'̙��?r�{R4�5iv�u�D�a��i��U_���;����<B�Ɔ0��g�?;JF9وQr�bho��6��GM��^r6�Y��[����:umc!\~ѹj�yZ�M��ݲ
öz����O��g���ӝ�L^�e4���.<��[Pc%���V�X$Tb"�c�f��>1�u%���sX+6�Z���A̙��j|���D��Q׶^	�B�o�RE�b<��Ǌ�N;�~�14����RN8�7�8|ξ�?n�}�v�v�����c�D��s��v"%h�3O²o`$S�l��hE¢#7�漳��P;��PV����O  �/IDAT/r��M�{M��)��k﯂�ת��S�f#8��C�{��+�
dcv�ݽʤVm5��@�h�ix���PY׊X� �%A��łE(5$�����z�C�+^���R]�ƻ|�-]��]:�ː49<�K.�s�G*�ƴ���{T����q��Q��H�1y��j�1��.w�+�=�P��p�B���S	��}4��v��k�h���嗞��j����k.��w�.WSR����vG͞���*��[9a:�~g�|�1�io���=�hU¢�\{��x���»�̳9�\��S�d�'ae�O�˗���u�0y�D̙�?F�	2�c��ǝ� ��"@NB�
97\z�怪���Kν�׬`@��J\r�4k,��B��}6m܄�^{��'L�5W.BSkZ��W]~	�|~9<��ӋE����"�Rb�8�`����|�O��m-c0g�~b�"��ǉ�~v�@�ZU��'�#^s���$^���m"�{���t�NN��;_}!�{whG�9g��寽ב@8���_!�7E�|�J~��6���!�P���j�I�x��y��=�)��7��	�N<�h���pWx�5�-�N/z2e���L��3�F���O?��S���ާ�H��8��eႳ�+E�k�	ܻ���Շr�hΜY8��c��(Q̱��3/���}�ũX�{6�l\���Sf�[�r'~Y���Q_�o��9Ys�7�h�\��2W1�żش���Y3�3�ؽ�Q'^�j��6�e%��Kl}չ��F"ƥ.��xOָ� 8L&�� ������e���_~�V6����.F<$є�駟���|A�	q�TG쿇@�0E� B+N>�r8e=��9�����2�sJu�Q��9��3ڕ�K_a�a�Q�M�v7ብ/��k�&�) v퍓�!�>�(얛n�mw���ZED���|����p�R�p��g���Z�������8\r�q`1������l�ju��I�'Y��c�;ब����^vf�.K;�"�E@łQѨ�Kl�%EM�Xb��޻��R�)u�e{ߝ��>��s����1/�3��/��{��|1�=�TTF4�y�&�������bkO�.�q�<,�j�:��5���'+X�����J�\TWU�Txw� ���[q�i'a�F�e�����B�g
�|�C��dX>a2f�|6��y�aڰ}9>_�3fN���=K��{�w�C�!��?�r�=;�5T�a��T�" �e��Ւ=�W��O�S�i�|�Y\���X�����مj0g֩���aV�(�)��O=�Pȅ��r�?��s|�����a�|��[��������E�_�8���L�ʵu�*1Ǚ�OEJ�_<w��7��o����tk��+�J�8S���z�٧�{AEM��p#%"�mL���o�ޏ��4Ur\^4u���o�}��	;wl���������(��x�ko�M[6+����[�/V���0[�P
���~�x�%��������=���Gq�)I�<�eRr�-������*�4�̊�qa{s'^|c��d!ƍ�����^���}��"I���G���Pm�Rѳ:�r�%߹���J�-i��+ƏESW�x`�V��^��(�u�J6����j-B�˅���p��WC�)�:Z1���x䩧�K���[���P�KgW^�7��k��UM�[^�]��x����PUU��;�B��II_��k/9�����]���uH��H��W�-�]��\���X���{$F�P9I��&����	��	s����3vIǺ��@��רj|Q"�I�X���l�Vȳ\(,.F�^V��^x�ކ���Mšr�n�/��q�jz��@^qwM�t��z�U ��B������Uzf�9w�Sb�^łSf�����6�~�Z5M�b]�(Gʿ;0B���G��zI�5�f���b` �<�n�寚�VVVHZG$�5I�K1p1����:�qH����!����;��#��C�>(9ߑu���m,p���w�W0,�K"V��\?�/V��SR�$\��bN�u>\�vx�ּ阶��5#q��+P3�AT0U�aܤ	���;�����-b��PZ4�}��eǴ��X-�5�;npY����rF徾�ҋ���a_�iސ�H/fU!�!|��L��j�0���]H<�ۚV&oΕtIx��ˁ.��;�A���[bl������~u�\(��n+:%,�k������Hj��f�G>뛯�/Ѩ-H�X�8s3�吒_����:�������7�t�K~��8}�	ri��{�=��/�zM!j��3W���w_���`U�v�S�
l��e�B�1<�m��<G��7����T����;;*9��n6���&$m�@��v,Ռpw��\�D��硂:,L��_��tF��Ƭ�h])N�*��!L��V���مڱ���ډ��g��>�d�'E]4:C'()���zV�\�����5%H�gC��@����=*����*�O_w�Dz��.�1�i��AY�d&�;x��zesc4��I?#Z��|�tRĠ֥�_�A���4�����?|�">ڪ/�MD%)����8��j4(ˠ�
t9�;r�7'iߒO?C ��Wf3�ۉdފ��4�}����۶n2`Ţ�>����];�0v�8�r���Vt)n'+g8!�c�V�<�Һ~YN�{"�Ig����<Vʾ�$j	(��6�;��[w�cLM}}�ک(�Pf얱V��X��ёx��+h�| ��8�z���{������F��Ko'ےD<�T��ޭE�|�LZ;�n(�-�V�<cKk�$<v��7�$E���|���L���M�+�}�o�q�=�6�����結�9��m�-[�qܡӱ}���n��U��(Ȣgdɰ��v	ه�Y��S|'Ki���xUD��{��nm�ڵ��*�+�l�!��R)��M -[On�髳�G��@8$��x� \��x�;,_��2�������{�y{d3�r�]rpb�uP�u=Jx��uz�ً-$8/��*^�j�����Oqp��W-�d�L�֊��)'����G�5k7��I�u1�ɔ����v�<�Y�݁*Zh������E��
	��zXK�Y[Ѯ�����pVD賻�ˠ�݇F}eAəaF�َ�gt��-�Je���{w��Y��Ԋ�&��\�!�ȋgu�j�<B�w�V0��_H<�+��)B�,"��]��μ�VտѨip�pDҰ���)A@ ��;�wb��)zV"�h	�gר��K>�d���s�9���S4ZaD�*#�<����5�E��w!+gBְ����]�k�=%*2ǎ;@�#��#
�93�ZP�<{䡠@6=/S��r��>�%�����~ZēCJ@�P�v���As�3��$+�[��aZ�����$�M�E�K���	1b���zVG�X͔����C��A���s�O�h'��eɤU���0�ɽS�/��ģ���Ds���,��Lgn�[~����SĶ����bP,���K����JA,����R^(���K�����^�)��7s�ɞ�q5���<H���u�K)����K; y	��e>�rry�-�r�57,A<�SB��;���\�R}X6�'����\�I.��=9)x�k�@Q�)g@<���E��J�9���A��`D�!-��W�%�L8�S���%���6��|���6��M�/I���S[V��T��$~�R�,�P��*s������1c��/m�!����q����95;�ۣ�e��<\<0��'�%h��	޾X֔HcQ�]�*	��������۪�ƴ
%��C�#^�G}er�I�4���H��o_"�t�bŵ��NVA,���1dz�0���X�q����!*���������HT?��j�p��VY_�і��_B�r�H�e2j�fU%� =vV��,����)n�`yĹ<u|�|j+�;R���e�^�l*��	V��9�)g�_�,)k;1i���x�I�B��3^E����#N��%����$��{J�wb��UC��;T�!�. *����o�Q���+DmuD�gPE�<俐�Ш��9�mڶ{���o��X��Y�~��En���/8Nk���:iEqKD:,��X~��G�7���>�O��N�sDb�m(��G>_]�FU��x��Wq�a3q���l�?�7��1��p����㨣G�압AΉ7��B`ЕØ���	�Dʰq�]�Y�䢐��"��V��Ov5w�WY��B�C�Ca��S׃���ˍ(++��"v�1T� aj'B��Z���r�&�9���*o�,����y
q�2�F�U�솝=��b�=����q�r�zT����Gi�(M�C�-y_2CyC(���%�S`K�)i��M{ED���zQ�.rY��=�U���a���?n��Ʃ�g�����{���D4_�<�a�u �}��\̌���9�3$-��_���|&N��t�[+����g����7���=�vb�ѵh��@o\�s]!�e���ա��O�Cr/�iz ����S��b�ן{�)x�o��,#n���j�}�y�TM�9/6Z�y$B˸�h�a�H�7��C�͊�%4��k3d;eb@2�>I1g(v�B��=�%s�C�?�?oބ����)�������3SW��[�[VY� ���i�f�`"�8s	9���")�]�ȴD���;�b�)'+�%�R�S�D��R�?�R�J֡m�j,8�x|��F��a�(A��X�;�7�R�����A�t�pgH�[��[����#n���9e(B�t�&�3�Ð�S�ڡ���g�t�^jH3��#�n���;4�U$2�'�35roi���	|bT���˙,���c�Hu��c��"H�32���ℇ�ǋJ�Z��C�`L�։�u8��ִU�W�s�/��Eg�釟�M�_"�t��z���=��gw⒣`Li�Ԓw��,*y�J�Bhj���u�I��+p�,B_�.�}�	x{�'7�-�O��C+]8��rQ��|�E&E��Q�?���i`��a���T��%�����ry��dyؘ���I�œd�v|�ŏ�o�q�H����r�I�0L�Ar:�刈gQ-!,^����R9H�\�2������.Qa�C����o*�]B��s�$i΀�_K��(KA�bPz�bX/���2�1���n�Ö]b��+���%�����	`�Ֆ������F��ڱ�~�	�~%����#���a�����/9��J%�	ԍ�C�}�P����T}�EX0��}G0c�;>��+8�L���c��8�!�)Ǔ�?�"�
_��Ϩbݦ�?�#�C8�����b %�v�q���bP���W痭���sʰFR%�\�e_��3构��/�m�]�G}P�=�2	w�^'?�hŦXlTxs��o֙%�6�4�lAOB�@N?q&>��3���éMQ��a�=&`(�Duu��i�n!�<��xa�}�{M�i����p6�h�g_}��5����w��b�$�Z��=W�p5��3O>�"n��O��	p����?�@_/���at��BEbr����߂���$�iW�iS&�}��s{���۴i��B��}�H�S��P����C|�O�X��Ľ����N9]M�p����e���e�89;�{4jBF:3Ut��w���UU�2��Wປ���n���͘!f�8̥}(Ko��Ѵu��1����O��6l4饝�d9��ò��0y�	dp���po'�j+��Ѯ�NIy�p�"���[D�$a��5��9'/��_�X�?ѐ��y[�[���]��"^�p8~\�F��]��LQ��,���n-����ےV�<�'�������ϖ�3��Ǎ¾ǠU��`"�)J/�p�>�"��~Ŋ6�7?�A]}=������W�(�� j++1����I�d�~�y��y�%����Vᮇŵ�;O��8N����E�������gH�>��l�JZ��+�UG�W�x��:U�N�OvH����YQ!�y��fPOBȧ_|Q1^fpȄ���a9p�a�	�"��e�P�'Ie��$J��G ��?
�xY�&2t&������g�2[R�~-��|���#���P~�svI{�~	�riAYf��'�˾1:���z�YGLQ�|����2,t汣����J.Y�Q{�ˢ`R"��^x/<19ȗ�� �5C���j���%k�ToA��F�+bA��9���G��5W]���-b�+1�Õ��V*�UG+��K��#���HD�Q���&y�K�ұ���
TF%E�1�õP�h��Dj�n�ф�����Z����'�
eQ����񷛮Ց}v7��;���uI�ŤF	��;�eUuz�fRL'K�u����ҋe���t��L���55�����q�b���M�M1=kx2h���c/���/�X;�ӧ�¾U�P�9)+������E.������W�#��x���}��:U<��:B���-�ʭ��7n�ۋ>�W���`�5���k��#�R#~��4�Ս�u��XOG�:
��/�^ۻ$�e�|��i�BҔ���77a��f��������㯼��.\�Aɥ$:Ł����5�? ��>���K�B��o�>��Ͻ���_����_�в��H�E
vu^x�	y#�N�=��S�/^~�-s�ab4F���{	M�0Pf&c$��|���#At�,���-��T��r<��38���J�P({}4��g��iO�m���-�F~��ZJ�Pc+��?�yg���E�DΦ�%���g&?~������$�N�!%��%�o��a�䒛6�Cy�\�T�� F��#x����Z���;��wAst�l<���8��Y(��0 )A��Fl��ɲ֟}�v�����\�{(�Կ��'!$� Aq̏=n:cY�e/775�9X/�;j�,E���/���Ԇ/��&��Q�-߃��^M��&U�����#�
�=���Δ� �����񷫯@V�֍[u������;���ri�|�AK�� �,�S�j��'��.�[�r�o�F���a����n��/�F���"m
Vœ$�G%��wދ[�z�
}Q��)iQsK�B⩹sǝwK4\�C��Kl����_QS���{���������J�Q-�˯B����MF͐!ӕXފ�xϚ�u�V1�5Օ�'xʪT�kSS���K�j�L�m�*�;.��p�Қ	q8�,X��H���ǟ�O��O��.��k}�)+����U�F�f���N$QQ^-�<"g-��Ũ��e�$f!�Uz^J����շ�W�`���%�kQU�=r�|�Y\r�ɱCb���378�F�5���a9���H��p(�8Aari_|k�?�P$%$rI��i�~y@��l+S��y����$�@�/��O��3��kT{+���߮\�"Ov�G)�x!��Egw���~��E�g�=��q9L�J�ۦu�$�hQ�S���K�v4�vj��$�F�����9��yKI�8������k���L
۪f`��������B��^b!
���P�B�j���%�e[��l���Z)LM�`E-^~�C̗4��0iǨ8�˲-�=����=^o)��rP��%9�L�U�>���5�d�ظy������e#{6����}a�y8���� �O:Q#��ۛ1���ښ���+�ҌP��
IwyAh0����<E�7��CO?�1��Q.S�Uъ��������EwM_���1�fy������e�im9ƌ��ؐFl�]ʬ?6�*Yo~)�2� �qM�;�(K�����0A�~����*����k��D`c�ʤ�܌�ha1S0��EcC�oذ^�y�r6���͖>u��V�����S��2mu�I�H#^C�u�1�^�y�$#�����*{ʚ�=?���rȕ���7Cbl#�SS��K��y�-�T�m/������y�J?�Q
�y�����{�9T�5�e�J��H�?1,a�ʫj̈́@a7�NQ�2������{p�����UzD�d@6����Ҡ��V�l3�㥕����~mѧ�(��Q��A `�}l�CBj{��Y�S>����
��h1R9�ؕ�i;�
[9�(��'��0���}}zY�����L[��V��J�E��Ĉ*��ݨ��̌�n$U�N��s���o�'�`K�A
�r T�`���' c7NixO9/$��їCv[��G�Z7�Z8�Fc�LfT�D�b1j���iY�@�H���W�pWUЋj4�_���\�(yH��)~�D�Z�ꗦa-w!�� �h:u�˕�����|w��IpɅ����>�L�M7�_�Q��CY�X!>&>�0�8]��<'�Un����G�_�9/RA��Sy:�Ŭ��e�v�R
�$�<g�D5-�׈7���O��g��F^B�u��d����T� �:'����v�*���V:NO���$iG�pJ�u%���E@"莁�����p�s��I�M]3�[H�hX��|�������g�AG�G��i����$�����a��@N9k�e�ցgF�J�47�xMS�jf�
y3OoQ��´�	V��%)�#�mF	�LD�Cl�ʁj�ҙ~9��B��ݦ�X�MQ^��G��Z�����6^���C��e��Ć��g7c�~����b�X����"o�K��E[6d)����h�Rs�R=��TNB��pP��d��[R���u�a�(���\6�Zr�~���0f���0�R��_Ga80hLiP�b���2���$l.�6nzAM��*���jD�sT��K�f%��-i�F�]/�u7�C�xp����N��eux+M�!\�F�6FT��-���K¢�UVCX�ZuS�L�:/bS����Ou�Џ�0x��r�)�{#�m-�?ԛ!���AE�ZJ�Nco"�v�,%b'~�/zΒUѠ��%��nҤݓ�(Q�J$6��u�X~wXR���YN�r��� Ϫ�,z�ͥ�K�E���
��t��
=(X���s.�7Fg����F?�5�����4�Ԕ��6��q)�h�n�E�H�`U�eA#:��.�΢�Z��+�ն,Ŷ2�m	 �25��UeUC��E�)吶|�����w�����C~����D2�uʛp	F5i���Ezu��i/�f7R��+E�a��+�M�he�v�*���D�9ӌ_��Ō��6f��xMs ��u`ii�X%g�	�J׍�2Ki�yY(U-�8��� ̳�,�'�ǰF���D'o<,�,S���J~*�[�@����	(	��1��U�'��I��C�:��h�׈oa!�\2�h���a���Lu;l��I�Mrx@��		'Y��ER��	cN�C�f?(A�2� *GGA+ݹd\[�N	��5����})1V���/�TǄe�EP7�8ӕH��i�	qV�;��.�s�E��p�0��m�F�7�8����Q2�y�f�<��3������I*��]��`?����ҵ�?�����b���2�}H����t���Z3�U=���2�1M!{�����p�d��
�H��Y�`�[�DrD%��8ޟVd,j�lB�zP��au�&R�h�b<BQ��$�O�\�|�QD�Q�&Z���yI�������kT^4�JPd��>��G���e��r�l9lm�@eU���B�]Ke�J!�ʁ�=ln��ڌ��NP����Ơ����˯��WÞ%@��$�4{&K���H#�X�I�����:-
u0b��Y%iqh7��9�bhֻƇd�J/ ���/Hv��k?�\B�l֡��A�\�<�&5���%�H#"M�����1q9�a�XI9�,2�%w+����0h�Vɰ�^�`.��ϩ��O�ڪ
��	I��H��� �|\�p��lܨ��x�������G���эj�y��+�����}�H���v�޳A���J�	���=M�X")�d��}	�w���&Y���C�yLX[�&��p���g�d0]�����_���x�p�9���ɤ\��bFb�8�S���J�b�+���?�^��2�����9'�SCjS!dvZ�5Gv(b�>��A�l�b	|��rt���#<w�)�\<Q'n��BrQΟ?-m-�<�D�صs�Z��}��E�I%��?���&cq�n�|T����oF��R=Y����98�Mj��V�Fv5Nos��,���Cr�W����!��q���N�el�+OjI�MSv14��N�8x
�=l��nA9E�'I�H%��uW_��ĉ&-�k!˝��U�/�F]؏yg��Ά����ڂ��_z+����Y���+HN�]�yd7$6����*9�a}�������!-��_�q��'"�)�J�ҁ���z[��s� #w��u�'j�D�>� ���5��5�$�T�K�S��)N^�Ǟ|���~E:9���۳�@kL#���³�! ތ�6'�{��?$��o��!�)�֥<��D�gbpj�A�9�=�Dp�(���4��ߗ��u�CCD�CӴ�������2�>�p�{�ffE�c���H���g_yi�WјJ�V0�^,\�YZq��9�����0�$+y'��^y�C�Q���(
G�M�������"�ɳ8����hU`?��]�?���F*ѫU�Z���,*��Ƅ�8d�	
�Ƿ�qpY%D,P?� ����"�2�S�7%��}K'���c�ɳe�{P��j[9㲠Z��:,i��oV��?R�$6�Rt�ܖ-\Kb'1�\\B[����ƏAWg�N�6{}�E�*�������#{N�'��O:#*���t����bF�^.<s.~��qH:��gg�F�]���x~���-�5�_>��1g]�ً�=[�B�Ն����7�����q>�_q��(��v/S�Q��7^�G�v���W���P�=kF)�{���oOL�w����1r\#ں�T���CcY��k7i�`�V�v���w�8x���Ed�R�D"�j�����6\��[P�َbQ��H@d��h#���3��_"$���*2:�s�x�'{�PWnޮ�m�8	|X�����^��v�¤�c��5���+�(\�������B]�(=�K��,�u�7]�����Ï��:����U%�kڊ��]9��Ck
��19t	\��d<��{��W"��ᴶ�84���8c�	ڦc=�['RQ��h����p�e��o���Ʊ��VU�2��"\�,�;�9�CC��3|��
bbh���j�!{�l�, /�V��@���p��=rx�(:�Z +'�|^����
�z�)�*�U��ϠN[A.�.���9�koŸ)��%=�l"+��%��?g�D������!q5��E�o��1U!����"a�_�x�@��Qi�w�ix@�蔙Z�9�!k^U�qG�\���v�"&�[6ۯ���x�s���#Ͼ`R"�O��1ԅ{��[d����S��{�U�c���:����1�G�᧟�$(J�KC�X���)
��VV�jŜ�ͺBHm�=z.��r�k4�z�
-��{1s��8�f��C�<�P0�޸��F"�>\p�<,^�%~޾K�Y�&N�%7o��Ux�$�ءR�e�h�� ��`���g�}����AȢͯPvM��<��5᲋X}�(�F��=�=�Z�����V�v�����[�K˔��*{���>����f����&��@Ήo�n�S���^�D�S��[���˾�'U�M.U·�UFp��)J�W]=*���_,Ô����p`W�6P�ދ���rԏ�C�Q;Bb��b���%jУ��7������Fmy9N?i]���S��F��w�b�v�>���!ή���/W#!|t��޳��,]a�:�H���b;Q&��������߀hy���h0�����O�5���?�g�}MY�Ə����OƉ'%F$A�(�����I�dw�4,L��&���?��>������	*�"%���DM���Bv�'��0bD��^a�6R�ܹ��R<��kp�4��(JTQ��YG��$�B�uX�j5�	�/?w�>��u��9����S1�*�dg�"ޭ��W^z����~z�s���?^WW���=]�y�{�q�����a��c6�/a� �;�T�XO��*G��'_�иu��1s&�Ve�:l�d�~\��m�r��&ؐ�`�~{�>E|H<B8���f��]���{���M���\�����b�f"Z4����p��3�δ�~�$�X�-�C�Kj��4�<\p�|���w��t�x�Ut��?���W�E�pí�H�ӫc��-8L��!��$��s���	���r��ؙ�5Ҍœ9f�[�)���4���f�VU!1Ѝ����/�ݏ<W؅Ik��a̜~ k�t�ggK'��MR4%���1e��H��a
w����`�bTS̩) ��Cwߎ�� *��-��{�rǃH�r�]�?�㯣�D�G�8�}�#자&��t���.Ԕ�%id�;��_~�Y�#����n����e�<t?���V�A���1�5~$�>c.�{������#碬<����}�L����BTF�P1�k�:�C�]�E睍ۛ0aơXp�e�n�R�OZ��1���K%J�c��������O�
IPPֺ�n������8y���圌�֫���O�P���}'*�w��o/�B�QPŘz��q�W����.��O�$픔$ނ��y��m��7^-Y$I��c�>_��^kb۸��?���h�7ߎ�r�G�iT�6 ���oW*�������}�#9�8d#N>�0�:�X��:q֜9x��7џ�jh�����30����HZv׿��֦V$�d�����^��߭:�Ϙ�/��Y�v�@0L�?�4��X�M��쪛4��c�6m�58���b��;��x˿$\j��FJ,�_$�J'tRu�/��3�Tm��v[k��x=���"�}a�-��k��X���=6�9�@�X���P�P�/�3�����b���y��̣0u��5b�u��で%��"^�x�t6�])���k6J*�D���Htr�Q����L�iE�d�n�[q��)��E_k�N=��z^z�~�s��S>��/X�Q�x�0�w�X�y�fI�.sN<^�؃�,N��x۽�����������c���8`�TH�)�V�Q(Fs��מ�M�����^��JFt���W���/9�~D�n�Յ)�Oƺ�Z��$��s�=�'�(�g��mW���$uy���$m���n��Y�Sf�;y
�%�P'q��%,OJ�n�'_-Ǜ�-�T��0/^����r�$�9�r���� R_��EN�V��d\Źg]�p$��Ǧu+B��r˿�k��8[�Gu4}������q�E�ٺ#'��O���ѣ�9f�`oN)�W�x[�Bȶ���j���'��:�32v�8���|Ĳ6��Cڵ�����O�?�?)��r�{QW]�x v�HaP.�^Bmtv�aѲ5:%�t�B�SXy�'�	�_�I������)2�;�N5TW��n�G�~����\�D�, �p��ރ�?oĤ1�$�<,}��Ds~1I4�W���J�=�\�h�H.9�I���|N>���lډw}&j�?Z�iʢO����N��"��r9�\�)җK�5n�HW&����?Bk�0|eU�Xe��%ULKJ�lԥ�6����~#��`A�t�x�����9D$��'3�K�����5���W٩#�	v1��!�C�|��|_y}	�rC՟5�1Td�p�2�9�x�#+�D}��S�j17���_D��D�b3EF���~�{O�S���hJP*>rJS�%�p�azY��а�neG�/a��7v*�}��2U���X�8Bz_~�Y�
�$�Dcv��O�O����S�BL��L��~Xo�L1]��5��FD��Z�c�?#�L�Ҳo��A��Q�oG���+s�Ek1I�jq�巈�i�=f�N�?��z�:a[IDh�I'pYq'��ڞ�u�o������D*�--/{��:�����O�'�\=�Ԑh�av��N,U]]/��.MM�_i��Qo�֒Oq����qKHT7���bX.��t��ò��<�2��bL�(m�2oWK���8��/>WVՎ���"�Ł;���p(�Ͽ�RH#�2V��F���J����#n�b �)8�$y+n��x�ʺ1JK�#k͂2CR�<W�l�)I[j�����=ۺ,�k++��S�ï~�p�t"	��(�_�~9'_����s:=��k���(zP��Zy�hU=bb8�.
6�%ʷ�%Nh�W�c��J:���m�UI��RI��c�.�iz-F�������́O{O\����r�9�F"w8 ��D��K��'���ZҎ�^Y��J���`w��N�l���ʋ���>7�O���:��`l�e����`��9��"Q��J��j̘>Ei�?[��tn�"���6����0S�D\:�
�����]�Ćb�+/;������LI�ܡ\\yI/Gh�E�V��y�d��6G���SS��V�6r�VH�����iC����bV1,�����-�VD�G
�&����c���hN/~�Mv*��a��h3'S�nي�S�ԙ�����ȦݪU��:�Ő����rٵE��.�P�E_s���X V�]SS�hI�Ϧϯ����$�+o��%ʠB<�IX
i5عTFuWhH��˾�5��Y[�������\�2�!���,��q��K'$�[��K(�(��%�1�z+f�*����H�4��۷�l��w��P�c�" �kIm

�3�d���	I�|���� �:�W�""��Im�3b$��F��ce��V�g����j���a�*6�lEU�X�9]6C�]��c�Ic���;e�%R�S��Q�.�b#?��y�.@����(��NY_o��󞲝�$L��ml#3M"�B�DЫ"OWV�8o�zԠa'@M�7.�X��2R�3]'#�BeEX�H���$p���u���J[�.��v�t0?��\���Vp�H�V��@�d2�S�G��������h�v�â*�|@k
�ry1�K��~0�.���G���F���y;C�j�	�H��ϩF�7����]i(f�&�ۃ��>44NĶ�m��$}*(!��er������`��[.�]���*I��Q�ZY���8TF�����noR���LJ��#I�� �e���P\(�A�VO��?���+c��R0z#���AK�abk�G����B�J��h��� �vi\��Q���_�H�re��#*���Me0%�
�ya�J�R_Y��1-$;�����b�'��1���8I�#V�d�,��l�~m��8p�<G^�r��ȅ�"�����li;����Cj�6�W��k8E`�W8^��6#g&87ğ%Y����)d��mB"ɐ�dMh��t������a�V�p�*k�a�\���Ϋ����=�n��KI�#S%gu����U���D�h�"�^�DA)	8V��L˔�U�gj8�i�����|]��R6,%Qؠ�w1�J����qj�E-U<2�<� Qu׮&L?
;�Rr_�1��p�U��؄�����"0Z�fq��N�#�z�j݁C�,i�*IM�j��$��K*:I�ny���z\6ū�e���w`�ĉȧ�CQ	��F�M�T��ȡh=�	1xiy�u���5� ��<�~b�%!�AD�Y�bx�P�ﱺ܏(uB$:(���Ǯ����_.iM}�����a��֞�d#g��rxe�3r����Fkg
vθrZ$�Yr�{�F�rR5U���E!{/Z�y���X���ɡ����䗟�x��;�L�Znz`���z�˰ �&���rY�Ց��eJ�Iu���~U&g{��;�)�:(C�#S��ǂ!	A����>X�1I�l�*��
�E�wco���b��C���ɝ�j����#µ"����5�1b�4�jCeS�/ə)�(^5��G��QrҖ�8�st&V�R7�Z��Am%180ԯ�A�HrZذ*�#�9���bۄ�y�Zw�`�M)�y��
n�v|��P.�l��ѺvzHgHk$�ʭB(wO{r*:EJBy�^���A��rIK��0]�d%�PW��*�<��ɳy�R��{�ƒH��:[Z����-ۛ�{th�J�P!����Xx�uzt^5�ެij�V���t�QW��e�gd6w�!�ꠜ#!��^�:�0�J��rxOT��A �e
�^���oLvvK���$-�w��iS������p2��dr�b����&g����9�<��v sr��m��b��˞JJ�R5�ak�`�{�_[]�q�j|��cDe��)���f�qО�8��iJ�H�c�re�c��g|���p��%3؎[n����°$`�o@�g �^y�2��C����U.��b:4F}ا�J�h	��9��pY]Z�*n
��V��F�D`��p��EI��*��c�q3�~�*mQz�^��Ȓu�G>c̨z��_�"P���D.����==��N<�M�Q^S���/�+\��,O �K���*9������!���F�M��I���D"����ܬ�LM���X��8�D�$��u�QX��w���s S�]����L�ܰO[�@�zl�C��}�=r��*�>6}���d��x�.�ˆWH�0�v��xqq�_�^e@5ri���~��jg�8�_��J篒��!k�؉�3���'�|��Ͽ��R��{��7��s�ᴓ���=��
L
xhon�)'� �C.�x�X���� #C���\�X7���<���#� ��99���h�Qcᕨ!K#({�IR��
s,҉m�m���c�8{�1x�Ű�a���DVVZ>{���IZ1�`�d����1�?^�.8�,5󎙁W$UKQ?
��,ڦq�ɳT��bsc˦-��Tɿ�WfqZuR5'Oe��8^{�#Tɥa1�}�)z��b��[��_�/����69�?�\�1#OD{K�;l:B+�ổ�5�c��3�#��VT��3�g@Y$����nc�q(���p�ygc�GK�h�"�9��v⤙�`�	c� W�}����6�b����n�Պ=FU�/���^��r�W��#�p�p�� cS�u�֣����,�LR̻x���Z�q����m����*I��ʣ$�봹e��i��E^�H8Z����3~�9qTz����Sx G�9����;У|��c? /��.j*F�A,�-�p�!�$�N����<�ʪF���%��F_���0 ~��i��ǟbGo�T֠w�'u�V�{S����3��W�GY���!��c�x�*ɹ���3���O�Q�\��Z��/8m�������W
6���`��݉3O9Y�س�;�o؂u�~������*mY�,���9k�� '"' �}%㠱�dC,8{މ�^��*��P~ڴ�.�..�ƒ�^Sz>���ŋR������E�����n=m,_��==�ˁ�TU�c8Xk==޿����Q�(B�x�����O=�h���Sx�)dd}���:�x3��
`��͊��T���a���/���i�՛���+��֎+V`�x�����۷��a$��bxw�gp����� �'�>�$�[0O��	�_r^CD)ֱ���D�����-�ƭw�'�VkQE���,��{�VV�*�D�DU�,��O��mr��5��qNT��xށ���ۊ`�\E��B\><��8��3еsΚ{��}����]�T���Ӂ��=���I��W�G:���r��ȓ��%�c�ۯ�B��.�
y$B�&K�[�U5���&&�8�֮�۲c$juJd1m��8��K��yXR�8��֬�ſ�q�S,R�,����\{����jL_�yߍA1">yn���7�tc�'K���P"��]��
Ͻ�:n��:M�Cr9e=��{�B퉪uy�Z ��/e��)ғr�v�9p��ុn��og؃��~���I�~��-���g����d9�N�#*��y��⹧���P��](��Q����*}�TΆX�+.:�-�Z����j�}(v�؁�q�௷�"�C��|dp�޴x�}�/8]�G'N<�PU?':��4Q]m-:��/*ѮU��:}GO�����=u����鳏�\���K�;�lPV�>^*QB���	n!F�UDvk�Y��5�d����Af���n�Y�=}A�T��ϗ�gE��C<�ܤ�a�fxr�=f\��c,�?},z�Ȧf�V���S�?g�J��2��EkO<�
.��x���|ġ����B�x��.�����A�WS���;T߭X�}�'iZg�9^5[9��&)	�J��
,���ݴMF��^�a{�����h�5w�x�!IG�8p����S$�FR��7m��u���U(�B����'��1h�����{�|�!$dݜV��������\�\Y��Xr��NDG��h1��~��'�%�<pox~s�6"F�b)����~A(��7�E����O������S�Q�u��ݦ�$����X���rYCZ�3�jf��[7�?�n���òCή��V�}[�2�����s���e���t�l~�DHK1a�H�%iL~x}4�Cq%^"�k&?�$R$��ԤPRzסBqd#{���p�e���ݢk��H����V��.�#!���&S�tF9^o���z�	�~��K�Ė.9T:{��ؾs'��.ӽc]��e"�Y���z�t����i�]1RC�������O?�rEi�)��&�G�e݈���p�C��xCb�2����,��"��G�>�$��x�K��|n��$B�������l?qz�Fb�8�,�s�y�|�r��e�c��d���{�Ҭ����G;���:N���~��>��n9�I}��v%�oݥc*#9��9��ƨS«��xN?er���$i�X�hE6�A{�R8�a��Ճ����
:t�V��g�P� 
���S۳������FY�,e�\�+���@�xŇ�x����*���ߏ��ݛ�p�oچ��Aŋ8346C�2N�a\�a��b'﷯^R��:�$���ү�����Zmg���/���mw�4T}�'8�#���y����_��\�V�Y0Ek�;lNT���S�c�9�R~������-�v|���ʹ��8��ڮ�.y$7����?)��&����LA55�z��n���M�g�����*:l�H�'\���?�ܹs�5,)��^����K>�FNX98�GxC� y�7�<�ݏ=�æM���#��ޅ4��t�\h���	���^yӶj�����S��K��e��������-���Kf�4>o$%�H�ig9�d��?�c���a�]�c����4�h���7H���)���-rRZ�/,Q��~���Օ��v�^$�o���GK>�3�Wz^��D��`mʡ"+蕈�ko��fk���0�6�l�)ri�NiK�#�����ˮR���.�����_���>�3���|sظ|��m�%^�P�WgL-ª_V}I��5�HO��*Ǝn��"��o� ���HEY`C�_�U�� �΢B�߭܀�뷠��]�%���o�c�O<���E�ڸN�6O�=����+o#�s����1q���y"T�2�I�8UY��p��_��~�&g`�N�*���-����a9�$#|^�L� �sIYrbX��.�����:x�ux���1�n|���͜Ci�$�=ɭm��D���\��)=:�j�! D!�'��Z
�u.[~�.��y ���{��Q�$ȩ8���SS4�~:�efWr3����-Q�c/���y�I�[�}"NYy%���c��fV3��c�Vm�e�.��܂/��Q�Z<�3��8��"�-j�l0S��_�1;i��J�賯h+�ғ:E*F����ьj��b�*F�֋���dK��Y�]����a$aeA�����Fe�������h���� �?�iW����$-"<5p��;X�PB蜒:�7�/�����N�O.a�l��N#S�X�I���g�&d�����ˢ��v�f�ZK�F�ͥ��o$s�:ς`Zvw�
N�Hə������A��Qn�|�D�>R5�ľ2%J	k�^���/�D �����pF�b\3�E���pH�{�@����zz�N����Ý͕B,�q�l���
?	v(����K�m��M�Ei.�ӧ�.-���6�"�
#�h1sSj����1�CjɤLGIE�94감�ޢ[^����5(,t���\ވF.pH"%�ס������DaQ�]ւ!g���]@[�,�f��MCU��%k���(�����#��%��H�R��I��d2��l�j<��:dƎKA��f���ٕ��li�]D���S3�kG�[����ҨyI:�D[�Ã��Ӝ��:���M��Y��Xw:I�y�4="l-�kTԈj�C������ ѠO��%+�FǕ��"�["/z*_I���5�΍��d�����9x�#��++u`�h8G$�ߗ��'�C�d?(����X>;O���)/��Z���g>���9@H��[��v8~5�ʁAt2`�}t�̜�<�Y.��6{Q��x��Y|��8IH�C�C�8Z(p���6��e����B�0v�r3�	C���3$���Ѐ���X�/�^�������Ɍ��8y1�䡑ˣl�b�(ɫ�,(�	9:�:�m ~*e1�#_������PU�F��s2�Q`�0���Iu&��S,�yu *�aI�Ĳd���r��&�(t���YiC!��X���$>H�JV�v(WR���[��b���}A���d��]�jY֪���n䆍�:���XXWф�L�xxx��j�&��R��X���Yٯ�h���s���ɭ�)���LZ�I�"E���ߧ�g�Cb+*����(1ly��2��qYDָ��� ( �Zе�"��"����x�:�<N���/.�&��I,�CV0�5�y������ᾐk��_,�K��Rz��F]J&CZ��=b���kA�̌R鹑Hh�c��AC%�/O����jIO�j�
J����;�f���3�[.��J��9+�
��*�0%�,���E��g�� b<I;�����S~?+�:�����L%�F���K㖕���5�ۅ�ݤ���?�I���Q��L��m:���c�p���Fn��a���O��*���J0YZ��2���1ԓ�ls�yJ�vf*�7���ï�Lą0 ���6�ץ9�M*�F�D���]#V�΃F�nM#A
<�Ga	�x����s�6q�9� .:ܚ��J��D��ȪӿY���z:���R�Fc�(�[Qf�c
vr���Diϔ�h��PFe�E����V���!�H}Fr�|����r��>�d��OX(�W���4LP��� &5$�i!�0eĚR�Y�+�����j Onz�C�jh4R�%�"�Z9�0���f���|�<R}��w�c������krȓC�%�����LP""����$w�K��Aa�"�JqP����<���=�����Ԇ#���02r��C�J@�	޺:�$M,W���[��+��H8yȇ�d��
}
)fH�u�NE��H��Ң�^0�"2$��&88h�����'iTɿS�g�M�ȝ�ұ]�Q,�A
$�O�ġOU�k��$=�(ӏ�R�@*����I�C�0�Vm�t��8܎=&L@yy�[�4գ���da{��^�qE
D�ȬfD�^��zS����~���r��P�vdǢ��F�������3�jo|��9�>yo��>�(GnJ��U+5��X�X�V��Sy�!G��"��u���T0*ux�kW+��!�Ħ���8f�a�S��b��L�F{q�9g��<���~�Z=z��F�����$�b�<��p8��)hg�i�$H(�zq�g`̨��)�S&������?�G˾��T)�С��(�5e��e�����+Q�W֠y�1���Jj���<��㰗�3�9�8�d���E�v��˯��@��X\�	U�ƍ�KDґc��q�F *��с�0ǲ��q�|�b�����kZ(Q͙�"=�PO7����ps%���]Z?��{䉧��Tィ�ba��j�K��mߎ?��<TTV��y'F���R��K��k֮�$զ��(J��!��ebYS��'�C���xA	f���+�km���Q��(ȳ3�Ɉ��X���{��X�~²���n��f|��rm�8Eb��2��|L$�q����٫"NϚ�(�ER��֍��c��䂵P�dԓA��'9��M�Q��Z&Q�y��"��T�90K�Q4���dF�1cځ��32*`{0̔A�Q}m����pk�j�HĢծ�ApYOG�D
���5k֬A}}�z�#gL�]?��LI�T��!�����r)Z�q�Ǣ��J���Q9I�nl��@?�liò+Q�K��ؒ2�&i��R61�C8sΩU_����������<���+�E�F%��S]��I�#F�R���\�];��qd#�q$cCjtgL��?���鼮1����vm��{pǍW����u#4������(�|���O��_���~�
oeZ�Ք�n���*�P&kT��+���L�B��y�!\��K� NE��n�F΀q�۷�ƫ/SIS���(�s�Zv���;�[�\�Y14�̥��̣���?���'�+�>��DY~�S�#+�p��þ��9��߫�|Q}؍�o����#�G[��^�*& �#�p}����]�8o�g��>c�+u��� ZQ�ş}%+,��A�)�<�������-���� �ף�����b�$�E���\����j�YHdo��v�\�����,�|��V=��@$���BWOj#^����o~�(�ө闦MLi$���k�����Dw�!��$�8VG������\��q�jG)��MU�r
�qX�w(�<��XR�ӯ���
T��\-a^Dz/�X�NM�T������;>s���!H��ax��:%��V����ᾇ�E9�b��"5
נ�6�5Q�c�k}��R�b����?�$<���ڮ$l����$Yh�w��*ñG�@r`P���V	���x��^Ԗ��3N��ϼ$�k�*rD�'�qh��W�a!�D�Bȉ���~:�VH����+~�[���(�W��ųne������
8+��u�c�t1tH]T�@lŮk���ڊ���zQ�F�;1E)Ab`�a�����������w�*0�<�?�^��j�%��!^5�����:���Ė��`� &��������,` ��6��T������xmc��RhkS3�QJwJ���#܃o����K$�s^�Hr�f^r�o�
��x�lTBEKBø.y�k.�Ͻ��J&f��ޓ�&x0��ށ��!�"T1IA�9"$�R��,�=�:<�����O;��z������x[�q����!����p�Q�L�{
�^~�:!��1�N�M���%�|�V,q�b�Â4˪���D.�����-�E����ꖖ���Y����r����ZlA}����b��z^���'��[�p�⺜\�%���q�}sv�A�e1eS}�3���ŭ,I1[�K��M�WB�1Æ"�R=���1vRޑC����\w5�%~bf=(ޞ���޴h�Esc=.8�t����ȇ]jڋ�ۋ��������w��ƶ�aqj����TG�3��K����O
�`�b�Z~��G���U���I�h<ŀY�pě��}�A�|�=�{*m �+y&-8�*K��-����v��q8����Gp�1Gc��u���m��T���.\(��0é����c�J��>T�1+�����~1^�s^]��ZW'�����W�G9B��*��ֆ&��|�*�M�8�`3K�p�i'��Ͽո��\&ϙ3*/��P ���b�e���������G�E2�)݅�μ�-� .o��e�R&�6��M��K���_��
��Q�f���(��mx��;q�O�9+B"��s@�v��Ǩ·����>��v�fp��OɻI��ѣ����M0�|��H���kB)�L�t^�Iu5���۶���qƌ}p�{i�}(O=� n��~xK�t/��=�&q�M��Z��0�~�n��)�?l,f^v2�i�]����������jk&���q��w�r�;�Q:j<�y�{|p㽊��
�:���0v8�(�:qх���+�L�e-گ�a~q0���e������W�1cFc�쫑a(a���Õ��YgV�@½�x��;��y &}Y;���M�*�s����i�y�)H�zp��[q�e���(�=L��}�->b�d/[�'��}	1�(-���oc�	�I�x���%uc��/H̶UQv�������A���7]�G�=#�â�	�3%�}����!���t֊���L��NL�0��|���~鞓��x��6
��k��ˮ�y�<pT��"��5�s�\eҦ�ˈ�r\�epGj����,�q�}�=Y��|�x�i�uU��{_<��[�c�Z��v��t�4L7J�e��G����S�h=v&%S8�c����J�����d���M��ݧL��� �����K�ˢ�$L�&a�Ig� .�Xq9���8�E����g,X[߈�O>|���V�.xK㗈2�(�"������"�@�H�lw̹�vkM�2�̼H��|>@.�������:�<J�{]m�#ԍ��[n{mrP��rJ���W�c�A��:X�W/�>�`����ZF�
������g�H�S��Ja֕�K(��
��_����O�g�qÆ�F�놼�:�\��$F:�JAA�@%f��6��>��ȼ�p��W)������N�g?/W2#&�(:<��J�=�2\t孲�N����Y���GX�n-�8�x��Y�z�Q�S�٤CkY���N?�@�
��w�y�Mb�혼z�_{�K�K�}�Iǈ�@O�}�t,[�IG��Z�1���� ��b�x\|�b$��y�dk�N�<�><pϭ�gb:	z��g��ǞE�4�Y.?�,����)-|a1���Kc��A6v��ɧ_ƕ���h��ċ��<��"9�c��d)� ��-x�����+�׳������Ko���c@&aK��b@�ʌ ڐ̮ ���zBeb�����u�u�L?S'���͸B���E�%�tHHً�'M�3�-H�s}I�Gi'>1y��҉U7J�;�{�<����`r:��Wc7f^w'�~�n��}��A��+�!*F*ƌ#G"��<��-;������lX���|��/x���S��+���`|��R�)���\b#�ˮ�Pz�y�Wz5�,u?{�3�u�����¦$��o�I�ܕW�Tf�Ǐ-��P�{�θx� B�sx��%�"�s��܄q��~K�����ۥJ�p"mv�Ͼh]��YSX��C��|���4 !�Y�R����DCu�I^|ml��RZS�i�n�(1퇟|�iS�T�r���`��!8���nN�v�p�z��p=�=H�}2R��zV����-�<��Y��z�����8>��������S�z�;T�_��2�PAU��)q.	k����;�}��JYm���jˇ m�5��x�Y��5k0��L�d:f�9Fν��E���Q#q����;��Ǵl�%K}ފG�z�w��a��| �#/��Ii	��%b���߳��d�]�q��j�ŝcz���dVB����8�I�T�)Fk8��	�E!�U�Z��lT��v���\g� �5���?���>1���L�7�4�g�Yg�V��cN��≅O�;nT&7��B���Xy������b>~*~Y���]%
f�/�x��_{�|L�UD��L�k?�ը�����y��G`�02kvi��V�8~_Y���X��xq\�"C&��(2��O�CYE��uZ��r���lVTU��7a��s$�iUD��ظ�.�s�<����(2ɾm�F�Z2�bן}�9��:ֿ�z��{ű$�%E��~�|�D.�^p������bq��\n6�Ț���.�h��!���������c�ÏKy=Z�:��R�(��7?�bi8ɪdu��~G��E�\Kܖ�Cٛ�*�����*��'��@�bJ<�S;��]�:�	4�dq�1�ҫ5���.�u�5������EJ�9���9L��@$���"�t�#�k��D��2jrbs8������#ɜ��l��������X���]B	�\����3&���r�S5Ll�H��bBD<�[�9ٍ�-�;`׾ ���15���/_���M��%Y��Q�` .�"��\������Y�C`�f�);���w��?�b�Ic���`�=6�^�<+)*#H�3J���s"��B�C�nn�a��*��ks@2=((ˋ	%�z���uM�(g��AJ�׭Y�\�z�

B�:�:��K��O�M�)�/����ߐe���-;�N�\[������11b&�c^D?�a.���,��6m����(Ek#u�]*�H��cB����r�F""��Y�W���1�<{D��sT<������eO�r}8<�!��X��o��M*\�=�"C&�����z1��$��IаC�/��@Ό���@�%%0y�r7�>2�d���?#!�ˌ�pl�ʊ�$m�ë�T$Cj۱M�Qò&��
8�;�	91���$�MjK 9T�/[ntI[�l��P,'��"_�G���T��Mny^"�8{��AX�b��cI�˺-�|� w�hgg���1�`��5���׊&il�xխ�+l�8�].XR@O8�@�M͝����6���wS��������]Y��bͲb�l���$P�L��U�战�i�l�fevZ�z���&('5ڣ��7����փ��pJ�c��	fZeC�|�����a�@�x�M��8|���tl�!��Qސ���_:�Ғ�'��Cl�l8G���9J幒P��Xrc�n��ZYCw�19���F٨�� Ge��$�$�����c`�)���~1��X�d�Lf��5��h�č�&{GX���Bǧ�M����/��o�%�#�wRB2��mgP˳V����������24Mپ�T�a��ې��/^2*��\�Y��9��s^�&���7[]�Ύ&8K�:��a�B�h�*K{ť5ڰ�Կ�bȽb3$���5�ż���в�68�M%���c��=�[���)�U����,�M��]�R7ס�%�Dd��81��QK���D�|��'NP�	�Ɗ���Y��F���2?<b�9RBF��ݢ:15l�$Q4g�8�l'�����o��g��|�11�DTԑaKz�gj*J1�3�F]�P44w�{����7l�((��V�\p  ��_���,j+F)�e��VA#�}q�G�!uR8<Z]S��p,r1yϴDf��s� bS<+ٟ"f�c���\`��8k� J���w�Nm� VE� �xU
"�dCKZ������_��P_OX.�,D�][Q��X�s�ŉܤN
�I(�e+�X=	`X(�����+�8u'�� J�rZ6���J23R�usX6�R�y��(��8��D��Iȣ-۔r�w���Q(�o�L���(�$7�%�J��%�~Y����`�-̆�SR�u���4�C��׿�%d���L@9������5b@�*~�R����MI�᭒'��sI1�"6���(�d��\bH���A4�E��~��ě�%<��e�P�"(���Gj C�*�r���1����v�g��.GyS����
�cy�ƍ�Y�L����eS�)�A���w��8��ͭ����\�twr��R��2��L�����0Y{&=riǏ�æ��t@l �n���J��$1{�&���+Y2�KPΓS'�'���[�"��NZe�\H��+/�Y>��6J�:V@�W��)vȁ��O�#��.Mv����?E%4�֙�����Z�]>)�*�2[:�1���>u�U4B��b4H��GM�%*-+V$o#�1CQYK�3�q�֮6�w�IX���(�`��^i�d0��V�˩�g��gw����^���S�ɒ�P\\)wR;A�.y���&̚y��4E%�������AM��>�I�8|�~���;1����#���hŌ+�3­ҠA����raR��a�ٰ�>�(1�U�?�Ջ��Z%�2��f���ȯ�!�D�W.���l�w�4%%!��ႊ�E;��̣�U ��v��6l�x>��HL�kJ.�����ĩxD.=��������T��hcF����C�l8���������9	6���������6^6���3��Y������b���xS��Ų
M������-�Ɔf%�a���(ĒWg�Nm~?�Z��"y�kq�q�b���b��=J��ZbY��`+1`Y9���aٟ�� ��C�;���wl�G�{<�ښ�I���*R"��x����y�'��c�[��=5	����l�H9����Q,*���K��v�RA�;�_X����E�s���m�1v���15Y���"�1����j���6��#���%?K��BOLں��qə'�%�Kh`���P��;����C��)xj��RW�����w�J����v��0�=���c��CB�#�k���ى��2%��mŉGMײ7U����o����T���+���q�h؂{g]�[n�G�9��.��*�>}�=���AvaK�V��I�D�����+��Uk����p�gaxu�rv�?JB�k����n4u��M��J���r6$t�ɺ��hTm9N;�@���"�8�X[]���oP�y��(���7i��\�_V�������8�\x��d�}{3%~�s�L���i���^���ǲ�u��AVy\8�?x饅�ik�+��5Wߨy�3ʗ=������W!k����m���=���V7F�oE^P��w?��uj����g_-��'���.9l��ڋ��A��x����{�	h����a���������Ack���O;
�&67�hU�e�|*�+�s	�{{�Z���O̻?`4�Y��yl>n�e����5k7���'������>��w��Ģ>��Ԍ�)gES{� %z�q±G�Ͽt�R�Jz�sN<�;vH,�ζN���+�jVy0�x�-u�~��A�g�$�F#���[��p׬���y��h�"l�ވƦ���au�����5\z�9J��a�c��zp��0k���7]���:�Ia�7�X����0��?����3�p9������_|��ͤ�_#���i�(�Vy�p��X��g���?7j���gz ~_����Ƃ^l~����X�5�B��.����,n���K��sNGFB��t3�9�~�1|^jK������$�$��[���o�J��tJC���6���`xm{Z1��3��ۏ��;1u�%0�޶7&�*T��_xu#�h㛪������S�g�-�&p��W���;[�4�Mau01��g_R�hu\{y����wK1�J���rs̽��oB�Ν��>��с~���ᗕ��`�T8���b ��.��l4o܀W�}�k7蘿�i���T�8*A�j�|��(��g�g�&�(Ƶ7ފ7^X�XG#Ɗ�|������h���;���Tw����΃7�.n��pz�������>�OD��/.|�۷
lEO�N&;���1��7�AMD;�f]w3fϾY��<>�a��A�ь��Mr��ں��SgL�p#�e����x���>@<�ݝ�b�����G�\�,��9�$!J�@o��%N=�L?p(v4�`�ڿ��7������M���������@u�*?�"	�~VK��o9d�=p�!H�mZ[��OI���c���j����!+���o��.���\�R�W��a{�(F֕c�Ƚ������GdcX�2P�^[;Z��q��i���꒍���@U����~��ȉ]/���yt'-q0QW<�o����=ʘ0�1rH��5KQ�ˏ�:��Y����9=l�@)�}y�}����8`�IڞO���.1����
�g�t����00d�0���ǘ��T�;yz���	�C���X�PMղ�Z%�aC����Q2 ���8>���{��*y�!��S�a�l�'w��s �|�#����"��9j�b��o��Kϗ��X�N�岬�j�!��N���^���6�`�-���ï"��ah��?��xS'�7�6����|���0&�٠�J�U����cΣ��+Ѹu+J�*$$.�K�t�R�a��_|���k�\���Q��a�aP���y��K΅���
8-�{�8�1�Iȹ_��j|��2A�A�8�������ڃ�|�3	���x�� �4��T!��JV.���A��Zg^�q�M�f�%|9��+���۲��GD���8'���~����4�CeV���|��E��/֞���P��>mҼ���]����E	��`�O��vZ v]~�%�x뵰��!�ףk,�ĺ���{��۱�Q	�����55n�%��O.DK�@1�rm�R9�T$�������Ü�ga�م���]�{Gސ�'�|��o.FPb(�KR��Ox'��?��\�LMQm��c�+�!��d��Ͼ�^90�$���}V�>KWw?�,Y���8XG�����}L%���h��1#��+o�pI�)�X�l�8��Co��%�v �m݂Q#����-�L^"q%jh��SdL6R���Y��j�`��)��"2Vvl���`�+T�w^\,��R�\언\���gLV��R�������8	��p�"���~����T�v�\X8K�7f,�yB~TYl�L5X.���,(��-M�4�I���l<��7-FO<����FN[�3���(���}�p�1ε+���a��iw�ϵᛟ���Z���d2g�,J�S�&,|W��h�JZ.!��`����5�>�8<�� %��)�9�����\�)q,��[�"��ݱ�E��c1����b,r:��v�5�����.z�[�rf�pU���%���#F3��A�����^�O�yu<>�VnMY0�U��_��y����e%%�x��%���������7�@��Mٳß�x,h�����'�`pgjj��f���vò�+侼��A\)��YI�z��&�2|�=qݍ��.5��x����Jf0羇�w���7���i��Py%^~����R�$�{I��ehmk@kg6nn�e��֯\����b�:���҇K/�3��9�A	��\Hv���Q�\kI�P���Y֞6���o,�M��P�&YC����;#a�?o�?RbF�5b��ۻ0j�D,�m�}�ET,f�9+/޼�0��FZB���?�9`_��FL^��~{�K����?�)���R.�ʋ
�Oo�hR	��mm,����np��q��#Q���AP�,�ϫ��!���O�����V�W�;Z�Ջp��ێ4�����!�\k\uU��H�e�4%/�~[�}�Vlg/�Ȩ��OF��ݏT�Jp���%�2e�Z��Ŵ*bd���T.��`CG��ء	�7>�Q7��}���VOB��\���
A��er`�n���Պ`Я|4z	�J?X8l*���8�FX�+FA�ϴI��5,��9������:�=�YUy�h"�UIX$tx��/t���HBY9p:'$���_P&�?����<6�a�O���m��I;A�Dǋ�/F�D<�@Ҩ�������VGl�=&�ޜ�qqۼU��'�t/;"�(��bf��9"3����g�D��G΢����JK���[��	g.^	`����tIK�� �E@��aqtdu�"�u��B�S�� 9�L�CGoo�a���B�i���ťOFb��ܧߒp���c8���$�S�\5J��� OY�_c��-��5܋��#b�N�#�I��a���{�$*`�>$a��<�<X��O��؇�d?Nr���z��_�$)�Y`�o�خ���<�X�l?'�"rɟy�Uՙ��@e���W�m�B�1���k寷��Z�j��e���4Kj2Hd��R�pg��cMi�:xf��=������f�:����Nj�
lt����e�{��-��PLБ9�S���Bªmmb��Zf$��U�sr����bV�AƦ��nm;GC��������_2Dٍ	��àt?Q&&fY�s�R�y�����d_K��_x��2����ݵ�lt��.�Q�-�;���Ցl��!{KTHJ�������f%�VpX���#Wr����VE�<%E���`?�Sa)�yC9 '�禮�1m\�Z��]Z�B����p���u�8_�d�����<?���(�cףӤ�:R������!J:��O�i�@�c�?�2?w{,F��@	�傒$oֲz���/�G�IJ�S�ư��w���%��ܵVԠ�D���:qrV]?�Hzau�Ԭ!��08i.,�;QI�����I�?Cx>�ʔ��?��$�|.����P�K90�z���	6���R� |��L�g��|a�g��38��7gu��&��VTi�G�|^>+��U-�!����0d�_��ٜY��G,�.���Q1�&>-��L5�D�+Y4��̣�m��g54?��������M*
�-tB��P+sh����Z��ٍ6@�Y�P2#��?�L��3��h�I��V�Y��z�$�H(ِYgf����Y0�"�t���0k��i!ъ�0���x�JCV~yK�Г��C���a��*v�lޱ�tv2���S�2:1,q��1�[i
h$�8�Ұ�R��&K��`*x�,������$G�*5���6o0����EB�ԇw*�y��d^�eU��	����Ry�����:���,\J�ɮ�~���Ԑ�.�2(�Iy;(0j1��IK�95�a��Ϥ\3
	���~a�:�k�|9����w�L׃F�ݖ)�3ՔU�G��������yE|=�z:���P�6�)ѢIk��wM��0�#ǆ:�K9-�	l�-d=�
9�=�-���9C"_�r���PN�DQ*�g�:LI��\�H����ɓh)�	�X_�"E����d 夹ͥZ1V�]m�<����"��h0��u�x����f�6�X
MF�7�pC��T6�����$<��4�"6��k��v���'B%֬��ұ~ne�6Lh%��~�e� �H�n�xR7��<Ӽ4ym���c��Z�`U�-kx|��+h�BD�u��jρŰ�f��i��VPh���H���T&'����jV���8)��n���A�g�fL�[۵ׄ(*k���%�w:W�� ��\��4x5��8lF-	��G�X�l�4�<�.�G/Y$��2�����$-�+���|Nw[��F+�jhUՂB��C���ƐG��ZV�w"0y!�u�|R�_��h�f�Ԛ��]f��NX2�����p��
����j`�q���?W2���ԩ�P��:�l zG�o�56`�Q�N`>@>7BBi@�w	���ax�p
�7�Yʑ�!����y����h�!�$X�p��pƥ�ϵY����yinj�qGO�>�:(xeb�j��v�*2�p��|��9YK��ӌ����%lv�]������|���)�g^ٴx��g�z�/��f��Y[��N���U�I\~�PS7Jsiԅ!��I-�ܧ����;��sQZYslIA=����=��5l��	kk�B%���t���'�E�C��]�__��O��?�*�)��5KnB�74��*�q����x0��S��dr���8��1c���.��X{G�@�VJvK,���fdG��ŨuIE3ټL2�����*���\VV���/�@Ye�6��C� �l.��������u�,t�ZyF6�쐐c��5�I���h���w,!1�ǎ��f�3e"��AGK�\��lRD�q���GJ˴\���
G�㤼���b��d-Z5�dh�?GS{V�\��ٽ�#�lz��� |r(w�؆�o�%��|��]m�D����oCfYlk�[�ДͲ'Ņ�a�W���;w6��r��{ �w��<���dd�Y)�.eZ�\�r�`N�1zT�̘���zF���s����=�#F�Q�Ng�9�:e�#��x�I�}��w�H�\�n9��0n�5>�zQߔ<�jظ��3��C��ϡ��Q�h����S\�%+~ŗKW�ޔ� GLN3�aY?g��|����g])(6�r	�I��&D�*E.��:T����X����ɟ�&?��C�˻ĵ����,�V3t(N:�<p�t�~�!��1��d;y$�կ�.;�]��^���I�8e�d��$�p�=(��U�P�M滈m���ۚ0�����"�a#93{����.�٧�����(*�T���0�N����&<���rV�`�#�~xq l"k�3q�g�'�z���(��KZRR&Vދ�;��ׅ����r���v���|Ig;���?9`/��ø�^��9-��K��y����R�)됑�3rh-���f�� ���i�V�Ho.�[�J��݄�V#�!Cz"��\��]���X6��Ҧ'�F�ǵx��e����'�;S���;���#���E�(EI϶ܲ�2�����;��e�F�2��gί0��%|��b�ȡ
;�Z;t���
�p�Y���wއ3P*d�x>_��`�IE.?�2�ww"&����D�ihv�0]�����<��@�4l4:��xt�l��������*Ɣ�dW\|�~�������@U:��Ұ�_����b�6�T����ɶ��q̑���O�D"oHE������lV�����=�5^yR(���f�q/�1̽�6<����UR&E�dcS�1�"�SO;۶��!���D�7�Cr�~~J.�7��7��ɦP��-�\ZC��`J��jl޴Q�3�Vl� �6fY�#>DyX���vA>Tzc���h��6�<k���8�f��X�ȭ���ŧ��+�A��/I�x/��f�|IL�u�����]��p	fJ�XG3��<������CZ��v�I�bHu�Ο�}�N�(	R^.$����{��s�D1u�Lq1�8���q�g�Z��k��Ce]j4h(+��wx��Gpͬ;d�]ꂙ>�,U{S3{�A�|���+�E8�	���{�/A{[f�]����S"�jN���U�GKB�{�9x�ŗT4w���.���т�.8CJ�1���aq;z�����w��f��/�G�褟M0�&�c�D����բ?�����F��T!��3N��o}$0�L���@gKY�tng��olZ�B,k��r��i�:���a��I8~�x����h��P5�P9ttt����B��m���:Z�NK�N����.AU�e8q�,��3�R�Q�_ʋ�X����ƎX��55��aayk�C���v��gb�_����ɚ���^�LO�g�|"��$Q�6T���q[S[������#����M[ŕ(Bbʢ9��/@wg���>�_�E^?��1$1�=�;�R��Wu�?_�H���jo�i'�k���UgeGCL;���"�WQ����O��]}zؙd�0��Չ�=
�GסG>k��:�=��^����&\k� tt����������j=��֝�'���sϖ0��#G*7�k֩�_(�5���e'n��*�{�eE�lv�	g(���7\/��@������AF�4�U��6HF<�>�M@�ć�|GqH��\Ɇ���LB&qer>���w#:qD���|�@u1��=>7̾6�s���0�����Um�ΦK������cFV�أCV�D_�ه������k@�y��=8yƱ�>�V M�xl�s�߼6	u�N��.<I�q>�\s��[�N�Ilv�^v��o�$-���U�[�`KC3��=x_\{���v�I����9�]���a��;�:q�m��/�Y�o�����XG2��*��7]�ɻW" +�ʬ��H ��&#����<�~�v�Yx��Wa8#� �f�}��P�b�J��Z|��
l��O���c&�Ŵp�:v�� �V���b�)cq��dN^�(�߯��u�dS�H��/�Csg�|�t���'(�*�Ϊ��D_#���${Q�/�?����_�!�1�8�����b��9������
)�YN�d�8�$x���������g�"[�?��.9��[G$�quA�}�Qrؖ�%�+�f��������b�\hq�����>�H;�8��������pƌC��'K�z�,1>>�'v��L�x�*�M¿Ͼ{J٭	����9�5?d�X�$�X�~����C'bݸ��3���P6l�d!�nhQz:�1�_��K/��P�%���1��74>�����Y'��/6���ٌWn^��]m�J�1���d��L��q���e�r{��Q�$=x�	[Y�3%������_��4$K���F����:��P:p�����W��.�(K
ל���1r�i��懱��sV��k*���mW�Ebz��}�L�t��p�Vk<��u�3e=�T�������T����!k��=7Z��ƾr�v��X�i�B�L�w]s��\��o�o~���K��y���+9��u�b4(�x�7��G�AD��+�q�>�P�N��*�wk��������}�l%��f�=xl		�u�p�E����p�Th�����1�!F3"N%��ϻTP�S�̙k\�z;���a���S:�0iT�V/D}Iq�ќ�q]pU���']��bΌD%zZ��z,Yr	>xc!��6q�8����+a�����C��x���mx���P�|C99�x�a�{��$r�ي���ψ��hB���w�&��.h�hjǡ��o�)��X��`��`���(.��N��I�^|/�l�d��=�I��(���:�Ν/^��В�p�	ǣ�~3\�b�~��Y���i��a�Xٿp�9g�8�B�ˋ1#��%�҄(��Gq��
:�~���X��.AK�>�l�������nT�0{�g�~:^y�#8�Nm��Jz��������+�Y9a����^�0m<�>l���
	�|rY5�/��*\>����$��ށP�<���f��>��=v�؄�R�M�8�ަ%.f�GM���}Ḏ�~��(+/��de��2�9s^��^�݂}���𫠁*m�N�Ώ0��o��&(��h���!���k���k1�߃�c&h��ɨ2��a����câ��E� $$r���_�G���gϒuϣ��O9X��ui^����n�!Y!��{1��v4�>3�T\Q�F���<���Y14L"'�9�!��1l������|�5�QY>�p��GJZ�p�}�qǭ׉Gk%�m�=��g���)�$�Kj��gK�qc��w!MR��z�pߜ�x~�\�Damm���ذ���v�﫮�Wrk����(%$i	��c<��e�T��94���G�iUU��Y��@Y�{#j��+145������ࣸ��a/h(���-�;�VV���Kq�C�(�5�ȹ�)Y+��1���L�2v�A�����K�cp9��9���b��J4tMg"��6�?��Cj����,A�v9�+׮�'jPF}�UΠ_~�(�xL����tؕJ:���6����ا�@�Dg�^�u�C0wέ0�u��-� ���!־��\6�y�w?_����R�v�yh�l&�~�)<��,�,�7ճ�|�H�;���G��N	_B������3�j�a��zL7�Xc�Aw}�f�?���/�+mv	lo@��Q�S��S��j�����-ln"�.ɉ�r�)�p:�)�6_�^qy���fa�U�+Vm�1G/�ա�TD>L>iÛ��A�_��k�/FqeH͹Ll�f��_\�O��ZP�m�)d��z��p.bW�ɺ�[Q>b�A� ���.���Ðe|�sO9mr٢nR�aC,'���Kk�٪e��.J�����~q��[�Ϙ(T��Q�[ s�c�,���T�<��N�$��Ub�o+����Āˡ��F-������~���'a�+��`uA�,�:�Ki�>�r���HK�L`Sr��VJִL��ʵ c��D���z쾠�{�xo������8�j��������O���pk����>ٟ�8��b���+�߿vSfq+ݙ dW*9_��߁�>�H�Q�V�XfL��c�aGK��Sv���=Z=2g��v�fı��j�L��H�%4���'kf���3D9Sʁ�����)�e�5jdEI	�ύ��~�$��4s=���������GCt\Y���a��|�¼��K�_���;iU�yKԩ7��������'�\���S��Ĭ�F���e��T�!=��Z*qA(���1,/��!:��z���S��w>���'܁e�&�`V�}�A #G�����-�E��� �҈�X!1��o�I�`�x3^TZiN+�"�r���w��������c:s˲�
�l�ֈ��x���Lֻ���n3���ۥ�3���K<�Y�:� ��C]	Wy�!��v9 ~�Y��ȍU���)oGJG9��9r�oo�A;YVZT�ٮ,��xR�����3�'X.��,��/�ӯ������I��(��s��b,
9��f�	�a?w%��em,�!&�J�2�˪��#�w�R��/�Qѡ����*�'��R{<،SVV�ܫ��A�C��ɋ�d#	{lJlU�'��X�a��*R}�D5y�r9��|���X�3�#����e�\v�Q��1@�ONnJ��4gt�"�)��%�>6���-�\���1���`��a��¼C/J͙1��9��5f^��V1�2��%�&c���D��P��4w�K6@;J-Z��ی�zI��n	����Uv�+�IU�`�MmF���K�!A��l��ay�J�'?K�Hq���/��T"��
oTؓ������%�
�N�]:]�J�ar˟���U���\���Y��ڦ�`¤ �ᾰv�z$6u�~fRV�3������Z.��t&GE<,�x	c*��>!��odyYS�s�f,�������ȣeFV�9�CgJ�yd)3(��_��B�^��d*�HH�Ͱ+R`�\R9�l�ul��ܠ\�.a�߳&�NR%FM��ď.	p<A9D�N��T��e9�/!��uP7�"BL�r#�-=�9bq��8�l����	�6� �5�e���t�F�z�z� ���]Jn��@Q�lu��Tv:���?i�?Y\nV��Gދ�L���Jo1g�&�;F{]X�e��hn32�6����R���%�"���<Z��咞���<�?ͦB�IV��(�h%�A	�(/
�_b�[����R0��u���%e�k�1z1�U��g�ܟ�7۽���z���}r>F���Լ(���WBw�#�6�^dU�xxj�X,M���Xŉ�"}(�Я��E�k�9,��RE� Q�.p�N�|���
W�	�9��,�Ҥ_�+P�~�9y.�K��Alo��/+��"!�����Ce������2g�*PZ�nKs��I���?V�H�W��I�I��`?FV����e�y|Q.��$�r��z0b�,X�ŵ:B�pV�X}p�Pb�n���]Xn�0YĬbp�_��/~Z�}�p�g�<b(P��8x����=#�ř���*�gK���Q���O� ���up��:m�ډ�O=Yũ\N�Z��p��!�bu��5ᤓg`�c�P��5k�/!}t0����&vG�E�I@$���4��٨4vᙔ%�\��9H����cGT�*S��X�~������j8L���<�^��j$���d5���E��I�k���*T������&U�f��Q���R	l�
�Į�T���ތ�����h>k^B�Tܪb�t3�_�p���lS��?V��G��*P�t�vx�N9���2t���'���s�������żp���,� �F�8h�$�5x�����cϊ!�������i�Dل��w��dCG���<���)�q�VT�ӵ>�K�w4= F��Ue��Т���R;/Mv��b��y�ޓ��oI�G���:��	�B����NF�+��ҁ.
	���!��_t�-|E�f�!R�23�T	"#��:��0�!�+��+ψ!ij؊�O<��ހ��	A���J|E(�
��j���o@˕l�2t~���Hc�ɣ�js� 7��y��2�F۪ә��u���ݷ��DVR%�wn�Y'���xG{�r>�2�ňt�ʟ	h�rL�~0�T�ərZ��%\K(^�1C�$��c�\������S�y��7�h:�j�e������c��y���4,��[UG��O�d��^w��IXΜ8H1�&e��kJ�W��#�0!�x���`���P�{��%b9��p�3PY^�ܼ��;TNT���,�Ry햶˹-������&1
	q�daoߺI��$�溷��?V	��D��%(��ǟ��3/��ѵx聛p�-����D�s��cO#!��kk�����P���|(�K�X�����m�&�Щ*ElJ����I�s�rN����Q\�3'z?��`Noo�΢�D$%�&��ˍ#��Q���?)0���m(oT-F�J�=ꠊ��	G$����ӰSQ���Ǎ�x{�<�>�j�Z�'rP6w.�0CH�]���A�<<|VA��4���	�b�xK��t���NC�O�C��/F��,<���d?��k��$6{M����I��hx,���Ǡ��M�+a9@4t��0�Ac���7��=v���9���/�߰E.lL�k9۳Ǟ�P[�Nq��-�q�H')�ǩ�Tʴ&�F��#�_U��t��3��?���x�HKM�W���nb�+�@���L?R)�N�q���'a�>��!��3�J��t�o�A)�O0��-[�N:�P�F�DskH�S^�B{K��Rv��j0�3>��k���x@��6mބ�&�E���M*^3�_Vo4:~�P�6��M����ۻ|�re��sxL;z�x졹8����0[q�a媭���p�J���#�<�SW��z,�u���DȤUS�;��Ξ��֝��3�f�m�c3^M�'��܍�Q	;�A�y��Z�e�����`��5�kʵA�ܓ�į+V�G�N�8�����@�8����h9�d̹/6��v�}xt�� ���+/DgS3�w��΁��Z�$̈�cP�̋��.��Gښe�َp�%�b��~Ep�IǊ�b�ʵȈ�:�kѼ�A�y<����eJ¢��9�[����q�'��u���c۩����bQE��ׯ���}w�Ͽ�&qu���:d���1�ц��G���W�V2��%���],��oL40���|ƚ�����#0�
3���b����'�w>�\�[�4H��q���p��'*��:k7l@�X�Z���k*P�K���x�o��	��Y�^�j���}��S��-/B� ��;4>a��Q,b[C=��~_���X�4t�6d��3�����8`�h8=6��A�`�:�DS�
�8y���[XCU��9q1ci��-[�c��ۆ���Q�ֶf1��\�Z���,��{�~��/���9�(~GG?��g�r,zv" ���C��d//:��ڻeÜ�a��ݺS���Cp���/�s�������N�x.\s��J�F���׏���,-E{g?��q�x�PavA.��-;[���C�K=��s��sUA��0bu���ܲ.P��M�z��� ^��s�4�d{����8��:�tw���(&)�Z�ʯ�[�v���k�d�9��J<��G����ݲ�'M�a∘(T�Ge���G�8��l�3�Q�dսt�-h��~��bh(�9qo	%�m��,$%!�rAA�?�ه���K[��T���G��O<���[0����w�VSb��E=�,�B�y�xJ��X��e�X%|���U8h���l�(��o��P4e�0�=�����Ș��9�'��p!e��9O㦙�}�_�B�s����T��8/���{�l�a��d�e�v�����9x����3���<m�:�M�*m$I���!1�AP��9����%��"ω�N��nA'~�j������?���?�����N<V<M�R��۱e��5�1�?� %��[�3$�Bİe�m�9lځb(����ŋ����B�KӬ�_����͠1�1�������Eo⸣�PR� V�ݜLr���n8>��k�sz��_�0%I����7b��k�l�Pj�����ukQ!��)����K�`��~9�v�}�Y
��VnX�	vC�j�^z�a����S���rǝ(����!�l4U1���7�(RaՉ�>V�C���Z�60 ���o�v"��B�1��-���$�X����o�`�5 ��+ތIƾ� bAzk��(-)Չ[�38��#��˯��sNW���5��0��e��ra��������ߘ��\M�G��j5�r9���lk���Y��v��xB!<:�ie�%[�-yMvT��x��q�駠��Ҝ�u�`�qc��V5�ϿlHn�����	y�7)��~�]�~��شm�" �����I!J#2���%�}ʱY�7��11�-��e+p�qG���O'���A<�p�������?�g�j[:s���
�o��&�s�M���~d����̘�ufq�]sP\;\�殌�����/��òe�^)�p�	I��r�\�#�����`���J�&u��oB¡�,xw�r��E	�p�v��_6�*�5Q�3�o`L�2<d��/�9��ٸ����^S�(!#��YB�y��X�b�!ё�)�����;��K��7?�ۈf���A�$D�&Vc��_tP�J��ޮT�~BG�V噰�a|H�o�ȑ:��̰�` �ˍ��w(YJ�jZ�Ƥ:%�-��+o.�k��}���@D�yz�8{\^|�շ����t^����gjk��/��#I-�1�e��'x� ҊU�U6�*�	[j��0��'1�o��)a�O�OL�ڝ,�%�}�}�݃1�U_��C��JYQY���Mk1R&ռ�:_�&���ȪI�w��,XZ��>�G~(L�11��>Z���xK��CuX�lhw�1��|>c�z��yω���k��I�i2lG[�v�pW<�Kj��t"�.^(�}��1�0�fx)�ty�"==x��O�-*Q��):�]�Ո��	l�s�x$;j����w�$b��o��L��兴��F��lL/+
\_^��>��y$6�o�x8��E�)3�y�-�tn%���kN�L�@V��&����K���hC��O<-x;�zz�~k|�=��f"��\K:�>ge/6�h��/��c���ϣm�6�C0�e�N��B�'8UtK<5��$6f{>�
�>�8j��8���a��p��@%�FH����I;r��u:�[H�.��ذ}�B��G�)s
�qG3��`Ę����(̍� FM3萐�<,\1Ks`Ѱ�Q'6�ȡ��F�8t���&�hP��	e&��'y��Ex�g$�j6[��� drƐ$���=c
�q/y�=�bt��0�����,��C{N�|���g*ݥ��&H����ەC�H�8v���(�2�^'��X���W��Vs�/C^�O����U/@��~��{�."Γ���8�?�4lC�9I��P	��l��㑸�m���e6����{��_�\��+~/Lf�2�gt$�H��قX���8��7��i�=�I���Nmɲ������\0��[T##{4���Ҧ��*us��]T�%?�*4^%�fl�j�9�KOb��+���pc^��mr!�{�(^�U�T:��<�dۢ�gٛ��g-LCU��%wxC�h��X�����pr����|����9vMW�]ʙAvlA�Wo��A�ڂ|��閃���$��T*%�Ʌr�j�}*9񮄢���3ې�i�6�9��#$c)7���f���)1�d+����[��Ԯ�0�B�/Ɩ�qNs��U��{4��X�Ó���H.�Y66���v���M'jM:ʟQ6��=I��p�+�G�k�����u��}n+�je=hdȖ�^��8>)��:�ъRo�_.qN����Hs�^BV�l6�?hc�f���&�y���h�ѿN0�lNm�$M���N��g���ȯQ�=$�C�Cg��,pl��!�k�[,�Z���z���ȳaQ��3��������e���۩�!��Y\���x�{!_ �Q^q�U�<��]�yJ䌵�h8��yع�(��6&���{�W:�m�+z镸1!�#�W�$fz-ʹ���#�%C�J�ʎ;~��dm������o� ������#�$R�u�ZS�rC9-x���$�$C�]<0l(�p,���1DA���v��9^墀&7uwL�M�~���(��;t8�C��PG��^�ٚطQ8dZ_�$������A~��$��F47��IE�v�Kwq�����Ť�cπ�d�z��%Ƽ��a�qy�x�P�nL�>D/-��\Z ���F�utb,�]�=��/4#�	��j+f9G bׯ������+j*E!�|N�ML��g�ȕ�r�ԛZ4E�̦$�xHh��Yo�ʕ����F����19��G�~��t����D���J��\��}M� ����QA�n�MPv�g͜�?˳�`U/m��X���.`��1���w۴g��a���JU���U9휶�ty}��ֳM�0�39t,�A�����(�Y�kڐڵy��[��qSS\^�>�hXu�篪��ĳU/a�@�@ߴ፬ּ���$�dS&��Ŭ�F��s�!��Qi�])08-�]��}w�����3;��l��]����?{� �&�����%�-�7���c����  ���;�;;��wf~�9ﬂ��u��gX����~��<�|�y�����ʬεa�F����V9͡a~mR#a�ǒ�4Q�䐵V���I!PZ��T�Ԁq�e���<Y�@�b\��K����Ez�cIk����АM�8�����'c��w����_��F��%���Z�Eڞ�h���`����N���rj��/,sH4�WteҚ���-�c�!��1�D�WԨ�5�e��$��J	��ߣ�!�!�6��� �UQHiS�1�b�iP�FBC�!���7˨A
CPɫ��Q�����[����অ.2�����9� R��J��F���H�W��GA��Ԕ��J"X��
)���5C#ٱg�"*q��煲S�ȰK�u���r%]���"՘B�����hE(SN\1d���V�J�85����
1�x�!��'�|��Q^Z�H0��9��ke����ވ2J��8�ln��\���>~��Z��I���)���c�wk0��!݅��/��h�
%�����^4�3�!ˀ�4	_�a�_^��摊�$ǖJ'~ȫ�b��6,~�I�Jk�{9JK�d*e�YW1�)�&���-2�<�1�P�:-~/VIY�L����U�Q-��Rd��u:;�X�2KE�p/����b
R���	�,2�����..�-/�D��Z�e�9��"�d0V侃��Ҋmo�6YM
	-Ũ���x�d��g/!u(itt�j<h���*K�4�Z;��VU*�0*�A5�aƐ�4PH\�{�j|\Rl)hO���2%{�0r�9#�8/� ÷����:�0 c�i�To�R����4������C�9���.�������_���J-pz������.�Ȕ�3�9# fE3���ؠ3v�ePo..D:!��Ù����z��&�� dԈFL3F���b��O�}�[v���ة�g�%�����9T�������:^�$�iWk+�����k�]��Cf�dp �4C����~���j�B�S��4������IftO�i>�pJH>�]m����0����u0�)r��`����/��zX��J=���ҹ-���zѹg��ѕ����g="_0�j̞y#�%Q��`�thug�1c�4L�|R� �>��
�,f^r�}�%,��;x��9�?�w�B]䇴�������2d��1��#ڼ��ޅ��|W^v��Ŕ/��r�K�|�oѢG	�kq�8�t�N͝����_¬�.����rL�0^������9��6��۴�,�]ӄ|�H2Z�/FF�����N��<
��1G�̜����[ SX��٭�̜�82J�$Yx���pΟ~&ꪴl?��܏`8��>��[{��ߜK@*�]�:
Mq���_|>C�A�+���խ�βQq�>�|%��!IF>@`_V ��{�q��	��*ҊQ�ruPS��c�%�W�=GX�Y�B�Pq�	�.9���\x��ڀ�/)E"BII	�3��֗���K�i@����tK�٪)�ݍ+ϟ�ۡ��wsKqP0��/�O�	!����욯�XS`h���c��Q��=ϡ��ߋ'��үVj���;JӡP�I���\R���a��(�Ϗ��4�W�\^�1�t��z<��ex��,4���eh��"�됟��%睭��k�+	M*��{�1��c�|�|��&��E�٬FQxO����W\v�;�"���ڴ8��Y�G���m�܏��J��I� M�u���b��M�oW�$�����5C��=�H�Ge�_��`I�Ra��}j��">m�����!_�)�Ϳ	���Jkky�f�Va����@��z"�j�C��V}�x:�V�S����x��;���'�E��t�� M�EN.�z
?�����Oq��`H�{��'�_R���_����P��̝��㞛.G��r��hAؓn�cAԕ�;�ă���[�fD�H�%
�2���m�sO�^�̥c�#
�AXK�ŉڑ��Ɵ�|7,SϚ�8�|P˪�Z�,�B��X|^,_��^ç�u�K�E��p��t��ůn��{<@��c��=:Y^��(�M7\����=J��?��e�)�T�X�ι�@cƸZ[������v�#����k7mך ��ƨHa�J�Hī.�H��B�8�f �ݽp�h�Hǽ۷㲙3��ko��J)��2v�VQ��|�!(-)�i�YGC��5D��V�s�9\�"�����Tg1_��\ c�i�&s�%+)C�S��ĈL��<�|کx��%((�2l��C��D"Ҍ�������=5j��܎�ؠf�M>���m�<�lLj��X.���O=���f*Z��]H#Y��0��-j�.<gz�	���%ڷ!���_f��Q�Ŵs��@����AE]�Ӭ#	C��(Z�������7��|�lV�54J2�4g1c��u:��+%Ӆذej�ׁ0>��'�e����@��������.��;֡�����غk/�'Ch^�V^COh�3w��w��s|�yJ�ػw��:-:���i�R��s�:��L�߻�݈yw��^։��5I���}���S�(������7�x=�4��8v�1�Qƣ�<x׭X��#pWV��r���ݸx��p��њwȳ���?�{�����}�5W`�(�����n,�}���I�[�:�:0��+P)�|���z�z|�d)eَY�OC�^e�.(؛��_���!���Zq�ݷ��ā�͋�n��r"�Nj��s:.�l�6���z��.,X�[��|���ֺ�>�g�uE-�\p7��v�NS
��ê�̢�1��E�������ب��ɬ.����.�l�Qk���HI�c�)��x{`!fZ;[���عa���å��#�֊��/����R��A ���u7���Rt��VA�ISݽ�4\6Z;�*�$��ʰ}�V�"Ŀ
J�)D�zp��b��8��hv�Z�}�X��ࠗp9���?u2�{�5��ZiP�NG����5�U�R�\�+�Y���bL�r*,D#���ꗳ��ҥ���|��^�8���.E�����K�����_ժ��&M����ظ~5�63.��T����0]��{�}\z��ыĬ@�}����S�P]Y��x�7��!�;��_x
J��g�K$��ig)����;0n≘7�N��n/�P_W��7߀��6bDM=�����w��)9��؎c'�S��گ^�Ͽ�;H��_d��;�q2�)�����=�� �D$�"7׀��������X���x�_�V��QU���__�A�哏�5�7oS�[�Ō�}�q㕳�����������n�v�DR��xuѓX��k�]���v̙w;ʪj5� J{t᭚`�8��g�b��@ "���<�@W�3�����PV���ɦ��L:b�*���]�-(�,��E���x����=���(
�.#�Z��2W�LƎ�ĸQ�Tv��9��%����̙^���ᕋ�ڊ��^����u#PL]�T���U:��hx3fθ�����I��_?��y���/����d6?�� ���9�`%z��_+�ȟ^ցH��(O�;�|�.�s��	Dc~�

4�9�.�β-�o��>��[��ZuƬ���u���s��T�wA9�z�O����[�8�6�$��k�@���2�dD.e�����&g��w���{]��T���B�w�YQ[LC���s�╿�3Y��e�{���q!K�}w;�x|>���˼�K/�'=�$�.�}>�x��J�XW��~�����7�7��Q�Gy(�Y��-�;��&lY�5Úhm��/Wj�Jx�4PG�q"RѠN���{���ta��V|���}�T�=t$��<��Ǔ�t��^�=b��WRH�n�N<���r3�D�^|����ϚF��COg���ֶN�T���aTvSr ���E�2̸d.�>�Z6����o���.�-�7b��s0��ߣ��Fs@r��X]���'LY��UT_u�΂�dx4�{�`Ε�����JJ��赒DI���5��\����߬^{��C��������p��E��ru�q����5�f4QYUFTB�X\x�������Z�.R�8��'�����vt`,�u3�F��c:�"�n��r#���ү����Ұ
5�G���H�^y=�~�n�vt����J��%���^�N�(�?�y5�|�p�J�������5�z�n��<�oŔ3Nǲ�(�AW[;θ�BD�w�����P�X�!��f��K_,����G��t�z�1rx��)1���c��:�X	8�N�<�ȵR��$�#	K��1�B<��B��h�	H!V��0�C�:m�$��λÐ��]�"��8J�kpٕ����_F*�K,�b�ϐ#IMœ�`��l��Χp����!;����1���e��N��haW��M�,a��c���i"��Q�����zڦ�f��������7�QTc�_~��e�h&EMv3n<v��7�����i���T��hւO�\�HB��C�^[����7�B�=�C3������o~>܅eX�؃���(�w{��ϼ�*��d�Nϖx�z��ު��~:��cPZX/�?_e�N�$"�g�p����'�#����B�����8�DUV��o��7x�D rl�,�VX=��`�2�5�`��FlܶM��")��cȽTV��?ԇ������&��9�s���+�o�n��M�ZgQZR�����0�72]����,U~�X�"a��\xb�sx`�uHh+'Q�/jbIo@l����j��&Ɍ�XE�9�z?^��N>Q:���"m���ak��3g�Qza7���
����F��	9�"���Gc��3����u���v�l��2*��k4����8�lل
��d�����&�gh�|�VȜ�cS�ո}%x�W���{��M�^��^�������b))�
D�z,��/!��ϼ���j%e�H;�$�]��/p����_t����������yl�qA�e_�)|��4�o�#Lh�%r&�d�����FB���ە��NI�A)>Pn�>�5�q�����t"]J[��@�z��M��42Ke��.!Ҍ��,?�)�4�ĳ����m���MdLϥ���rh���BZ
.-�ťVĢ}���������2�����Ñ%QB������D�{�
�+�B��y�		�S�C^;zc2F���E��	���W�}�2�aɲ8d�t$��1\��$�H�.ZfiW߲v+��k�&�xGj*��G�-��<��F�$�L��)񬿬{�`<~.�~8ڣ1���m�|��v��q����fS�d�� 9�к)�IB(YL�󗤭)mAk 3�G��z��f0�$4z��En
�A[W|�rD�0fe,���JԜ���;��P���dF_�,�D���tz�FDe�5��<	ޏ���+�⨱MjH�yܔ��5&o���Z���MZ�rXt�xذX�a+jJ���5w8�z�&�RR.\�w;�����D��/0�H,:2��)3,��Xj" ���:X'N�(]�k�m@	�2�gWB���Xt̾�n�ne��I����Y�Z�����a蓹CI;n�A��o9�K{GJ�e�q�a��0�΋i����.�Z�/�g(+�!���O�~_G���ZL��ƌR9����f��:=�a<�?3i�JȜ%����R�1DJo(C�dv�Ms��}��hUg���F:�uMi���ϋ��!\�=��J��g�$]���wӓ����ý4��2��Ak
|:--�i��%Ǻ�J�;i�ǩ!��i�h,q�t�*�
qut��Ce�@�b�����Pݳ9�t։�J.����	��p��6즞�)��9��N��ʘP>�Ǚ�0�%�]�R�p	�E��X��rqa�*�A�/�C+^U_��K���ԫ �i�21JN"*�����g��Th
�����$�l�b#Q�&o�Qh��j��L8�y]�*�v�&��8����9��ɇ�fXz;��%&��$���}Kܴ��N%[�dyQ�~~tP�T�(utn9y�~�T�(�UN.!�0?ː#�Nt̩�
��\)^���KQ�a��)�
8K*��wk7��'�.^6͉�ɩ�6e~�*�0!��ϘrC��^��l�A+)�gi�̰E���8�L���6��XD��\Z
?�����{��	���WT�!2�䰙�m�"��4��n��š�sF��w��X;ﯤ��I�#�TQ���"�H�����=��m3����Bb��n�5�d����K����� =m�_K
}p��.�Q%��&:�H�G����R/!�������,	��=������tʐh:Q�+�(�p]m��ԡ��[��Pɽ���9ڗ�ݼ$N;�d=Ζ�<��.^{JɆ���{2��i=��L��%Jm�*�t�#�1J) �O9$��OA�R�1���/"��B������m����c�Z�P���aѰ=�Q&�ؾk7u%��`�H�}����u��v	�;v`D����`.,�u�:*��H��:����c�b�::_�E����;�PuR�n�:}��˄=i��dS:'��'`��/@�0��"�r~Vn,)W�I���H��x^8i�o�@Ǟx(`m}$�9n�l�a�Ç�� ��걫�G�OQ��?�{,��{	����Sk��=-FZ�lB�����c_�ι�S

�z�Dj����ݣs@�Zw!e1���V��Q��A�.�î��m14yi��(�Xa�
y��7��ʘ��V^i�T>���0c�ʒ*�Ǩ,�qH��`5����Dz~T)���&�h ��]���c����{{�0��`��f�̽3��u~��� ��%��1�)�X�M�6I�d�a>apr�P�=F�ZZ������ܨ����l"�)aWOn�qh3S ]�1�6�V�Y�-*/�#G6�����>x��*%��0Q"*�����[o��,Ё�y�|:�8�b��.Rta��b�=�Qp$!�NW駡0��ދc���-��~�"t�|;<�ǥ����K/":��c���B���c��:lf��V:A����=d4ٛ��|��� ��E�i.&4��8�:��ڎ8�?*�P��P�<В�Tr�����|�)�qa��ߏ(u�"��U��PB�"B�J`ֹS�\��� I���,Y)է�^�z3&�q<�Zp�����?U�k�UN ؉�s�E��-p�k�_�1�N�D�:x��E`�V,�n~��?��K�چ�"98����S�(:ϗ���ڔ�F¶,�Gu�m�F��r�M3p�ܵS�X2�0Snlyq�~�mJ���"|��F���X�٤�.�Ś���0"���B]��w_��Jmaxr�ԟ�	�h�|��e����Mʏ�6�J"e�`���+�����b��ס��M��V�h���"�~"�*\Z��=����&���-�6�j���_y6�8K�XW��C8(�#ޛ�p"�G������@��O�g����ϸ���Ҙ�A���W�T�V��J5]0�<Ҍ��أ�aU����0���UAD�j$Ċ9��I�U4~�]pñ/QT_�ػ�'��I��5?m%T����"�6:���_$�`�8
�ؕ�A�J"�^
j��D���q�'Ӫ�U��j�2�׹�+h�c{�D1�Qr�x|��s��M�k{�N#�>��"��Fq��OB��M<h�;�L�hL��q�-jc��N	��b_E=b6*WA���.��G��?�i\�ۑ�����e���^���t�D��9
��~V?�݋@�=����'}D�u����sеjR�-���a�i�Ɨf?b�Bl�ъP�I����S*t}�x|��ۨ){e�VE��G���E2�Fsiģ%�=}l�4�ĐE牸B��ǡ��B/
O�c%�[LȜ�����ga-��ְ1��s�V�:l����|<�����2lh��Is���|��5�BX�#�ш5v�0�!WY#�m1R\�	�jܭ�pO�2��?�1�h�!:�2i�������b���M�C�v�jN��e�4�M|N�� >�h	C�rD�&�Q��Q�N�[��g07�����K�Tq���M�:�j|�9��n{=]��S�8�V�/載W�um�|����:|K
2��Y��?+0���R&3#���y*bDVB..�o_J�ua�{Kay����S��E�~�����>���#�xsߔ��[�� ��8���K~���=��i4�������kT
"�=r?h��wo��������K.�7���M>�������8y�ׇ'��?��O���	���K_0J6�����GH�jvҙ0��������u���g��.���G6jP5��iT�p�����k_�$�<��{ܿ��/�~D�I��g��Ds_r������0��_�g?����곡k'�@i��Ce%�{�����7�l���I��o�+����SO���[���ԟl��}N �s�z��{��C�=�3����$Ŷ}��<��4$���?��~ߑ�*r'�4��{_������m�:t@ׅ<*F��3-�ǯ�܆�qK�$����}M��B��B�z0r�r�7���z��`�f�)�A� =dͥW@�JA��|j�u�5��jY����O9��5?��ϐ5�	����������pXe����!�(k.�<�v�:��jW�u9��f�)((0�����E�Ņ�6H�    IEND�B`�PK
     eO�Z��I2\k  \k  /   images/35c60fd9-1fb3-48b8-b3d7-7968b0279531.png�PNG

   IHDR   d   ^   ���   gAMA  ���a   	pHYs  �  ��o�d  j�IDATx�4�gt��q%x�!a�{ｭB(o���ڳ�dS�(q82�Jgݏ=3s��3���h�E3�'ۻ�e���{�H`nz�S,0����ｈ�F�{e��pd1��ｃ��v�y���?��L����h����@rL~��ط7��ߺ���5�..�t~&�郯0����_�#��60�k%���N9Ʀp��)�z8��}�^(�O?��%~���g����x�r�僻�\���Y�KK�'O*����yـ��~d���օ|��^?W��W�{p�)qx��9��r\>}����֍��0|��e��v9JrR0����O�!��?��������_^��z��`O�/�{�7����n�ɇ��l=�_�m�L�ceu	�K����8ğ�{&��Z:p���w��[��n������g�x��y�����5�v�y�����?�=��|���"'&f��'\�̀�vl��#���������;p��� }���	�����#3˰�wNVgxy��a������q ����
]���'g�a2���{��zW~~�8�?&�	�1a��t �ח�>�����?� X�Vi0�����?��3B�C14����0lno����l#+=k���M�ᔙ����GxX <||'�;�XZZA���H_�\\y�,�,#1!ɉ)�y9! ��]��ݱ�l�
���GG�����[�0L8q� Ss3��IGKs����l���+�04>�����s<;��uo�zU�C8��w�y^V'�� �ַ��iUF#0�����e�������W`q�`av
�c�pp�ں���k�e�þ�E�h�"�x��YL--����M���Է��3Nc�~ 7�O��`�;��%E8[����<�i��l�W����|�g���ǳ�F�Ǆ��V�++Ɖ�T9��U5p9�yΝ��޸���Fym�.ncw.��o��6fO*����@k�0�=<�o���X��6̭�������7^-�'���cs�M�Ђ���\Ԯ�4u���g<,��e�`uK�'������~��7/�$3#�#x��Fl���wo^���ct|
�N�!guqcC-�Gxʇyy��W��o�x^���(�ӄ%��ȤV�24���E~n���6��,Z��(��a�8���G����JϚ���ܜ������},3f�������ױE˲X��k[�]^	�	ۻv��}���I�y�����]�tǳ}p�;�k`�d�pRa2�ڏq�Y�8�z�!'���D�:�C.���G��/n��ʛ{G�58�#�w�� N��`D��,�6}ψ]B�!�Hc�<��9��L����V8�93����_|�ق}"��j�Ǵ�����ǜ#�]�C|����oo�Ǝ��pv2"<�_ރ�Ox�D� �-F����:�|�'�3����`M��?���^c�7z_�?������Y&�7x��a�1l��z_���A~�02fm��pD|e�!Bx�`_w,�n�b��p��� 6"3��蟜���@؊�Ch�/��7�=<�*���X����z�������(Z�j{�hX{z� ��(5^祥oӄ7>�>6��̀����u�r��n��6\;�WwZ�9�=C�\��bQ.�9C��i����iL�\+�dx|� ���� <�lT+�ɠ(3$��8d�8S��	s���N��g�U��%9�p�����"-6���D�8���� _����\��6�,�!;))��XY[GBD^zfV6Q����d���">/5m=��A:'� #�3���pZ�M�����D,��"�A����=���ق��#36���'|v$c������C`��<=���D���&tyy⍳����3��N��?��1B	���S$���{x�b)zF��g���'`|�ɹE�y�K������b��;�G���,sNzf�q�0��Ղ��[�0,����K������s�\�ￆ�`});]���p�֟}�&-��|�;��~[���o^��7(�|����|��o�qq��d0�
	����kdP��aX�R�#��5�����0+���"."�L�	Z����H�A���B��i�Qx��)Z�0�bQ^ׁ����8�u���ǐ�O���Em-
ӓ��/�YCb�<{����� ��{7�M�M�
���,����|W�ǿ�cxy���:2��������pQF�]���M2��8<4!<��a�س�ӌ����
���čƅ�`l3�?���,�Ŭ�4%ɿ��[[4z������~�,���d	;����l����ܽ�އ���3la�xm����i=&�y�+fJ��h��9�`vU�#�&�L��ǵ� ����1H��	G&�221��`dl����gW/��{j��x!c5:�0�z�B�g�3Z�h<�'7O?�|���!k����x_W��җ�p���u�B��i��H%�ŝ	O7+��\�M��M���ALR*���z�ˆv��0�ғRRӰ���H2���A�5Y�Յ�+ˋ��L�����6�L(#1c@��I���7.1(Z0��L�����&.2��e���\���Y��#lp��{�"a~�N��Z��A��7_��m +�XES���^�7.�&z�𬮁񊟏��K�8I��U��^t���֕2��"�W5��`�@=q�(�q𳹠������;�p�D>2Rb�+<Q�آ����3?;A^n���u���������/wW<�����.��q=(���U��yO���V����g�W߽E�?���5�<�4���n���xg��44Ɵ�v|��3��.Σ�c�y��˗x�|)���$,�*�9&<���s%�T�L�Y��g��nwH����I,���:uM	��dI&#�����d!BDG�--��\@j;�7�Ť�Yݠv�>�hǄPf�ܾ�z����54��Jnn&e�&��z3������E�v�h�gg&w�=����:��$�p������il��Xe v!���s���nr���.cՆz�>��ыZ�E�Āx���/^�r�<8GX�\��I����͝�8&+�3���Z����0A��aeN�#4�a��C�0E���{s��/y_Qgf>ׅ�0���_|x�������{t'��I�fHS���C�*�s��V �p���Ͳ@\��E��$xG������	k���ǚRq��p���� �F���������{��g��M�f^g������H����Kټl0l�Bc8����y��Л�`�6sA6	e|*�̓КE�E�� k�&����������0g'���fC&I�����,�j�و*��i$>F4��e}O>�\a&��<���3�kLp��?�Gc����4;:��f�Q\�6�y�b~e�k%p�����<�k�*�q6/�P�7�$�|N|�?�G)!&,�O�����G�0ۻ��d�"�q�K�8Ľ�F��id8��T�q�T5RSl#):��S�C�-���Ay�^�Ġ[���{nҢ��[�YIJz23��h�ޞ�i����"CB���'g�N�G+����p���GF9��y������N�cnv�!��f\xTߎ@/w\-����2�|�QV�O	%�V^�T�I�#3����q5E��](��۾�������,a��ST�;�'\�:_;�u����	�*�y��"ѓ��k'A)�QX(.�p�l��w?� �>�>�Q��JgW�?��
δ��S��ē������vw���W��ΡaĄ��g>��_�wn�CFt0^4��%�?}�.�÷Hs�Q��ɿc��M��	�M���rvRAMs/��\.��O&�V��a�TV"ic6Y�
�7�q�-5!��)D��4-=��ۈ����&�~��94�G�	u��ן�%����_� oW��=zFɲ>}�.���B�e�7�L/����"�������\[!�������A����hd��{B8�����.�����	���������~G]�NRrDz��&�zw77���ocg�A~�i�i�.�͕6u@(���K��q��'�a��3`��P#X1���y�Y�&�6S�7�O�X���?���
�"X�[Z��s��ye� �| �
]��-�c��}��<��P�Aؓ���D�Gs$lP�vP�X����D�$ɧ�+ܽ����� �MD�+� �Ãɦ<>�m�^ApY'�)��¶��!��9�IʜHO�0x��GG�އ���r�s�\�6�ɂ
{� �����9�:[������YD�}-�,Mx=����,k��Y0���E2&gl>fW���}�
�T�ί�[����Go�#Ut��n`0��",�l�Wϓn��͉\���k���"޹q��}	����n��"��A����Q\@��C8!;����?�Kt���4ą����L��&[;A�Gk��2�o�Pz[˿KOf#:2���L�Х���Ջ�%��H��/�����38�3���o߄߹�����dY����u.�z�F1K<���w@����>��(�%��q2��&�R�12¸ӏ��C�Ե�/�}�����<�������w��0f2xo��O��=�ƛ�^��L�Ih��++]q`hjF�(Z�qe+�����v�%�i&��@bh�ZxsG/ֶ�8�N���E��0��47��%��ه��UX��磣X"m�Tk�0����V�v�a�lǙ�qplN=��ᅚ��Iq�P狉��p�5=����f�m|a��}W:�Q�d5��ܿ|\I��ß�����]f��#�>�����D�����q��rb\�B0ɲ�%q�e|I����Y�x�仞шڹ�|}��
QĢ��@���%I���\���<�'gVu^Vy�C�2Α�9��Rz�`e��t~m]��}�l��γMW���uZ9Ap���A��'I豳u�GX���?�;�̂q_�%N���_��¤��	�mr��,��@c����B�����F���߁C3�vek� ��I-s��@���4	��k�S��>W���1J"�.C2+$�&�'�戋��cV�F�����I��E�(��W�zaA�Jww��k|?~��11�$__o���3Я��W�rzr<����G106� ~�""Bh��EtG``r�����'�#:8H�sln	/�:scÐ���yeu�鞢�S��Q@���ϸ���)������T����M]Z��
�Enz��D|�l��,TL`0N�&����/'�̯o ��%y�J]Rk8Ή�u�Zw\>��E���;h������^�X̅7b�L�cx\S*>�V�.�T5�̀�;<���~x�:��A�S��<\�J�����:ɀg��.�2c#q�#�x��I��\��kg��J�߸r������n�Çw�)���(���)�<_�G�h���+��2���9����g	�ǻ��%?��|Up@���G��V�}�1!^T��T����O�G�>�yrL��mvR,n�ע�oQi�D����%����%Fgx�ӚT���Ǆ��{/115��_9�L����4ꀗ��x�ء����$|���l-݃��I�j�S9���C^zZ&q���i�J�y��_�ٿ~zၾ��+��K���M���Z�'��E�ޓ�06���|t��u��k���p'�Z\����aˊ��*��IR�ļ����H����".2�3�L3����[�!��n!/9˫�!�����sSx��Y��gk,M�O����O06>�Yb���!6�fH�65׿F�YcpY������hafZ��ؼK�4:��2�1�'����ʁaz���&f�L֡r������m����u�������.ۑ�P�_���r��V�E�3OL�K�H��=�a ��U��R�ϯ���I�����5PD.��q�j�v�
I��ưZmʰ̪�%gg�����`?�[�L|�C���������vS]=m�����jusr~M�@rh��8�o�f��uܱ�;�u%_O/�39HLv����������E���,�X�\WR�o�c+�n.�X�!��k(�.�TF�

7;'kze��3��@R�5u��yoo^)� ��n����$����t�*����Ֆ =}	��� �����,'=��^�N�����kl�A!!1��%:��{H�3B�r";�W���::5�	Ԟ�a���F==,����a�0~t�{N��{7��I(����O��C2NW'#f��15���0?���y���DvIX���"c�!	��[e4T������q;����42Qg|p�BsEm-a�,�O%��`�p:"����&������jvb�~�}̦��u*t<��n�V�T6Q�ڍ�xɈ�et�Pc��pQ���O<v#FW7Ma|~E�H��b���6WԌ3�i���Dlq�n��k�Soq��OS�l6��u�1h�V�� ;A!��Ԅ@oo���c�
ܕ�f���IM3_�E��$.��X�a<��Ch` U=�ynUk>�v���zmj�4��D�H��c�(|aVc�~!&��}PQ�@���֗V7�yR%������3M7c��G� y�ƞa1�	�8����l%����"��;ֶ6`���;���Rd���mR��R񊸳s��F_W	��共�mHYT�<��Eb!�;j���*%� /)�K�h�]��X�#M�O/p���r�ɠB�B�@�&Y���L��vee�� ��P�����v�h�P��H���a�qd��RS�z�2R�<�-FI����J�P��V.��\�$88N�9B��������36��`s�hI�5:Q �hQ��6T�J..���T��4�j3�(����;��,����#:)��U�fǇ#5&J��C�ɒ;��I\��Q�N���&��}����!75A��'�ec�� B�=��+Z�9Y�Ă@�DU��̫h��K"�EY��u�k��4�%�.ϕv��������,��^��d�*H���=k���urD���L�w|6Z��L��>�Wa˅�y���ك���l�,��Y��yp���,�PA�'��˧r�����$�����g�Zm����+(+��������X��А,,.�LQ&�����d!+5�דe��߫��7���u2�rU���/ӝ-x��i,.�&�N����:u�w���B�=2��xR�̟'��ǅ����Ih�D#E��3��N�%����b[�(�{�'rP����9d$��K��IW�V�Zg&ģ�񡪹�s��A�45ۈܴd��%��4�0%��$	�<�EbT8I�.>�{14��/�PtN"6"����W��7���b�#12S��?|����2\%|
c���	��?�BY�7�j^O����� ��߹�82���i��E����i�{d_�!'%�um\���=�}|��(�BL�K�����!L~��30wpB����YK�r�vb�6g7at�h�������54���uZ�<=]�&��ͧV���0�E���u�Mi������q�C�3�͍��/nh:):\�Xz'!k�1KTxNZ�B���F�m0X���`��,�[���.&	Y�����T�����b���HO�3Y	�Ԇ�=��_��yx�A8��hU�Ѣ���I�d"��'�wB�7��@Qir�nAXgBOlB'x^���)5X]����m�ۡ�>d������D��OR4��\V�������F�����k�M2K/�^#Eն��p��)b�"R���{��։��(v�O�V�g�oPpI.*5&c�s�v��K�S��E#9< =C#���38A���RƑTL�I� ˺T���i�'��P�089M�LB �nrt�ΘB�0�'��Z���f��+�ı�Ee�[��"��+|�����©���J�E�0:I���*�}vz<~D�!8�k���-Mw����o^���L��a̝�r�����k�\��K��>cl� �}�{db�$�yD�oGk{;��Fv)��H{S��5�Զ�k���[��J؉V����S����D��AX�C�VmS7&8�V'Զ�"�4ؗn���G�]Tk,�%	��
b�N�q���:|������e�-���a���G]�M�9�	�܏iZ�$�%k#|J�t�ZhG���h���4Y��kml�EM���9�C3��=��%[���[4>JP�����Ć���M�9G��>�hBRT�4���)ؿ�?��E<!��"1gFY���S2���92K7�E�8�����V��i�ՒN�]^��Nh%���!���.����YYQo(~������n�z�CrvuV��&d�v��V�Oa&�`����5m����|�����J	���KJ��!����dVB� �@Ƒ�z8E\�]Z�f8)��f�B�Y�.�x�d�i0��u
YY2�Y�WH���+$ǌI,\�S(�����Pi��Ci�[���U����"ܦ�����KV�I�[$�O��^�����Ѿc�"֮�T2����2���H�u\���,$�m~��\:��RBue�Q!�ڞ)�M�=u"�h!�~��q��]�*V�BZ|�`Z���-�KF��EX���+YD�������{�"�S���G��`VM[���_*H����3����vj�]x���$;�J�J�._�5�Jޕ�����U�T#hq	�f+�e�dKlu� ��2��B(�����EJ��QWOf""П�aD[���{5R�)Hg���@�ZX^A%I��ޒ�d��s��N�إ�,'��4MY�:Y�gO��Wq&;i�I4�-eV�>�ԲD��bi�fz}�`��i��q�t68�B݊��+��ʋ^�r�T������
�,PȽ{��B8��H%�7u��}���#%U�ǩ�<Ba�C^�rJ��%�X���FB[#�YV)�c�Μ�X�t�O.�1fd���dg�X��oBV^z2�W4��Dy#���}DE�bI>>)�!EN@��EFR$���~��	1��=����I<|�΅��@������_>V8���.jEҠ:Ȍ��������5������v��?���"�cSH!3�?��r?x�
HL$ٚ����/����ӷ����B.J9�JN���%(�߹r��q�=�&�k[���.��w��'�k�a@��d��:����Ur�u��N���M���#�z��0<�@l ����I���&��"��;Q�K�ub~c��S��Z3ӵg����M�[�AB��6]�;K�aü��eqQ�
 �.o��s�֬��q�!���=��d8OB��v���Xi�u��5N�[����6TҊw	L�A��=��X��0;Q�6�(Wb��'���������C���//���M�%�ށ~��?Mz�5�fu�ʦ00sQa�><}��3>�-Xr�O�7LK�U�|H~�lV� ���R\���M�2�fĄ��o�0H�Z���Q�L��z�!n�*�JI��1"126}\��u�h�)�ON|$�Fp��]�����7��T��8�E����g&�j� 6ȏϙ��D?Wiv*��L62=��əY��G~����xjְ����Ҳy�6*�c��IZa�#�6'��݂��A�A̒�H���d�o��&��pf�dL\e<��a��[籽����PBV����y��-��߁���j�A�jj��{��0��b7����L+����%�Ȋ�6m p�B{�YӚf>�Zp2+!�h�dI��D�T������Fc�'P,�~^����(��%�M���_7���}����3Z�Ĭb�7yz3U� '؍�'��-R�P/O���NȎ8!B{ww��GG��?M6�t�)c��C�l�_�G�41��%�<�jD��7VfI��)|u� �u-�
 E�bl�����H�Z\h �v[�MO˾�����-
K�I�i��� �����qN���Jv��ϝ�����	�&�t��Ɗ��.��.�������gV�p��#�P�9W6�(���KYWJ��Y�8�g5]0҃$h[�R���C#����vp��)�Ւ�E+Y���/-Ɔ���������y)k��ࠗ�c��d?�X��/ae�\�ŕ�PaR�̎�Hu�0���9,�;	d�����dق AXJ������H��@X���V��֨%������dM6H"�F&�	�9���!����$M��*�Wa��J��	����IY���v�R���+WW�=J��Ƿ�q���H����3y�1����8��DqN*U��?�47�1�=���Fؘǋ�~�ݑ暄e�.��%Դwc�����8��jue\ZEy}'E��Ȋ���8��դ��d(n|�b|o��=NJy]'�c^����\@Y�����wɲL�I�Aq�p����.GWbyiV�M��$Ҝ�"�j��𠸔����Qe�R�-!��	!�"�6���upTc����pi���=�9���>��Sy�8`���ڗ����Tf2Rⰷ��F�9I�2�Rvb9��(d��~t���2�R�q��I��%�dBVyM�E���K\�����j����21=�P�⧘��������맑M8�c�-��eОE;�ѵ����:�q*+�o�b��].!ˊ�ӆ..j���'/P̅,H%��kD^V&:���Z{p�$�����i=r��Nv-�۹�YJɿx�HvOj���~��q�8�E���N�&,���W_�A~j8J
��aZ������K��@�r�3��^�njp���l�{�/�7�vm6O��O>������Ƴ9b�>R��_~�������h�B�����.'x���W��>�jAI~~��������Ù�||��Ε���>����!�u�4�5�8�ݦ��#�1b�I�x�x��O���h�ɰ ���l��EZw�"�]��P�:����"-)B��Y(�j�G11G��5�Ei������T�#�R��yĄ�i�A��F��k���_΢%Q�5���m���[�s���G�puG����8~�(��dU��X&Ď,l�4?����ލ3bC��Z,vmˁmȎ�=M��F#I�/�9n�`�>�Ĥ<so�d|��R��>WV�u.��Cm?0:�`������f㡶�n�]�l�� ૵!kvz87͸b��

��1`�M.�u�U��U-�+��*�Ec�+gO`�� %>�,gJ���`)��?�I)���6~�2��t�e%`�lG��v�p2A�QH�b�Ls����/��Aj�*R"�S&�����3������iEP��C�p"+�����n���&S[�.�DhH�B�0����p�A������'�롵���l�	}�x�r1<�h�dS�k�����;7N����b5b�Lp�
�J��&��������Zm�Xߦ'k�FBx >~R�y���o�>��3Ȍ��˖vlom�`߸z�(�~2��G�J����^>	�����JK�lZ>�Z��wUk7�3��C?� 8��k:��R��)Nj���E7kQ�%�Q)ϡ�wHsJ5dY�1H	�aanF�]�蒢�4�/241M+�����Q�>ّ�I/�x�F��Ӡ*��%�k7�$�{`|V�:�Âi�1PRS����D��`�����\rSۄ���vM�K��YO���c_<~�B���ݶN�R�ٹ_Y�Ҝ�長�Vc�Fh�'߫�E!ӓq��ǕJ�%�����/O��9B�.�?�l���i۪�oS�jg;Y��k6��>|�p���d'���b֣���Ik�$����T���$�6? {t��.�:��Am��ުj.�v��	�USҀ�I��b@��rvqR�#�����"���p�����0�h�0'�R�Ѥ[�9��O�;Bք�	krG'Ⱦ�ևu����
�F���u�1��\lѢ�\p�Ni�h%�����<u� Y)��%�Ml]ٔQat����tW�s�_���
y�v�4��h��q�����s�K#0�&v٤�L+ �;���!7-S� ����7��MdM.("�b��4�q1���f� Kqvr�}&M�D��3Ey�ts&+��.�]�Y��%)T��W5�R�����N�������./[�e�I��<ޫ!�(7Eu�����V��$�x� �|Y���L�>~^F���T:���W;ŨN�'!6�_�����M�i�����L������}x
�m=��eY	�(�J�r���5Z��)с�x��bsׁ;/�	q{H��3E�1O���n�vU&�[�],��$ˢ87��O�M����n��8�����{��|�1 ;���E��(�W;�����P�����$6�Ny�"m��4���9��|v�i�n(�d<�n���$�/]�(��Є⣺6��H��[(�n E���O�݊z\.�Q����WJ�E���H�l�o>-GQN<!$�?�CVR4��a���L��I���'z���D�r�bp�4��P$�0���'����S'��WT7E���������Λ��X�ܡ��ů>y���>���1hh�AfrY�=�l����<�k���"���G��	���PB�E8<w��������M.��a]?��f�3$�+�́��'-C\�%D�#�,kjr��� O�z�fF�(Mc�:�g�jtg��h��Ī�Н�7��00�3���dc�݊*���{�ѻ�t��r9ɡ��(�A���-����Ƅ��MjJe���C��ؠ@�'� TI�W��3:��`xf%�ч�q�-��Xs�1���5z7i!%#]X���Vh�vB���d�,=ka�Ax�����b�@�זNWi�.�d�4��ŜܼAܤ!o+�x�\Ê�p���w�Ɖ�L"�Ɂ$�|��dʜ��>���Bք�,<I+�^���e�B��8I+�	�\�,i�@���!V7/Zm�ޖn�[$�!1�B��ѩ��,p-�'`���8p��e��+�����:H�0�Uzjb���:kp��t�B�OmD�	�q��db�1>=�R
R?�@ąxacsKk3�E�	�~���v��˄�]Z�4W�v��ݭ��%vڑ��o�M���Ia%�����2��RE�� |��J)8� ���O��M�Ň��f�5��o�RF�����`��ek�����F1�i��0�E�#����q=�X,&�I�V�l���B������L�clFZ���f�&�r~��bّ��PQK
�09��7C<��KM�i	(N���N��8��¶�S�}�073����c�ſ���0owB�
�8��
�#���X=i���D��b�8Ş�������Q-,ɦ���.$FEb{c�Q����]�6u #)N	�}B�^0�U5�h}Cb�}2�9�讯^T�0-Q��O�0��
}PU���dx��p��CDi����s���A��*ϝ$.B��?�A��&��p�I̟?�Uvd�58;�Bv.o����%U;���DU|���t��RJ�&�e9��#�23�H�GY�������G�ʤ�Az���ĠU?�&
ŭ�rX�ɓ����\����i��;Ўt��{��+���5�?Z4��[����M-(#�����Aa9J���0��pi�3�d_���o�\�;��=Dؚ]����FM6�8H����#��YC�
W9���u�j�$�y}�e,a���w�ܗ�E�H���)/&�m�����C��&��|��S��i�CS��ks�e��j�10:���	��V
򒵃P����0��5߂��R�_!�ֵ��
�w�d|=\�9���DZ=�%Nd����ʲ�wG�P�wg�&<��&i��R�ϥr(��kIֶ�:�'Sb�	T�|�ʶA��$�BS���g3^���֮�&Γ���rom�
=i�(��J��U:.{Ȳ�v�C��I�������2?R锘P�2�nZ���.m8��Ǖ�\����q���#}+����Wo�'��Ƙ�@�+����2|��a���9�xAn��Gy�2����F��������8}�������B�XFt�&ℭ��_t�+�J�%�Fq^�Z�4�%�E);zTۆ)Ѵ2W3'"�dE���Iy3Hsq�y�s�P����/�u1�l���"�"�(-w�[��	O/��A�	��
���<�,�jq���$�Ĺ�T���K�� ��ǵ���s�>{ZoOW�D��_=������e _�!cBNJ~��.�>���U�r<ȩ�<���l����W�����SI8���Z&���_Ge�M�q�~��}�����%d�E���s������D/�ˍ3�0߯h�v+#�(�������y�#��CP�?����7��V��;�'��`2����}�dF6�aл�|lx���X0�V���pZΡ����ft�M�c��!��愇5�&+s�������v�Ѣ�w�y-〄#=)��L���16�m��)��,����x5��M�5���$28+�Ȧz��C��-'zi
<9_O�h�ó�p1;�p�(�Rf�1��P�ޢ`�����n��S=�R(��^s�glp������S�3�G�E���t�vh鰗2�Tݽ��[�͉�	�XCTto0��%�S��J�0!)
c���$��@�n�BVf<6�� �-�˜"K��'뉠u�($H�A���`EVl�n!������$�橋���#�U��ߟ;�/$G�Fz�7�D]�@yhrBZ���u��,�v��I�>��E�/���]�FJ�=�4�-P�,*�"��e�k��9����(ܢ�f��g�P����ǉ��컻���fr�f���.�������h"[+d��7y���&�c��Y��X[Z��7��52Wo�H -s��x�R�W,��`�T�ȕ�`��s�/\X�O\�e�a�1�kt��iE�XJ�9���+4q�+�{Gix�\i�,U��fhӋRp�d��MJ����J'���^͍��4���;1���.��ό�
��p�NK���EnbJ��6	�/����H?����eD�@��ԭ�:|��� ������Q݀�z&�m�m(L���o'�ە�V6�����[��GO(F�� cA�'�i����>�!<���fCek/�G'4���S��}\\u��&���<ù٪������_k�^����|�}�	�OT��ʠ�g|qc�+�gg�d��R�%�s�/�ۈ5���Ǻ��ae+�@�}��V����5%�NNF�$s�0�%)�4u��_��|,�*Z���'�M��Dd�r�����s�Ɨ��!UwS�(��B���	��-<D#?���l �(�2�nN�G赦�-
Ւ�'\I3ơV�yI����&�t��@N2G���:n?���C��j��h�A
m���*�v��N�Ɨ��u��	��4|����=xi<�Q��) eF�Vj�R�J��"���E�H�L>��l3�3�F��Ƹ &�qNF��n�����8��&����'��P�>�]�r�s��{�n^�9$]�\��0��>����A�N���,+���ty�\N���9G��磵��]���8����"54��m����M��
S�� I�I�����^BD0����%�-������	�n�8��>�!(�L����b.ѐ�d)�c.�Ȃ+��<E��F�3�y{�MB����P���)�ɾ�9�[z�t�Y����Hg��i�ޕ�\mz�%��O�b�3��u�8K;+��2N�ee2.4�/�������W��R"PC�*̊!4���/���DZ�I}�?�k�<k [KG	?�K�<Ku-���*�Dz�,�vU;�KKv���<'��<�|��ѡ82Y��ϐ���|���D2��_��@��eR�����ClT8>�ϱ���v�ei��dYܭB ��+g��Z[�L��s�X@#޼rZ��J1a���*<���K�[���jY!�_�gR���o���&G�ܸR���!�u�B��\?[�O��ҙS�'��l���'a��y69Ɂ�6��+K�l���G�IѦ�m4��IL���;����T�T	E�Tʟ�7��t~i�_>��4�2�K��kTvM�ֹ|ZW/<\]����227zϫ�"a'�n���&W�l�FRB�n��%;z\׍�a*sR�o^.�%{���sj	{G�ZB�S�̛h���U�W�B2�~�Җ�)}�4iz:)����	� 0�yΉvJR-&:a���?�g�>![
v�һ�����Umk�Z�Fi/�OL鑇s+��xbfV�iܭΨ�$�l��{�T��+�_��>@gw/�	q�_;z �,1W��d����#+����lEq)I�e2�Y���w4vH�zi�Lb@�߰#?9Tk��v�]V���/r�#���v�ߝx*�TF�R�Y��L~!���P�X\mȋ����'��� 3����	���+{ɦ��-Ɣ����;L�4AZ���'RC�&��%풙��҂�z����Mz�BY|�RC����~��mZ���.�΅���`ʂ��1��.�{����3d�kH�\�fr�&�������@v|��,��j�k
�;4�˄���qƏ]=���k����&J�����v�sK�.�tBuK��NJ����dER��c��F��eNn���տW�B(��7.�hZ���G��+:�9���^��IZ�� aS�A����I�;�Z��\�����h\�O ��&.�jN��w ���x�,[�z\��H$'�zP3�ϊ�i��Cȃ����t>#V3��� �k��\n���j��=��Gh�"��R����')Ix>���Q�j��I]��=�l��e=ΐ5y�y����#cz�ԗO�p�8�����n�uj����S.x6N�%`���E}ٗ3�<��؜�H����_<����,N��G�V�ԫ4�$/h�$ʶ腍]|�F�@B��`d'�7��g(�����ܔ�vv��`Ma'�����:R={�ء�R�rr���d�����1z|�-_z�t�
.��!91��c2Y�]�:�Q�9���Μd� ,$��֊���Po��12���9�x�Jg.����3$03�O�!�y�љu�3FIN�N/�J�(�0ˀ���Z�c2D�Yx�9�o��8Xz�I��=��>�<>�s$�[��_�F���0M��g��(Զ�
V�9��à���]0J�����ךM��Λ���j�4�q�ĲmdM��s�6�rd%��^rĆ�q��'`j�7c�@FɃ$�䨍B�@?��u��+��ּ�ąa�X�ő3����P�Ec��OZ��3D��3b���V3`� ;<$k
	@bl�nmn�F�J��Y����eh`��[��s:~9H�X������32�	� /�<_�Z��s@�n���p��	�/��:��|�=�֍��p�c�g����I?ƪ�^� ݭf��RE)_+��}�J�;_�//o���X�х�i�!�Z�F;��Bq�6�u���Y��4>S+�H*9u]�0Fq��K�H1YH�Y�ԋ��d=丱�%��%	x�kryMd` *�����dS�ds�zv�V3@��Ba&�z�D��4N���NDy�:���"���$,r��5�Ə6w7�!_4��x��l=�T���{=��&+����c�J[a�J��Nl0��q��q�]��+EK��.�ʥ��3.���B
�^�����\E1��������<(L��p��v����r�� �z������e9o����eđ�om�"2"?��Z:z���R�(�,�in>��~�v-��"��?6���@���K�qA�����}h��I�xI�$��~�z�֔�3���w�H�'n�%�B/��7�I�J����L��������}蜜��w6����IO��h���A�����nh>I�W���{�D�e�G�P����������ψY�>�z��yJW"�HM��ҒE�n�+�W���O��/Gz�WzBPd.���06�"��o[$:��H�	���I���<n���%Eyz2����VGgW����A	���l�Y�R;ř40��#f�~����N�@�	��� ��j�e���1���}#�j$���;��V��E�^ݣ%�讣C����IIZ��N�У�$�*�&��4�A6�'$�V�E�])a�D5�᧹$iё�[
��&\�y;��r���ZD��+�.z���3��DG!��4��E�S���!���<q��J����_��?�
�~�1V�=����4�˿�0�����Mִ����o\-���8�1��y���]ݓx�lm`؛,/Mw�JsanW)���P�����,-�H����NΈj��+�)أp�%�S���O.}Y�dk��6ٮ�`��p#�gϷ�^�E%��[K��\��b�zl�$�u�Q����4��^�2]��QC(,�|�t�6j������q��u�+�IZb�l�S=@��!�^/L�����'����y�B%�&<o��:'wc~��:���5�R�:�yj0!
��8+	O������#��ӜX�Yv��T9���*\.)�kZ4��uO���>n���eȏ	D��8��:(^M��,���gQ{B�ZEc���>�WN�yY�N����\�Х��d��D4h'����"�i��M�PB�k��R&]r>K|�O9@9BB��L_��.'B|I�6}�E$�Dٷ(�R����RaX&�x?ă�V�=���Y�X%�I��^e�@ /-�2IgK���}P7��Y��29cˌ�\�*�Ci���4]/��j-ٲ&���1=ܙ7�'+ծtix���D
M������pPqN.=�fra?��?�;h�^�#�R��~���&i����� �I����4!�%=�����P�:k���GL��c|�T��C����LK�X����TMG���x�W�D5/E���px���A���F�}GdA)�!��mp]��Z�K�����O'و4��o�ƞ� o�Q!w�Li~��.�� b�?��:ƨ+���ǅ�#��K�C;Y��H'���� �Ek�}xRi����	�Ҽ�98��PL���:9f]2ٓd���A��Y��������Q6�x��(+�q�L�"N��D�	PZpB��R�hwì�q�$|��G�-d����[���q�ݽ�0Gz���8ww(vV�vp�*7<0�X@V|���TC���zɉhS�	_K�90>�S�qRWϡ"�Q�4�O�(5Q$
��S��0=���} Y���������i]G��a���I�GSW?b(>�?n��b")&
5-}��$3�ã�D����Š�����+'2���&{7R�Lԓ�Fy�eeQ'5�:p���;*�рKder���N��wNcc��?/]�7ˉ��N��o���|���0��{�L1��$&�����rn�/F��*j���w�*�$���EL2�>�W�7����̸��o�zO��1@&+���������{W��I��@zR��ww��3����P)�mr��o��Ek�։S�+e��2��]��bgRT�ʾ���{M�h�Q�}��ˉA.&<O���pʂ��~�����׶�au �����)�}x�${������ԏ�� j�mW�]��9�����S{��1 a����;�U#	��\��o�zNo6�o��:|S���p�ӿxѤ�@?O=�_ח�彊v~����D��$��P^ۡ��M&uW�><)=�V�E���NB�ĘP44w���_~�f&'�l5���k�V1Y]	��X��7��
W�m��-��U�
���BhX0l>����9�C��`coaa���	��{���V�d󽜏��IB���]�G�4��5��� ���"",�/{�i
�qJ
���p]t�'�VI	S��3K��?=�G��d'RfjH0R���ɿ"[��£���`o�$�;ȡ��	qHKI�3�%��/�ןT��zj�ߍ��4һd��l�(;%)�uz��D�F�GMW\�y]����$=�+ZІhA�]�E,�`�0�Nb'�����N�ig�i3m�N�&]2I�8^H��lf�		�о�B����s�#0�C����}߽��{�A.����k�TS_���V����&n�T��~k����������c��pl�^�T����_]�M��a-t��˛M|���#����K��p��#B�MRJ��0ӄ)�^�gGO�?�ק�C�r�ڐ�4K��b��P�P�3 W��b�<k!%����\�t�.���\�v�-�2�O^/+�|�V�eS�E�N>R��R07�����	�xk�\$���rVC�Shni���b+���t2:�ߔP�LC\��61H��<�\�Y����'@�M{�f��@��䩉�����C�/�c�fxi���]�cL����������i��`Vk�ى34a�P���R7�[�D�QL;^���Uh#�s�x�2�z��k=�+����ԛ��Z����s��EM�!*��ǧ�@#Ģ�ĥ��|��f)X�4����i1/�ghTŬOT�R�C�d�����3���V>�ʥgF
~�/S]���Qqc?g�|��&tRn?j��o�j�xV�*�꧸��1��`�v�&�����i��ʴ��I���Jp��55�t�#��`�B��&�e���/���aZ�`�|q�����c'�b�0�?7k�0!�?�qhI��R��8�à�������v�d(�)P �;(ЊY��#�P� :?.��v�~�K�i7��I�DrP�DA	��I��NѨ"�Ni��\+Tj\��<S�~��R�)����dKs<$��S�/):��!�$1OL� [}��O�1]dp����Kr�d���T�W��m��)�hO� }T�Nl�k	���5Kh,!��#�����?�FPI�����~=�KBY��h���!44��CJW�3�S�;��6<�k\̢�+���]�XE'�$;�R'���&?�H�S�M����Ӎ��tܡ#�a��3?�v4�ݝV�S��Nm+2�������gل��A�y*3��QR����N����9ˠn��({�Nu�=�5KBq����{�V�����EE��1O����|��>���z!�^����W�		u9�����u��Y��"�6td޽~�տ{�c׶D������bl�n^���175ӗ�_��o�K��v��������N��J/����߅���x���!5Ճ���?�m���_-#�:y�0��ػk��Kk���?~sDJG�n��(	�/�Y������ؼ|1V.ˡ��1���'/���z���F��m�E}��k��aQR��W����ĕ��8s�r��q��hJ��-�u�\\�,|�2\}Ѐ��t�",���-,H�Ʒn� v~b"QV=N^�I?���I4�y|��#�Vt;�7�܇>���p�0�=�W(Q��f� 6�m�)����as0�ND�V�ɫw���u� ��g`��||�,<<�����lhWgWN_� �����J<�Q]��.ܩ���3�}���mbiR:�}���4�RpD����~FL��	a���EoBGWRM�����q�	�d ^�~��D��#%Ճu23�~��3�IMCRJ��a�`I�5H�,*6ʗ!`�+�#ȅ��DDФ)q�ԉ�=%p��/H���#�9N���H�g�a	?�)'6�~~jj
��n?#�J�HÒ�L�&/�K�L�W��njrq11��m�6gM�Y]��	��Ą��.��(��rI.F�{��GMm�eV��}C!��Z�q�qS�-��v�+D�^a�"�fm������Eh��DI�"8��.��TBt�^� ���1m���֬h<%)��{܈�ŋ���hl?UЦ� /1�XO4U� �4̯��W�N�Sʵ�;_S�q�('��;/,�Ar|$��zy�#�w��)Y�8�	�|#��D�x�*�e�R��u��)�}�T��J�r���`����I#�%�D��-KL��A}�ɻ��3/�����ƘEQ�L��4�I=�nYm	¦�~<��q����[��
Q�[�xO��mt�{��!A�h��滄�߸������l�)]���m�(_�����c��T-��O*T����ؿc#�W/5d�lj�1&���U�N�!��C���q߀��'-� �r:��0j��Tqk�� MZQ�w�dƕ&�#�;�rsQ��;13g����i��*�[��#��
#�{�߭&7��9?J9����9D1�Q��wf�i�`7��i>(��u���.߭E(���eg�����[z�J�H�@2��]N�*�H�c�\On7�5�j$�G�q���#;x�ݖSQ�!�M�qs�y�8�4и
�x�45����oO�h�@��]*gK"���;�}y	F�J(�% ����6�O6v��V�e���!�O������$�ꬍI���p"��a�͜��W��t��+(�6�/W�NպbK'%�v�d���Nɛ'ӌM�8Kw^I@�܁H��7�@�uص�9�EٍKe��c8E�"��CA٣�v{��찌� �ڵ�Y�n1<�����f|�54j�V�K��_h��1����aC�a��Y��E��+�������s�:Q�-� bg�zk��iT�����=�wrM����Y���v�j�'/߱&̕�&�*>nj�`�υ��LBQnFi��u����?������J�ݮy�:uE�+%����m�5Mt�1X����z��"�4cH��[M����ˎ���e��<���k�M�'$ԁ^�蛡<���.� Oba��X��r��`��p�M�ߵ��\�m���%�a�Z�)�`=��VZ^��]�o�|��5#��޺�4Mz������RG��� ���ʋ�0s���)���N�ӇG�]8�c��i��}h�K�vw�b�ܨ��ΑWw�Au+���˛����'����#e�!�w[T��_~|���_?��"�$e���cV�'2Z��NG��Jk)8q����DXk��r�H$���M��Մ�DMt���נ�AzL��~]���ڞ�E�/J�ї�Yǭ��l|��%�;.|����MI�'4���|t�>ʅ�݉�P7c�����h�g�÷ Cjq��Ó����-�4/�S⬙S���M��2�ˏ&9��y"��x�?8�9���$y�1>6CS��N���@dAz��@44�������И!/�@���!42����;@ ����.B�Vw0:��Ϗ��s�"�������>JO����6�o^l�E���^ڽ�M�z}s?T}R�PdB��!H��+�E:N/�[LR��6���>������g��%\U�BQ�>���LMKGb\�	�I�Z�F���N�&a���%�,:�e�Sb@�f����j-��Z2W���#��]�A��5a6�'��5�3�|�U�DE2F0�di��G��H����C#�P!�0/�?H��^�O{(�塷�3RMIH�e�ɯY���z���O�~�Nauq�:��
r�<\���2�'�_3���n�߼]}}XLHy����1u�<�K�?2n���h6�S��8#y��H"r�xPg��l��	�J�5ַ�K���A�[V	16p�VM���i,���HM,2���*�G�-�+{}�2�pћ:�@�V��x����Nс&�~ƨ}i��n)6����oy(e"�b�q�t���*祩S��;�{����h�5�U~Gu�^*�fG����6����m����ً�{��t��f��b�^Hs>�s7�Z���/Λ�t����?}��|����62vX�k ʲNZn�Oա�A�.�VUr3F�Xn���i��<�ͪ��A�j��ft����d-��F\��Y�c.	T��7�)K�^hG��!�X����Kq4/�7ˁ
Xh
υ��
����0�:�f���y�mT���nMΑ;w�>�3Ȫ���ƟR��k4O�N�����l`���O��Z,�����]���K�J�$��h�ʽGF�Q�8�|��Ճ:��X�k����`����PW�d����Q��@��Ԋw~�17���#�&�ͭ=����G��s��y���J�zZR7�7��'����`Ф���r��#����О����(X��?�2�_�N<;=b,v�\ u� ޔZ���,����������c%����O�#c029fܬ9�Y1p
x>�O#�{�>���,�ʦ����E��������9AQ�g��-"��(pU�Vm�w�s"�'_����18fp8�k�~e��UO����6�hi˚%��=T�6�O��}8�}��߻t�**���O�������^�S��}��-�G�nT?uQ�<��K'K�V�Kғ��2'˺NCi��^�D/<5.V䡟'#��^c���p+]� ���j�C�nK�k�ZGW���I-������/a�'@����}�'KY޲�+���B�-A��W���i��]��r%�*��%���s0&�'�=���VBRAgF4($�����ly�t����$����/�Xgؾ�k1Σ�y6���-��'.2�Þ� xx�ނw?��L��vmEτ��{�JF����kG�'���C��$��Y<"�}��>�2�����-p���&���M���]����8v�:j(�Q��K۴2t<��m�чx��kI�"��J,/X�/.W2�{����XS�c��Y錾��jPR��eO�ܲ�Sp�������!�ç��|�qh&����UӘ����D==HK����{��CR\���N�y�J 
��a��WˌO%��Å����0����o��w���o?G�s
��>,�C����:?��G&*���ްZM}s�B���w>�wz?��Dav&f����7�����k��Z�B#�������A^k�UM�x�1F4%q�ŋ����A��3go�;ޏ��Ip�����{��jA�� �]AƖH���H���a�	��.���ܹi�.7"�%��`��s�����NLA Q��s���U�22��S�<P:�Vb�<k&uH����������Hz>{�ߚ�������&ЂC��;�)Q��on��j.s������J�մ�:Ӯ��0� &@�:i%&0I��v��EɘG4Os��ӄQ|���a:c���M?:&�q��z[:;�(U�L�wI�C�^ݝn>��D��wӿ�����@7����\W�	�g�&2�|hzCk;^\�O�<�%�zU-��@�qm_����y6ҧ�ӫ���) �p7�te����&cq&�x�<���#^__���i��Ѭb�k�A�$�/]j�:��e5u��H�o_cC\ԫ2J���vo��V��osg7�G�,5?��.7g����!��C��zY�AgUD�ۻ��f��҈o�-��W��)�ӏU=�Û�׃ቱ:��Va�3�������6�VBdWnU�<��+�8�m-}�j��.�a,��ş.�،9ާ��߱9��~|�wn6���R>����ś�hF�KR�X��Q��T��5e>n�Є��]�Q�c
n�>f�+��2���	�6��[�]d6��Q��b���oW[J�3�J�*1�`B�	|Ej��jז�����W2����Ҭ���8��s�ם�o7-:h����bϠ/( ���������[k��ڧ��"E
��k����|6`�S���7�Q��T�T<#�JMq3#v���ߨu�z�N��J�ω�χ/��i��\�	@������_�knx�q�5�oU4cGUhJ���	���ֈ!_�T����ӎ���Ú-�F�K�^�ii�E�>*g����&�'E�oc�%���E��wX�Ȍ58|�.y�I�;�\�k5y�"��S��L��v�(����7xg�>�h.\����+�H���B]7b���n0���D3���^t=��p;��O�,s��v�����)@H���j��tZ�5.*�_�f!���&>�u�`��������DrXe���؄ɬN����J��{�V\eui�i��,�����+�u�>%�6E�� ��{�GXd�O� w� ����ʢhg��xJn��5v�����x3h���TM��	���#?/.�l�~��Zb��j~IM�Ŋ*�[W��Ѓ��k��*[Uh�5�Hǝ���]�{۳e�@0��4V�\����K���������S��O^@7O��ݛ��xJ�Z��l���ϣ�&W�����=�x��n��/��҆���@EuF\�qh�ua=ih�+�������N����p~x��iWl[���t\�����E�Pq߄�voX��K0���6�����Q�2���:Q��LF�u(g����`�*礧��'���X�d!vnZ���N��t3��ßnX��^F�}�m<���{���X�[�POs8�J�<N{��_م�H�a�9��o�}n��￹iI	�������ǭ���sq1���E��q�"�����/��8�;���0H��?�՛(�Y���m�����}H�>���íg�����ѯNV{L�w�2�4�!Q���y��#Le���X��}u��CXC?���h��	o�z��8JW/�s�I{ʈqx�;ڍi� �O}S��	OB�M�ۋ)�@���x OX<:��y�1��υ1g8������7��&n�y=JL�3Gc�~����L�ET6N$7��L;����M�����1:cҭ#����@D�Ϥi�b��~����tc��LI穘� ��D�%��aL��'��ٌC.S��1����K�j��w�/��A��ϙ#*��ώ�:0�?S��,�����e����;y�A������	��%�mC'c��i�e/��`o'�C�v��\Z��a��ġ�Q'�g�"B]�� ��Ց)�p��'��M��X@�����_>�D��a����~�\��N�R�&����ET����S����}I��Q�hb&�I#{'_/���Kfpj�9a���n��fRG�A����1�����Φ��[͙�wL������Q5�hl��V˹C�0�:l�1�Y��
�vʈ�����\x�(�����ǌ(w��9"q���]�{�1�����y?Zf��r��{� &�q2:�ol��f�bL4�"�����K���7v"pr�"����t�,N�����+�s������x��3�,(���/}�M���n����U    IEND�B`�PK
     eO�Z	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     eO�Zd��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     eO�Z�Xw�s� s� /   images/49baae61-cb81-429b-96a1-6cfb8f124b59.png�PNG

   IHDR  7  �   �&�>   	pHYs  �  ��+  ��IDATx��	�Wu/^[�3ӳ�fӾ�F�-ll��1$��;�'���~�|$$�@H�%���9��`0��Ɩ�%[�-K#Y�G�f����ޗ��z�ܪS}�%!�,��O_�{�k�u��=�:��0��`�#0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
Ln��`�+0�a0�1����`0Ƽ���`0�
LnƼ��8�/����#V���0��$��0��������p8l��i=��j�\N�O>U˲�L&��f��唀���w�a���ٚZ*�[�U8��۶M�F3MS�/�`��iZ�_���J�H��u݂u%�,�0�R]]�����TSSS��ظ�ڵkm F��`0^50�a0�z�)���=2::*
���� ��,�l1��{>֚Jf���ԛf!�8vԶ�0���������R)X�K��S2���zER�!�qJ�RR`+WS��F�4E���pT�<��&e�� *��	�"a�5C/���em���9�P?��@h���_��Gft=�jk�gkkk�`Cܪk�+vǻ�p��u�
��x����`���LC�)���Q}||<8�L6�L��f��xb&�M&�=�XK&�[��fہ���h�L�ֲ�0#�� *�8����n�w�������Ă䅾�P��Ђ��'��jb��E�c����a))%�B-���?UU���S8|����)���>��\$����>2��I���d�&�hji��m�o4�P#�x�b�;���_Ln��
$gΜ	MOO����Լ|�k_k����J$ҭ�T�9�ɴ���i�Jg��k(����D���l+ �@��GW$$H6���B����i��T��|� <Hp�x2����
�߸�C��q�@ ���������M+�E=�����C��X8�
��Ñ�T}c�XC�v�����M/_�Mc�+V�����`�J�1�;4�0j��D�������['��V�%fWX�B�i���B�eY�}-,1`&! z�h�����@xv ������O���b=�KǑ56���
rC��@�>Q�Cǣ�H#��l;tL�d� 7�YBҦ a�?��9p�j|<��|O�@2
��6
��jjkG�u��O~��4/�iYؒm�mM����6m�:��a0�`r�`0~!Ȭ4::	 �Y��o|u����T&ٚL�W�2�E�|��y���5��f� |�iU���x���kT���ք kOp1M�}��ɑA���k>q��˟��Whm���_.%�WP\�Z�Y
8���1��H�����#p��b.�䵌�B#d铓E��q�z��Hx,������o{j�XGg�ضmۆ���&���]]]h�2�u
&7� !�?~<:11����n����R��2�Juer�e�lv)H��|>WcY6��,��A�k�9�B�B������Gh�m\�_���}�����Y�"���j�K��2���b��������&0E+k����cym�~��K��ר��i���� ��dR_g�5���944�9p��X(<[[[s���q�����~��cK�.M����,Y�W����0��AwϩS��'�����[<6:��\.��P0�l�j����,�2�n;�_G^�|kYT���TiDׁFS5A� �$(нm�*8�w�#��1!2��`���Dl�5E����ǭ���ۈk���!SZ�1�GnȜ���x��)����#H95�bC5�d�m-�1r;�W��{0a�*@r�,o���1SG���E��Hh���������t/�w�碥����Ln��!<3S�������Ư~���FF���&W�3���|aY�X\ �6V(�1�Z�PȒ�MB�'�]-_�2�K�3� 7��n�6�Y#��"2"G@ѧ�W#������վ5�KU_TDJ�o�v>b��ST��D��$b��-�)G���]���»�$�
��O�>�����un4���q	��.
�h3��5ΜcNONΞ=3�?��!?�����{�w�����رc�V�B?Mg�+0�a0^'@B3::����MgΜY761�6�N��e�+M�� BS�2�cȵ���cq�f=��p�D!L!�A�5;�.��"�����D�@G���e?ܖ�Ѐ聊���Fv��v���.k^\�u�4�XAl�^I-	�&ks|m�w*�>��JS+�]$`T� ����D��KrBA�zH;&�|�w�Az���}�����`:�������_v�ԩ�b��d49���o�h;���|����˧`���͛�W���c��35�}}}�ӧO�~�K_�z���Ԧd2�
���N�	$����
Uv�E�E�UJh2BJ�"D�K(���D��IJm���vY#��B�G��Ed
�F����i[��G&
2��&7����
.o#�����<°���w<>��p��Ne{}'�{9u�IX�V���lan�����hʲ�B�*���9�D���8��}]Ŝ���Y�=�ۤ�f��n��p6�o�{�RU'���>u��?��Η��k_;���Kǻf��^�5&7�<jg�������x�������GG����ήO���AN6y���
d2��/���
W����\����@PW¡��Q��]�Q��OnP#AA��� ��(���`6)=H�`Wi��=���7cY^�a�#N���H�:�A�JU��U�GF���¿�	�`H��7G��%d=�k^BB��*����>�G+y���Dֆ������������I&�@�5]�vQhy�~ὀU��C�3dR�bmA����Y�U�js�B휑Z
����9y���C�ښ;�;^zꩧN�Ituu��G��Z�c�q�zz��|��ԩ�����^��RXV�p���!���y_K�ڗjGY�����X��Ǖp8���ħ@\�l6fN|��Y�i�%����- ;�h��-M|ZV�#em�A6�TGGU��P�#��m�o�o5����gu�����"�h=�!$Be�d�:Y�����v��*�� V���l�BrD�զmzd�#tZ����<����7��u��}����u#�/���K8�H�O�̬���������=�_ll��Y�l宭��M�uӦks;��0�A��ԩS���x��ӧ�>��_299y-�� P�r��4u�dB�W�`	a�rGV���D�-=�P(䓘��6%�)�hT��4)�����Rff�yA2�N'��؂�
�e@�M�$3�7��(��v��Fv��>�l9ނ�*�ЃX���l�l�n�/�b�ۮHE߁t`y��4�6�M�.u��8�|�qS�Mu�H+�̃�-l�c6e�磸�ڢ�A�K$B-�H�&&Ҽ���i�|-il*������7�������l�#�JDG���{�z9�1"�	���ద+-F��855qۙ���b{�{qk[���q��GV,Z4z�UWa"A�5:��Ln��N�<�f����_��߿nppp��@d�8���X4Б����!���	hJA"�������Yhi��E��dfllL��z!����J��б�3�0 C�E��z�%jxPH�"�;�aCl��-4]�`�H���
�`%���T�X����C�º\0��߹��䢑h:�e"�0��#�H���.ה��i���#��2���p.[d�J:PŒcß�A_%\��1�miE��M3�g2�@6���� �u�6�h2���M$��|-\;���7�ŘU*ƊE3
�@fBS F�!9���LM��x"�H$Eז�a��&9H�6KQh2�I�Y����!�dZ'k�<_'�Ta�aؾ��
��x*�z�ٳg=[����~�o�ҥ����7�y���`\$`r�`�p��S��6|���088p]&�� �h9p��B���3�L`�8�YIja�����6�455	B��zP�7;;�LO�ňennNI�R�(��dj�E��+�,��1W#��
��p�Q�������f,��ж".@ZR@Z����D,����@�&�3d+Q__7W__���i(��@bb���ڂa�3��!���)���	��+d�B���|��V��!EƵT*�[�&0�B�Ā ����&#��H��@���%��@?6��Kc6W�C?�a_Ch��f�ղ�r��+]�����K�����QR���aE?�P�9�Ldg肄��/���}Wӄۡ�'�Ϣ-���4��WfR����>�6/<����g�-[;~뭷f�l�x��������1^|��رcǖ���Z���}�Tr#�n8M@2�����t���7�#�immU�$(uuu��(�EM̙3g�ٙ��Ҡ�$2Hj�!�B��h#���(�C�H
��^RIhJ%����t8��s��DWw�@<^;��l<�<��T�b��6"����fW����⽈M ��Ż���C�ƒ�dpjj* �����kNL�-휘�lK�&Zs�|<��5X��P��˴1��f��҅:��q�R??_�����O�)�_�C�+��
�wn�AS�p��0�.8==��#�@pU2�x�����Ç��>p`�3��ַ^Z�j�ئM�0�Ne�#����q� M!G��>����?����#��o)�+�M�~G!�R$�Kd���dn ��d}f�̴��	a�
51��R2����BMr�����I�\��#1&|G�I>
���3����4�6�6Nw.��X�1���<Y[۔hh0�L��x1�wQ-e����	� X檷�{>�(��33�����tn:4�7阚�i�ߖ!Z
���I-.�/�"$~�*�k��T��[ł��x��_ْ銶w}�<�fȱ}�U�(��1�
K#��u@�~�����v�z���۷�衇z���3�?�q!���x��B��k���<q���cc��d��K���s��jz��rF���(dnB�����Nq�300��fc$45Q�>������A?<$3ؾ��p(:��h�o�kni���^8���1���9�����W���<���f�r�����.fV>?p��2�Q�j=���p_��=���0ٙX&;h���|Y3�g86�9+tu��& ���O�݃�Su�� �������;vd[WWǮx�(��+V���U �S�NE��,����K��O�����m���QC�%~��2�G�������O���}������I
"�I��B ��Ba���k#��J�����z ��b�	X=�&���ӝ�m������|�PWWK�ЁĴ�)�� }jzzz4 �j4:����T�O���d0m۱b>�2��>��0ܧH"���=k��]����~,D'e�O��75Q%��_�tQ&3�Y�S���KH�*j�0�@�֑������=��c�/����O��6l�p���kr���E�#�� ��0���������|�3��<y��SS"�	A�cEmz3F��Z":�A�/�@P��Ҡ���2p?�	J&Go�x,
�ƿQ��q�ӆ�PB"II��O����x}���Ovww�.\�d��k�Lss��d�\�6�kph�@`rR������L��o��o�3�L�i��i��V]�*�[�b�e���������,ۊ ���߸.���nra_��Z^�yx����At��ב}x(2O5�5z���G�%�+)�V3`�Ս##�g2���������=���#H��e��
�;v�����M�c�7 �xS&�^Y��(:�b.Ҧ�~3�ƲJ^�Y]D�Æ  ���hjjQrق 4�䘛fjJ�Ԡ����ͣ�Q2FH	xO>�5{9m0�:j)8���MM/uvv�X�lYߊ+&0bi�ڵhR ��������{zz�Ã�c��|p<9����}����V(�ڋ����2�(����a�ڒ�D`�0"�^aR�ql���˓��AU�d����~���Y9��AA�������l��sFv��&=�G�yud�i}<£�8aAOX���]�Je�ݻt���v�ٹ���cz���i���3^0�a0^!xZ��}��wɡ���''Ʈ��o��D&$r�(����!�B�uQ3Co�HD0��A���Q�������43�t��ojg��e,�n�t(	��Cu�����]=+W.;�t��i 5�ŋ^ς�#0����ԁ8���6�e�b�����!ݘ�����2�2���
}�;�5]Y����`���ߦ��9f�D��9��mS|�!kb0d����y����*�#�dd��'�+YTm�\��q3H�IFZ�b �5���C�7�����������466?��Sc����U!s����>Z��.��0/3����l����������T��i��${@@0	�of��͊�]7����DB�����53�T�X��pm"7��@�iKQ׵��j35�5�����6[�|�u�֝]�h��9�y�z��@ڱcGȌ�H$B�јϧd2��l�����.�.uA���=�����m7�~� .����c6c��e?���3������O��*k`�F�d���]a=������ي���s=�-�z�l�rm�3O��!_ʕC�;"ŏW�L��㖏����Yeb437�!�m06�'�'��}6��b���H�x$�oZ�r��<�;�iӦ���V�����x@a���ٳ��_���cc#�67;�F�� ��E�L���	�Hm��Bk�d�j7�@��M�#��Ar��X�A���f�@45�I�su����Ύ@b�\����'��k�@h�דό��Q����`����5###ᱱ��]w��+_,t��� �%��"�Tj�T�$r-܃���|-��R��$W#S��[�䓛��!�
Ѐ���F��3�H]�V�_��6���)������K�,��s#�P���V��M=/���ȹy��ѱ��
5[�<��O50�;�_6)"/88}zp���H$���������ε��d���Z.��8/��0�`��3�<���/|a����W��Oޒ�fV��k��o��z�R��~�lo�F�d�i[�dB_���O\��QK�@�TRK~)�7��M 
 ���L4=�����ʕ+�Y��DWצ��Ж�/9|h===��ՠT]WGF�m`=jQT �f�����l�؜�$�䲅%�B�ö�v8b��
zK@��E�1Jt�J������p��I@u�'q,�
_��e-�8�B���a����L�Bsb�E�=�P����)9wQ9ܻ2N�FY�69�YLs�zaJ���MI�%jz	������1\`U d�V����Rnb|l��@���z��p�}�����ߏ5�\9�e��¦M�,&;��W 
�]�v�?��O]�w���ѱ+a�:tb !5<����O�I�5q%�ݲ^N�ACf&r��p��)V����&�O�`ssþ�΅/�X��Ě5O�]�0���^|�%�{��ux;Ggk�K�������W:��`���>�\*��Q	C7�A�E��AF�����`�d�@ah5��Z,X����l��:�RC�^��s�uT��>&mB�����AY�H^H�c�-��
X����)b�GV���}��u�Y�H�-�e����w,H��T�[Ǐ��f,""�7i�ߤe�}��&3����F��ѳ@���:��������$�ϧ�v����������M��g���P襗z������?���}n��K/�^w�u����xy����%!���z�B˽ﺾS�nN�2���
�-��A��HL��+ݠ�Eē�eqk=Ţ1�4-� 2C5�p�U�("������jjj�B!?�P_?\�X�\wG�sk.YybŊ7��nJl�$�5_4��d�eǎ*\/���������&#�N�=bۅ�#���9�˷��5ؿ�4����P�¡j4M���VQ� :�a���R@	�b���Y��h�d}b0|�2�i�!դQ��1�M[Q$ӌ��Z�y!_`+��ZWx�.��߉�`�-�N��91�q���) 
����ȭLn\Qr57%S�aA���e�����H��|����髤��,�t�	?�I	���+� ���͑�MH�, \�Ui�+�Di˒Q,�͎W����!�3�P�*�a,�	WX��ŘP�(&ә���������{�߿�����u�{���E�%��yg�oUvJ~=����K �q�{��ؿ�����r��� \�s�|�¸剜rҠ�@� [���GorrR�����|p���&��"L�	X:Y�lٮ�kV��]q�ɋI;�o�>|u�5�O��O��d�)�KקS� 7mɹ&�k�� B�FU�Z�,���� ���h�,,�&&�l����Od�Xt�`����W�eAh�����V��#e�%�} �(<g4V�h�����M���x�L6D���W�,f�N�nn"��9���|�^ ��?�[\���T2=R�) �X�	� Q�"��أ~�%-I�ϏlB�6i,OKC���HZ�okYd�� �Z�s�1�H�p�v4L�㕠h��͊ZZ��B>�΄���#=�'����~���?��S.�Y�vm��:�Ln��(���=����~�ʱ����
��
�|7L�Q� ���槑'g�P}a�:w������Go�$�h�v���a�|fB��T,;����Ժu�nXyɉ�V�tuu.���#D&466V���u]"��6�fK�`u8�� YZ���Nu���4=!ID� 0�����b����WZ"�X͇��,9�"H�cΟr"<UhCQ���|2��?W#�τ��s��$�V��$ryh�)��"���)o���}D.,�2��r"H^�RQK���`��K�W���z�i�̛�I�S�\�PNHU���i(��uD�d��kFd���N*Qa���TDrQ�eG�K%/���72̢]�V��Z�>]� �J%���O��?��g��|�G5/J~�����Ln�� 55�v�j��w��ebl�3�s�aN��\%�lV���G�<krN���0C� ��
~ē(Ri9�n�9[:�jaZ�}�`=f޾|��g7o�p��.]������ړ�����/4��l��km~��e3��]Z�k�"��v����}"���#��4%"f��JԤa��D��Y��w"ԗ����fs.󾟊 3�+�K�S���h&�'<r�~�y0�����ܖL�T�"�J�O����m����(��`>���QL���J�A�
�E�8x&#G�v��������H���(�סu�<��Fqo�9�&,oeET�LN����!�S�U6~>�S�jse�8Ƽ�h_�v8֦|���������̡��ٽ��]�;�:��.]:���P��;^7Q��Ln	Hj�������~�ꩉ��fg���l{A�XQB58���8��3�j^n����GA�� Պ����_C�'+k'C��@$�Y�pў.}���/?�iӦ�����2gΜ	=�;x��x�/���MO':�z�����`"�n�aB�Le�U��/�BN<H���ZY�_�tc�D���{2��S[v����5/�pLh0P3��%�#kB����s�f<3�C#�hWw7h��Z���!D���_�<v���$�l��yI�~w���P���H�B��\�����~��6�>��N�ܔ�Jɏ��cT��跲vG=g}u��M���=�9�&��7(�8(��|��˛a��\*�d<W���.>�w����g����/��'?yj�%���~�E�e��`r�`(�6����o��׾����o�7�ATv�y,����I�.�X-G"4_0�
ArFm9�`%m@,Ca��`��l_�~���KW�^q��ɮ����oEB�{��5�=w"��H�����t:��T��k��e�v+\O����b�`8N	�Y5�="H>+�`"����:%A*�~��.�HX��	9�ʚ ۩$�Q}�Ё�Վ�>1x�^����hƏZ��G�%�M�Y\��&���dF6�&ڶ�0��Ne�F$ζ��`��j�
f��$D$��F�`��N�{�*~�a�G�*yZGZ/V����9��v���Wk���KW�
�F�B������؆~�ȹH6����[o��}cS/;x`߳��}�s�333��ۿe�����0�}�і�~�������{��w@�V��~Mf�p(�	�3i��7IM�b� ���M����������m�F&�3�g�.]������nذa�Bfb�������@___s_߉�?��?^�J%.�_�C?,/�X2"�&�¬$¤�p�&�%B�QP	ł����}?�5��C�I�20S�	�KK �AȡѲpv�yn���6B�m�5v-�;��N.�z���^�%e61�-<���U<�Ԣ2���"�� `�$T��-Ƃ�*�#H��*k�L�{��p��'9!e6&b��"0��\/�H�����5T;6S�i��#rC&$�&�9�
�;GD+��Fu���}A���fٖ��T+˿'x��OI�4qm�N%h�_�b�`��b�c<��9���as�$��"5������?�W�Z5
;��l�����0�����}�cW���ߐJ���	q	�0���4Y�B��ތ�W�}�W�7d������OZ	0p,,Ti��ihš�֖=k׮}��+�ܻbŊ$,��Hhb��˱c/�^Q(���viM��t�ﵘ�C$�S�0_��C9P�ܜ�g��N��D��Z(�%u�����9�k��Ie&��Op=���<A�&"OH���n�g���52�wڇڃ(kl����!--¬e�D�.�+���}nd_�ܠj���ԇt\ٹ���dd�ze�s���q�����N6��~U�1xn�4>ϩ�%k��<�ߚ�kE䍶!BG�#j�J�3�w_05&��m�4���Fkjn����{����Z��}�_<r�嗧7o��_�b��`r�x������������o���	&�Ű`Z}M�O ��B�$	9zKF���Ȫs�HQx����9��iX�-Y�dۺuo�~��o:�iӦl�&Kׯ��{���egΜ��`����Z�X�9b��I��@�.r %SE��Q2�YH8�B?�v���J<��wE!�	,��=�5D�߲ sM}r�.[��]��B����
X:Vɓ�r��,��Wx�|���rz&-�]cu�^�o~��|�6��7����>Bd��L�7"�31F"��Q��Z��~V�5)X@�2Q_u�`;�3�$E2�A�E*�
/���s��3.[�[�
�F�{N�`��S�VҞ
�g�o@tt�[�{�C⣔��ggk���U(������w�����җ�tx���3R~���u��9|�p|Ϟ=�>�������č�h55��P��!kZ(�*��B���5���G!Ǵ�Ԡ�i0��Z��7��M=W^y�8���v���'44Է�ȑ�K?�ɏ�!�N�M[��	������t�$0�`TkdH�� ���kƿݨ�rBB�д���j�(X�Fi.��H�����vr�<2/��1X���]�bTHҰ�vG�,�Ʉ#�tP���Pi"4�;��������o�?��O9��r��6ˤۂi+�� d�C�5�W�/i�W���o�2ñL�p���}�d�,�\H�G�@ji���t��}�Ҽ��W�2B٧1��L����:Mՠ�"��a�h��^��f�=�J�{��ч?�O��q�ƾ�n�	�q�͹���1�188y�ǖ=��[N�<�k��]��ZlbjRs�REvZ���5u�*�`�̠�FM���ր&̺�:���k�x��,L���/_��k�ٻf͚�ezB�ӳ�>����|a�K�^�ljr�j˶���6� ���F�6+5.�r�D�ܸ�F8���[�	���"2�a?,]���|ۡ�#�O>%��7�~���Bθ�N���g}��q�\�+2��*�`��lK�(2EV��-�'��j�0	#�k���r�*͇ⷁ41�x>�q*�W�1UaS�ٮ�&QUE��e�9��xE���B�kj��oa?;��E�ʄ_W�:�T�}�k�C�i|��>��)o�)����'�f����.Y.�sl9%����R�m�	j���Ɛ�+�������Y-��l��"<��<���Zg��7�LO83xf��޵k��UW]�R��0�-Pc��O�~��_�������06���s�x��s �r	�	@�I	g�0I;^�(Λ�	�Lss��u��>u�U7�x��WL�i��$�����󞿻�cG��Z4���eж:��kW��!A����k4�_ԗ�}Ad!N�FD�P0���	��2{P���d� 	P�>Pn���	�-��Y&L�p.��MV�2C��+�]QQ��w�r���,��J�Za�����y�T�[6���"��i&��@�"u�tPyV��q���!͆N�R��1z�5�����}��L�t<'rU!�oHCc�4\h�����(�M6A�f͊(6����9�8j�Kv�h4�还P$���y�N��Z1�T/QXMO�td2��ӓ3��w������-[�l�mo{��c�Ln��������|�3o:x��o�%o��]�w�		
7�|e���{��A�=�8^���`%n������H$�RWW�s[�lٶq���L_u5^��^����]����7ݚLέ�D�-�C#Z�f�je<ӛJ�7�D����F\sR���d=g֘0;!�A���mgf�|�*�m�#��^��D�0�T��S����������<�8e�^�|B�z2I�{-Wr�6�!!2�P���	^)?�r���z�ㇴ{�J�L'��U��5�فX%��>,G�Y�H+�L����G�l�}@f��k)�C��TF���9� �wl��rV��~DD��˖]q}46(�̲˵�d��k��s*�M��`�=>.zf���N��*m��`8�����bG�)]���=7�8u�_�򗟻�.d� �Ln�(�������wߚ�/�x}2���l.��
�R	��*ke19RVZ�pI��i��A�ŁŁ���Px
V��[����k�9|�W��]�6s!�4333�G������ґ�+��f6��u�S�����I�����"14ø׏f)W3�:Gn��r)�rx�{��,X�@hk�^2��Hʂ^��p�e�S�+i̪5'�&Ā�������o��f���o�|��d�V�?F֔HcMlSD�T/[���Dv��wƅ���Ǣ�6�y�3������p4��)9��=��.�"͙�~̘-�C�>/k������5��zY�V&�����G�$�I�M�WBP�#"j8��I�$��Z$D�C��ʩ�<<�NYK%��v��֌���pr�jl�4�OOO7ټ1�ͭ���������{��Lwwws��&7��<�Yxtt���޸����g�H��+� #V���e��(q��m��'ri'��P:}
�ERK1��Fc�u]����K�o޼yx����k���~�I�����& r�|�������U#��+��L��E�����u���OD *�Y\W<g�r������证��ѱ�?��쬟�Ld�"Ti��!"�����[x������%P���P���O���B��4��t:#��=����RvJEIU�K�%���2�X�-�I�Uը>�q�n}'Oc��'72��I�!����&/
w�dO�:$������`�f���F�ı�<8�+��#k�^��!Ⱦ6��F�M�#�X�$E�'F�Oږ�̤?ְ��%% d$�3C������&:[rR�JRb@�vm�b����`!�!��:W�W������Y�N��jk�.�yi��'���O~��-��2�^����;��0^�p��s�CG�\�c���������dr	����ry��꿍�[N�F�M�T6���r��BB ��7�aat,�I�����mm�Ͻ�Mo���/Ȅ�������3;vܴ����:��!�L�����^/�V��l>�Jg3yO觡�/N�2)�I��!.LP�=����C���H������˕���K&6�������ǡ�sM��,�-�|¼6�T�U�/GȔM_�&ZHK��ρO>m8v	�Y)
��RQs��唊�(-�.�-b?�J�;���PIS� R@t�[�Ȅc�H�˙�m�8��&�.��y�R��-ԼP�:�>�V��x�T�js��\L��Ll�Y&��T�#�LĂ���v�8�OJ �4���zc򺹹9?��ȧ���'m�_r�q�D�uXW�*k��
S�L��H��D��H��/4C�4`9?�K�`��ݚ�X��'O^/"�9r�={�`)�Y��z����:��׵}�ַ�ڵ�7O�>�&�z۴utN�7d1j�<� �Ŗ��e�E�M�x�w���f]�	8�N�\�uww?�ۿ��C�4�����\/��q߁}o|z�[9rs:�\�7�1���iU�ъ�0�b`z�t�[��QK��9q���C�鴬�A3i�܁��&'�}!V�UĹI���J�6%��Μ�G*�Gv6v�g�B��!	O�>�_.A���7��O2���h��D�"��/��*�� OAq�m[-������,�3�%A�Mi�>ci&	�t=���C��c=�3W��!�,F��Zu�i��p���qM��\M���1i�j�N�d �Q5i��UL��|K��N�ܗ�1��bA yA�*�q�hՈ��̎��[j½�HJϙ6��U���^�7&GT�r�#j��%�>��n�Qk�փ�Q�G-G�a���;��:�N�:cMMMp!�Tf�L���r�d�T�����i�V.u50#��α�q/;Nc�?�̈}��]�m���!/Ɯp���/G�厽��-��>?��إ �����ٷ�K����Qoo��u���+&7��P[3����К'�m���C/�&�Nt����Ɓ2㛜�;�
F]����s.�:�#�|bE�P8�o�(�Ƣ��X���z�����;����7/ȵ�G��ÇW|�;�z׋�^7>>�&�(�M��gA
�rR8�1�fX� 'bR���obbB����$	���x�컀Z����=�����$�dg��dx��N�'�i�|�섐���9�0f7l����e�X�~:6it`��A�·��/�si�>g��?����`�o�\ccc���ٌF�r��F���\��+W�NNN�����E\Љ'0�F����X29��SB��\�6��0+4��6ht��8@��٥0L�&2t &���A%-�0�o.�@�}d6!��T��g�R�����l.�f����tdv�[%-��k���q�#����D5U]�'����E�-87��ـ��iu���'�M����vQ��>(7?S���L�)"��:dbû��1#����gCvȖ���0��G(��N�Ŝ�mI�
F�A{��%�o8{��w�m۶��n�Q/pݸ���0^3��&8::�t���on������\��X��}�/y,(�\В���$�o��l���H�(�[�,L����\�|��ի�������/_�kML���O�����ȭ0��mx�4P���lo�w|M����W�Pl�\�Q�����W@9�V�����OC&%ޓ��ɂ��^�$mW3��&'����!D�Ȝ���8?��(
�+FFF|BC�:.k��7z�	q���p�I۶�A��6g�\�����pMM�p,�[�~y�A�^���1q㴼�������l����@<����3�tP����p� [��:�X ��~�E]��e�2��B/2?"i%_�p8���B�X#���h��.E�*HtI�� ���E�ښ��H4��|�>��$�gg���Ba	P��~Mɶ;4Mo��Zm���θ�]%?8�C"�b"eD(��c������h|�x�>@-%^?i���5b?ʭC�פA��Ȅ�ֻ�����c`���YN��q��I
�`0���v�С�ccc߂g�{p\��z���qу4/�߿�gO>����X(�g�� �Mp�����͋rf HAoq��F�=B�r��`�J�dx$����i��7_�=�yOZ��E,SJ�i�S����O�H�X����y���'N�K6���5,��(.����}Np7�%�ބ+�߈��Z��%iGH�TV�V}^W;�Y)���/�:Ⱦ#D�H�"��He��{w��!���r4�O�`�p]Շ�M�a���t�8�EN���L�`�hmm�hjZ[\��ق1`SZ�x��G�������8|���߀��g["�i�Dԕp-�,�2�/�����=ŐdM�F��A��P�4�#��_rG]_R�Ju���{"B��4u�&���Z*;��KDl�~��[�\z������8x���M2N�8�Z063��셪�/�gx��V�}������,�!;��}%jq,/hm��|��@��"�Ns epN$g}��(wT��њ�n�@Y>	�����	��s��D��~^���o����c�������=v����	 _F0�a\�@'ڡ�����{�7�~z�oNOO�Eu>N8���9�e�&u�(��,C�5"5~�Йl���(��J0��a����lmm���W_}�O��O��������:Q��O�:�~�֭���{�O$���]4C�DK&"���o�8�����^SAjI�А�pZ� �v�I���A$��¹�����B>���*"Urh5E"I�o��2Aq}������4^jj�C�'\�<I�*�0��֡��t02�(lw����$���dV�X� �g�~��¹�b2xm1���k��7~<����~Y���a\�j lmp)���a��Z]�\��fY|~PЧ��三��Z`����m��VCq������~�a̬��~����3+U5�������9B��,�������'''k�5$��u�b��X��, M�M#,1��y�@#"M�/�:�~�;E�ɡ��+�~�ւ{=���zr�mQ#'=$�ee8�^�� �q?q�0���5gJ4��u�}'�&'�ϭ��O���C7_}�8;�<`rø(!4�T����/۾m��/��^��N�/:̊� ���E�d�3�酟I"�clׇϋ�pB�H���@|�.��UW]��G?��	0��z��UA����\�uۓw��L7�1�O�I�
N�T������"���F�677)��E����9\��\�Κx<�!�ąDd�6� ���}�mii���ތ��R�o9D[&6�.*�H~2�v\P�@�Y2
���� 	Ǟ�>Mӏ��Ԟ���=�u��K.�����}�k���Gxp�{�$�>��=22���>;�\Z,6¶k�?��o��D�� ��Q헂j<MN��Ǳ��	�2
�S��>�(���̜ 2eE�B^�($RA�{qϾ�������~���᭷��}h� :f{Z*\��2���~�T&������Q8vw�`.�VX���)9a|,�t�A�4��h�RI#�:�of�*�8�(rI�AI�K&N\򅐸fܖ40��x&H�Hٛe"�>�L<�ܜ�� ����f�=ONN��N��f#,�?���:f�f����wv6����jk���;��<y�c�>���� ��X6 '��@X�w2"��9J%��]��T�|&c5�}��>�v��W^y�it�����y��C���xb��;r�˶��`
%�s��\+F����$8a��o@�O��@RC4�aDN��/�m=����XGG�0Ea���"'JZ8�ӛ/i���(@�ٗ"W(���iHۃ}��	2��s��1�7l7��������普�,c��h%�ga��"�������E��nذ	�5��6K�,|����p�v��N���Ʌ�L~C ��7-�R�.u;�Fn	M��ؔk��=�D�F����d2�;�"���b��CrRA|���6��T����w��ܷϲ�o���m=���V_�}��MZ�$\�|<}�t 怶d2�iY��B�
�hn2���` 5t=Df8�Y)�5�;��P8 ��5Q�����3B����cҍ+ki�{�6�<�O��r����Vb�`��x��>o�w���~G�,�;��D����W���^�º�Ln<�L����7>�s�=���`m��G�.hb!GA����%�Y�yM\�W�X�)#WNE���@T:����M-߾��������g>�y�Xm����|���Ͼk`p`3L�5 PTl���*�t�QyR���0.4A�B�)�	�F�38awww*�/�+Zˤ�LH�e��t�����K�	��߬�C�Dl��"VHK���dz�4< �l�4�a��qh�0�?d� �CHd��V&���5��@�b�Gt��2�o��п��'�6��ˠ�6h�ѴE�BZ���g�>�8��h׏�Q�׀���s�����Y԰���|��;�ڝ@T~ﳟ��/�x���?�l�r��%����>���{�������a�4�ؽ�U�䬆ߺ���0�j0_�xT$e�V$b�6ҲT�T��׀�>g��$��lrn�M����ʐИG���\��!���'>�ccc��ƾ}������C/�_�M'�c���?ٸq���T���0.
��@�����߱c��w;~�����(4��{d�>��o_��'�L\FB�H Lx&�1x�{����u�W��t����}����S�y�'�ڿo�;����j���ׁ93�e��	�!^/�AD�����V<.�>08ac�5�4a�t`E�߅�@[[��r�Jo�� �r�Ey!�
��)��}(q�����"P(c.��������4�[�u�qP��`��@lN�B��X��Pcc�DWW�(�?s�wx�??�~���9��~����Y�J9m�z#P�7��Zc#���dَ�"-��\R��D���r�G�PW爿q<"�6}a�w}}}�����I�ɓ'����w= m��>�K^��)\��wMN�����lf#�f-��50~:��Qx�BDذmx8')��J/�$Ҏ� nKZR2��vd&��U�<��Y�9���>4�񜭭�J{{��	��̴?����@4G_~�̙�o?�`+<#��oh&��Ln�:����������zf׮���V~�S�MCQ9�m=�h��7��NJ�d�-p�J9(�`�9�j��V�X����7�j�`����~z���<��]gΞ�5MU�u9�������&89"!M�-�k��"�=OMM�A����j�@�,�������10O��ʹfH3�����q2�{B�0�ᖈ���f�n<.E�Ph:j �M^�%S�W��������L��@ ����m7��̲e��:;;���~�_Y����R�^���9@��с�����\�I/�B�50�.�~oT�RXUb���*�\��N!����^�U� 8D�lL��y�a���g~�{�n�����Goo�ck׮���8�B��V�=w�}������<z��'�V$�����%]������XՑP�?�[�8��]�ь .��8E҆��2ˢ�2�]���J���<>�i�%#�'�O>ADpP���$]���\�A;CE˺�,�~|�%�~8�Lp�{`r�x� ,FW�����o<���;a�[�M�4�B��nS�������&_N��b��I')%Mq`"A��S��>�����_���{ѯFQ>}��U�����G���G}�=�&���o�Dl��H�o��/���L�%�E61�:t�K�bu,l,�/����j粹D�2{���S���Ovtt����0����677#&SQ~�+*H���	$~�j|K�1��&�+x���%����|s��w���1��$�;�2P1�k	��Jc@���o���w,^���K/�tͅ
�e�g�A5�ޑ����{fg��Ύnr�F#���j_�p?tx����;��	��.h�%�/,���%
yJ�G>)^I��:���ݻw-=q������#t6~ɋ���!E���6�8q��n߽{w}��%���a��]Z���i��3��%�w=i��Y8OQk���a�gϞ��U�	j||Td!v�L�8h������Nh^D�[�]��𒊢6�LVH����٘�E_rj�4Q�"�Ҵ��e��<��"KU�׸�i�����`r�xU����6���;o۹��w���B�l4����+ȱ�B�q�D!?=Y�	��R��`��bw�dm����������{f^�0K$q}}��>����x~��w�.h@��]Q�rF,�t�@8�۰H@�Hz>5�dw�&X,�-xO�9��嶯^���+���Ѝ7�=|��[<���ct���S��Co��w
�Ɖ����)���W�����`�ľT��N�[�����a��p_�ֳjժ����:�y�f.0xp�}�a?���
�������L&uܫ��>��{]�&c*<���1����l���=.��k�D��&��ycDmii1`]w__�|��X�gϞ�Ë��k׮���fFo?�\�o߾�m۶�ٹsg��������ˀ8l��dECUsa�ha�%�d*Âd�J=�8F-jn(	:��k�m�����{���+�tR��!冓�Ĉ�wgg���`ppP�K&|�<;��8��'<>55��^���:��6�2`rø�����Ǐoٺu�=�����Ǽ�&M4��S�u�8��#-
X�p�<.i�ԨJ�Z�������`(�������{���:P0���j9r��o?�~��MЦV�d��L�+O�*��9J8��dB?����H{!�%u���@0r�Ȕl�D6�����]w��{�q�s��,��|��#Gn���B���'T�*"GЁ�5)ilh�|,,AHp�wO�<ݯ�MQ"r}'?,=��mvn����|�	�&a�c��3�h�Z�[����k����9>^x�	����<�H=
������[�/�����!�~�S#8^�P2*�@��(�q;|~�7u��E����7?��S�gϞm|��޷�=�?���1js��?���[w?y���+GG'�m���Լ�̦T*�1�R�E)�� �Q�y�po9�PDc��.T���7+۷�p�BzP����&f��5Y�N�D�0��59c��h��K���j����ͻw=��/ y{���/��j0`�ܽ{���v��SxH�[%3�E$��@�981��ON��T����y.Dx�p`�����[��|{Ӧ�{?��e���Sܲ����n{l�O�ɇ����=R4~.��x��LdĶ�;D$�uZ4�$G��������|>�:�Fv��6疷��%x����g�}杏<��]0�n��0V<N��h�w��7��H�|s~�zz�t�5��Ihb�qAj���L� �c%��X�Ϭa����@@}r��U�.���q4;=��C�?��?(�W@n���!����;���$�H�d���B��f��M���^=)��☡0gGh�A������1�������`�Ԃ ��������G��v�m�<y���+V���x$	�3�˃>���Ƕ���\c��H$�yzzr	l�"5���O�`�V�D�<.���]^?�Y��曕G}T<7nj
��CGmW3k��t�/���X:���퇆���1iH������p�[�ٱ�����+̝ۙ���`rø @����g�}��w���[K���s�������>�����N�(8]����J�.)�j �ɀ =
��_�x�#�ׯ>��U{�aҪ߹s�͏��?J&W �	������QU��h�l��q�E�/�m�h)���`��(�2�8�xc����^}��믟���ە��sO����zv׮�f��V�a�2-��c��=�̇�(���Y1�S~ ��\.<���ȑ:?�dxxX�ǭ��@[�p� 5G�[��P�����^w�u���rK�#�.n|����9��FN�1�J�P�����K��\�p�w%ό�����MA3U��q�`A��|�ϱ;FlQ���~�Ǥ����������׭[7�r^�w�!�4��/>�[�Ϳ��50�k`�j8��a�|.����sB��\Qz|N0���E�����g;���ry�]��O &�NZ/��y�O�F�h]��@�	��{g�:N��s����P�6����������\��h"�)�O��(8qR!�7Aݜ�(�ə&�����1Y�������K/}�3��{������;�u�Ooz������1���Z&�%�+��PP45�'�����oK$%����Ng禦'�k�ozh��O�ٟ�Y?&��җ�d8p`Ï��?8�{�6�p�=M�hB��4݄���"
$5^}�FU��D�:��p���z�F�ێ+�S����	G"bVu�۞�hݶ����k֬9�e˖�������k�r
>���GOmO��n�M��@g���Z 2m�qL��EV�8��1�G���ċ>��`��M ����OvQ�����n���ї�Y���+s}{�?��?����Bu-�Ԇ/\T����[o-�W��PpzV��u�;�-�^�l}�g��/m�`E�z|��޼�b�&��*��,�,�C��ل�<���
T2�D�r�������~������z��+O������޶m��w�:u���G��rCJ5ŝ�,�C��oBɀx�s^��p�C�A,R{hN4�D"��b�xɲ�߂7����w�j�oa���s��'��\�p�=YFSt�*�i�- 2�����Sq'KG-	��@��~p`�M��T*�ӕ������F���1�|ǎ�>��C:4t��0�FM�Rɇ����A�����N��j.��׸������n����Fu�7VLL
,���p�Ӗe>W[[�tGG����nt���`^����~���o��9����`��1t;Z �C��8��u��+)���*3�s��dI$�D�/S$,����������%�Q���w�%{H¾� �,*("h��n]�U����竾O[��Ӿ�V}Z7�pG��$l�@ �,���e2���|���&F[5H�{��3��n�s~߳}ϴ������}kj�>T�tk��ܴ����޽�����{�|FbT�4�s1Rm87� ��!%sh�07����}Ŝ˥�7J���pQ����<nI��^.I*�,#����z�x��F'�:"C�{"�`���>�𭷞�e�M�i)�΢�MN� j@^Z�����9�y�P��mf@�����ydco��`!e>���:a$��b��Cf���h4o���Z6{�읏>�h�[o�uFϹ�Q�|�'���I{��aTCC�	�N�P��؋�[#����J\pg�E�Ճsеh!�p#]ӕ��rS��o�]�o�>�O��,]��[��'y˗�v���,�r��wwp�D����9<���:(\��7���#D�牓��	).t��'�J�O�8��N6l��c�� s���;�&疼��Ε+WJOO/��/� `~�.��d2����h���5��8!N�]�E�������В�G��w���bSee�"�t{�9�I����u��5���?H:3H/�P��a�X7�^]]� 6��%��NB�'����G{�L8M%�����PDk����p퐶B͒��\�N2��B��n4�f9|�������X��t�h�������1�7'ߙy��ݤ���I�W!��#d{�@F��hXM�e��|d@+ɸl���~��(�3g����TԲ�K��8p�7~�o���l��!�&����
�0L<�݊�y�Cd��d,���Ř1c�<���'xV�b������ɹ���xz������\�J`�E��"c5�2xd ����u`3F�GE�)���\�i{)t�_�)���~�0u�T�VOsn���\�hѢ�G��).>6����I��t�b�f#�Wt�h3/D����1�q�!����U��_��w_�?p�������_(((8��Ɲ�2��z�����ޫ)..�t����3�1�����Y�y��
	�p�رc�7���3��ù3�AdVf7��h���:�����L���5�V�������/~]8џ"�Ѥ[�2�3g���������$�)�<��M�}ra�QN;E)�,�Pj�>�������3l�~�:�x�ȑ�?饗ʖ,�qG't%Gi�b6;Sw>n6F�1�`�0��T���#<3|穄�.�����^�,X�`;��fx����jժ��=zy�	��q�
wz�0	 $��``a���������6��FEf� ������1^���@���z�acRR��C�)&��
@��Ӝ_��x�ת�:��X�s��r���K���n�a�G�'G/h���_/9�-BؑQ���ȈD9>l��_��~nnn����ۺ�<0�L j�|P���I*�E�;�z��P8~�RU<��I0��� gaҤI�9�B:)�=�2f����[�.ꕘ�'M
�����z��=�|V����X�5:Y4p�I�	
�w��q�ƍ�-+?9�:J
�t��-��/bj/:%z��9�W�Px 08 (F	���r�����~�Us�~��8ܜ�S��G���.�ؗ~��l�	���S�x�t�96r=:KRMU���q��MMud趑a{������裏��UDl� �~�w...�M/Dq63�22m�~\#í�����U�N��7'22:<�R0+s��ԓ<G*����-��	;i��:th;��3�!�I�ܣ+W�<J ����������t]F 9���ݠf4�Â��;�D�t�5<n���ʠK8FQ�#ה��Y�x�	sZZZ*��O�y 2D � ��K���o!}��t.�g��  4�� ϋ��9�#���7��\ ]t�E�iCG!"���.Q�>��@w9���b��E��S�_�j���E��A��������uWй ���\R���k�^���/������t��$U�aÑ<��4�H{T����g�� (�"f�\�U^y�]�� 5������3�>Y�Ɍ�{����42P.��9K<�����|[�;&��1��}m��$_z饟�v�m%J���gس'e���[������kL}m���M��+�p�p����k�a���	�P�Px�Ũ��*Dǈ)�M ݣ�n���L�8���c��!j��^�$���������I�o��g�[&0�rWrRw���kԙ ���&ɣ{Žq����=��׿����_l�馛��<�{	��Cv8p���ҝ�UEz�gfaA�L
�3����2C� ;B:#͚5KZ�~��tR'��O�Ց�Ck�!��6��������l���z}��}ߖ���	0.���H�h�F�$H��9�I�[�������F��f�GΝ����F@o�4PN��ؘ��P9D�Ŕ�}��m���I��!����{MOYP�zژ���͛7��t���*w%��9q�7�[έ[���������w[YYy.m��;��W^yűj�*��̻w���k%�=���,��gc�]N���́}4L�PC��IH����fcӊ�����ѿU1=o"P�qҤIG���?5-[�L"Z�D�� ��׼�{�2+++����^���jO��7ʐH����!��O(�6@OP��� t8���+/�/^�x�/~��q 8Gi�/�۷�V[[v��=s�@��D$
�
��P�����#p4�&]r�%�p(�z��"�{�E�G���
u��ɺ
�=A�9p  �3��I��=� ׏��>���5A�tڴi��\6�h�wȺ�n=t��=͎������U*�Ɉ���1�KD��ୁ���q�F�q�Jk-���Y�H�?�����Ν;ǬZ����?}0��<̑O �����A�Έ����g:�wx��/}����@����<m�򥏻=��hv���	��lq�q0�̝���X�gcm�0�8|�n����6Q���������o��^cD���%-ҴiӦ/�ޭ+**��l6�9��_�\��ȄA f�ffc�� �ʌ�� Vf��$�?�hћ��_~y�c�=vZ"8��SRRJH��LOO�q�D
HU��W�Vؗ�Og]Gz
� �����R3{8t��i� q-����N�tcx
9"���Q5Օ�Hޞ|T�O:oi4p���Dl�{�zͺ�e8p-�}��Wͅ��	R8�7&6^���v*E����^o���˩&�^C���9s�EK��C)����o���7�{���A���.��&�#�C����#�cH�,H�����6�Z���Of����?�ڵ�M���W�hni���a�i��S�!\��'�bJ��Y���o�y��4ܭ�]+Hп�_�����6[Ē!C���E�=	Xjr�f��K��'�=~���Cn���t�]H�ot(�����4�eܛL=��IɎ��o8��`��իW�/^���{�<u&H�gdd�c|)--��;�xIm�2{�.<_�f�<<|}cB���Li����ԩS�)((�����J�'�9�>�A���\b�m�<��H���� SJ�J�o�>�f��-����;<�����+V�x����g��q ;^a���#F�V�����E�.��~+�,�V(�R�ቈ���x5y8]r�%�ꚓ� ���ѫV����|=(�1]�2�H��
�1���"^x^����F�m�^������u�-]�����Y��������'3+F���}!� �}����d�>G'�������$�䎎��1��cc��ϛ7�xg���&�G�Tr�ʕ+�o��%��U������8��C�y0��)�h"�0H� 	
���ut?u�<�~뭷,��>�O��#�C �8���w}_G��.P��S��x��27�ǎH5 � �	�/L��Թ@Nm�c���F�S��pm��0��ZWW77==����B��t�n4�Β��5�<�_�B{skK<�����F�����B�9\�E�̤�M��[&�S��������=eʬ����=��u6o����ܜ��uF}�vO�!���
fVw`��>l2���C]��H �������%y������0�@�}!ua򶭿kin��p<���]�r�����D�v*�T7J�0>
�U��K�~���-.*�]����wY,�h�袋z�����e8�v��Y[RRZA���� Z��X������9�8t
i*�b���)B�,�z�������|��g?AM��8v�%]z7'''���U�����Gz�"������v�����&��"B
Gd���Ҙ1c��k~�FGtM*΋L\�G�8�-R���n�<��O6%�H�v�=9T:�9����iiiU�^���Z��L4p�ɿ-���ݻ�/��?~�.R�p䂽���=RPD	��\8��������� )3y�_��D�1eʔ#�>���xD�I G�=u��m��Gا;�.�H���6P��0��f^
6XHE9����6]<��Y�n]i�"i��6o�|��W�����t=M�T�gCn���%<=�t��n�)��J�����uDD�����O����O�t:��qq�����+�@�&�S�Q��<�̫������t��]J6"���q��yee�Xԑ�B۴��a���l5�����1�%�����~��SO��� '77w�믿BA����h���[.6��B'1v�9�d�.�8/H��ѣ�$qڦ����\�&�w�b�J��+�Q��-D�aW������@O�PWW�����K�����:� �n4���f߾}�h������VR�8r���B@xF=f�xã���K�mR}#fD���Dl��勎�,�Xl����{�M7ݔ��=M����mܼ�gn��R��h�`�APF.�V���>����DE�GSSS][[����|}͚5':a����'OY�l��t-��6��P*��?�S"60|xpk)�OU��ǿ�(86ۤ�I}�w�;��ғuV�egTd�'�F����O;u7�&?��i|����geeU���0�{W�#�M\��a���a!�=��N�m�b$����`��o���FZ�?@4�t��(�MKK�x����*��m���`�đk�(�_&�3�(Nd�Y��=�mx瀨�R� ,���P��Qf���a�?\�l������U�۷���+A��u���Տ��]䔖*C6{�}=��M�-IMM�jժ��븇��wMM�ކ/�g�-!0LPZ���2'����U����썉�9j���;|��5���OU�z(o
���~��9L��X-����sF
�;�8�#��`xV��_"���X߰���S�}��G�2�){RF|���� `s�i�6�#F? ���:�(��� ���O�~�XN�<���f�-�ק�'s���G�@#����t@.Z�h��\t_z	\�cP��{�UN��^G���ڐ2�I�̈́i��<�t�͛7���><-m� ��/�.]�������(F���&tQ��z"�#�ؙ��ћ��.�ƍ'edd��8�a� 9��ʀH'��T��ItP�z�Qr���}ˤ�nL[����������t��n4�VA$!%%eyD�����Io���q���H3��4�&%&��b�ee�2.$Z�#""�v{D�Ao��x��)�������Yꉂ:���_4�����DEEklv�Y���GtEq:J<zQL�a�`�LFScEE�q/xzÆe]Dl�������r߀����S�+ߓkl����2��\@�8���&�I�Y���"�{̠�<b��%/��t����L
:�X�'{�?Ũá�}` �3p�Gr�_��#p����v�o�^���>��s�o���G9-E� |饗��۳?TUS�_tl������b���A$�i�g 6 �E|��I����Cq>�5�⼡�4f���r��R���`��>c��/h1M�7oO�^[TT����Û��@4p��7
\2c��
��w���xRZ����,)��e��D��f5O���FD��n�@�""�k�S���^w�չh�z�����Kٱ�&��4��]��y���#�8�"�Z����0:m��iN�pѦM�ʺd����{�759�q��q��1�h�p~���6h<�^"<HDl�E���xv�m��/�`\�O>Y��>#i�ə7��+W<x�]Z��j��1b4�8H�`a���(�x}��\l� �#`�U}H||�}K�.<��s=���e1��_[������t��<9:���6f�L)�u]�q)���`zРA~�SWccS�P�6��� I�~[[K8������.�V��"���$�;�vpFu}LAaт�;w��o�}�h����M�Ю۲n�͛nw����{���B���C�S�h����f����B�k���:��X�,6Db���Q'H���?pŬY#`ӣ�WKJJ����A`���=��]g1Y	��$tI��^�^��t��>�U3�8Qtp�Ё������6eee�.|�Ϊ�����xxiF�^�!�*-�v�Ԭt~��2���y���a��.�F�I�~%GSS������uWlt��]vI�/���P��/
�qٟ����;���M������x|9�"�Dd�����D��J:]� 
��[���o��b�59g�\�ᡇ�v��4:s�#�<��%�u��j��H�	@�l	���!"2�� =�U8$�NvN���#F;~��!{��m�R1t���-��~d�*�h�t��(�76���
�%E��O�)3��N��~7";7��/S�D��Q�9>>E7�|M��Z�v��5�V���q�DJ�!B�A8���Lt���m����a!�
傗b2YB�U�,f�q�G���?�����A�꣏>SXXt�d�ȧ��&���t�|�c��U�WW�$&�y���������)�>���kJJ
�}@d�`B@�X@p(�x�k�r�x�BCxo<
^y�YdL?����Ob>�sڠir��bʞ��Eii�'{?QWW7��79�:,����C�yK�̥Czz�?&ze�X~�|�r0�9L� +W��&�����Q��Ek���A����n�3��; e�������'7nLJQQ���֖+�V�4��߃@�9J�r��TVg l�x��e����\_�p��#�����4�$����&�O��t�5��x�?%O!Z~_	s�Q����rG [p4`�G�pCC������}�pYz����ç|��O4?��RO������۷_���`0�-j�P6X�I�m�0&0��.d��>\I�n�����UW,�����O&��K�?������Ձ��y>w` 0��qN��+�u���3ν��Ȫ$C��o��K�O�^L�J6��xA��K/��qǎ]Q��1�q:�&���f,�p�����J1b� �Xđ��d��=����# Ҍ��J+z�
�N�6m:��~J�:�l�`:N=�� �_#���>B������L�e襗�X6mڴ�nM�,((����T������]\�V�	{��)Do��.,|<H�ͻ)==� ��幜����&aA�bɧKF�n����Ʀd@0GE����u�QoO�56���9�R�FFF$���i��~����l ����Et>���Xn�T���Y:<g��w��!��A��n�aI�YQ�>t�vm�n͚G�:i��6�&���v���yz�-��ǝX�
�0�0�d�t,�X1y�ď�z�J�V8��Y$�?���t��{}>�c���B���="R�@�<<ӎ�hZ�{S�����H g��`ޞ?~kNNΖݻ�ƶ��>@o�"P�c�M�0��pD�q�v����kjj.8v���I�.����_�z��̝;w�)͢�Ɠ2pd�Et��a�
��l�>c0D�1��#���٩ʒ����C����6�)��DRQ�~�d��/�z����V2$Q�8딉��'�%<�^�<�9l������8d�[��;w���4�_Ijjj�������r�zt?q1#��V)���;��k�%��w�ԩ��z�o����������t�_�Wz���eZ���X�e��'%��ʧ��X2Z4Q�D���� ���/��!�u�s��D�D�o8K�.]�q��Hҋ��H0���)\ၒ��a����Zѭ���!Za���"��}��ǯ����3gN��#�y���������	L��@N�2.�	<� G��xF=]YYY,���źsܸ!�-Z����Z��ӟ���-�SEzo���`'İa���l) %�>��W
�ʹ�+�g�b�w򻕕���A:�&�k�FEX�dɨ�۶<�hi�)��>(	3�rĆ������;>��g')�26�M�2%�l6h���_�
Cx�w�#�g�Q&�bb���'\:� �����K���̮H	Q�L�{NUU2K�K�|8�&_w�/����P��y�!2l���,Z^�=��-��w_3-�&���B:��t:�<�9������ɶx�� 8� tP���ۦ�Z+��euuuͯ��z�2P��Ӵ7�0�������Ҳ�t|*����`���K tFṢ��oll�u�w�>JǘO?9>r�7�/��Xvv���|�����j��5>�.�&L��58���5�m��~b2�"�


v�9�JQi��<���;�u���555�HJ� �H�[a��O�M(�<�V�<.9��VD6�2A��d����~��e�C=tVy6lH��Ͽ	Ž~�F6DzQw�-�\��M��
��F�N,X����>�ӊK�gd�����Vg���t��n �l�h���9���|6---^��ބ���f͚�� e+=$M49�:ER�z��w>��� 9��hlt�"#�t�\���������j��߱�����b����?O�-��t-�/^��ܼe�P������)\DlBz�Q��%��6SQQ�����\r�����Z�Y%���~��rӦ�w�h��0�V�t��'��]b`o{�S�������G��w���%��,V]s�#�����������RG7� �|���#�����֖[規�"���7 ��q8�.�V&�#� D�����ܹs��t�΂�ʢE�.#�q	#;s���m�~�;2��J�������7bĈ�O?�tCW����X��.��T�g� I�|���`L:ޯh��yZ0>�T`���SOCC�~E�^q��۵VoM�%Q N����m����rذaqz�0@�-$��%��a�ŷ2OL���!݊����R���Ͽ��v7�!@�D`�3�����.,�]����9^s�Ϡ����w�ر��"�RRR��ET�~�:v�ȼ�>�"3?�诓��FTWWZ1w�Ng�N M�k��}`��)��]�!C�ܴi����dw�+58�9����!�S��kw:o�x�����e%�S��x�EĀA�У3JQ�QRdDd��lNILLx��;��O�Yl G��_XXx5�~����ɢ|�}Gk*�&w3�w+�Ȭ��o�ו�xz���	�� �,�
N�l�"�%w_E8Y�r�ڝ�pQQ��V��P��t�E�&MЀ�&�(�2e��a��$z^@ ?��L�$ױ��S��Y�9�`����"1..涵k�@�u	����ǚ��[Z^^����'�9����=���ı�p�^�q�JQ�����rX~z���C��je����ڷo�ҷ�Z��������UUU�8g�R��b�3���̬n	���5x����I�+�oߎ���2΅�n�CA�iÆ�6lX��vg�]�}1���+*(����P�%5�tll�n�;,6�椤���ϟ�l6(�{�?�"�6��
C�6��-��(x�4B��������o�}�5�\��b��W^y�'O��f�"��G����6y
�&���\���8���C#��#ÞI����ٳAT�M�Y��NzP������ԭm��N�?B��&A_��XD-`����͒���v��''⁵k�֮\�rMwwPa����˷/[�b*���	�D3+1�������������ݮh����=)))k�̙��۾�KZ<-���OJw���9<���Fd����6���*�\*��l�;���#���]�vY�wo�-K%�M:�E7� �$'''nݺ���ʊ��!oZ<�����F�҅��4jk�ĭ�PDzEEG��c�һw����sO��i�|�Y(�!���˻�N�������VJR���[��p�~2C�]��/Խ����k�����֭�w�Q�p8JgS�Р@[�#rc��p�{�\.�X9L҇龴��yg���O�&��4Q"8��z��m�R�I�n��#8��E�
�fx��h!�i�pf������{?���]����;*����gg�^H�y	"�<2�TjJs�3c�!�b0ѝ<Y�7::�#G����S@i+))��ݶm��l�U�vF-�����Bz���85�d0�&�����VK�~��ÙV�o��o8�ST�9�����1�7o��ĉ�X,�>mm-z9b�S�-/2a\0�z�^��@��ѭ�yl:t؛W_=7�l6������I��5��0����5��C�T�c��PL�~y������Q�IZ?�x�\��8��K�u�`�+Q1c����tp���Q~�� ����+&���O�S�O>)i��� J'���Ez�~\cs1�h"�=��."�nx`%�q"B���t195w�Z����Yԝ�7(�ݹs�����m����q|�#�}�PnNP:��c��������Ǐ��w��"	y7� xTVV��o�k֬�����Ц�وmpg%l93�C8O�F\3t�6��������<��lk!���l8�9�7����o����/R�1(h�vP~p��O��	�<b�\\+�����6�M#F�6���������?������5�K�@/�p��9\T��\���!�Ȑ5jԦ��s��6���D2PwGG���_�.�A_D��)G�07��@f��&�r85�--�:}U��4��|D.SRR��.�_NNN�tdnDD��G��S�)\��V��r�W�"�sӾ}��}�YR�u�q^~��u.�d����f�Sc���^����˺���� ��loק��紐w�>�����v��f�ƍ�C � �������evԸDy@+A�)>��������7��9�"��9O$--ͶnݺY����n�Q�h�y%���͞�!j��Q����נ�64`��^{Vt��A
<%
ڸ+�I�`s�SLg����Nץ�~���?�yNW�d���l�tmLL�4F�����5G�7�'"6^���0�����B�f}CÆ>I	K�L�R&i��y*�;YYY�P�)..N�E|�	�%����z���xQ��z�]���͛7�lڴi}wwy^��'��r4:��~����3��Y2�!��ب�7JM����v*�笕+W�uE/1p�@���
�������Z��;�pd`����5��9���ѣa��>3�홒�y�w�g@��~��H4ps�./��´������@��k��ߡE�yV���� L�X`{��o<x�����/sǏ�y<��̃�ɦ��z.���3ө��X6����h:6u�����sO�����a۸����ON�k���{4�6`l<��>�D�N�H��\����j��nOccCfLT�b��a����&�L�4���);����N�8��V����1C=� 6 j�c2��#��(��{^}��└�#��!���'����YSS��h���n��#:���0�a;̅���f$���������6W��>Pd�x��G��K�|&���-N�q������v�����
�e����l���g�#�qq�%��=CugO�J7�@�Iag�M�)���Z�c�T�e��ψ^f$��0)}�K��K���;�#���YYc�|�kkk��s�Ŭ���燴Vs�R|��B���g�>�U�~�Ν}���C�t,S�-1��=!u��_\��F��I�A������s����hr6�M7�q,[�l��؆���Io���ŉq�>îa��ar?�Y�{$�s�566�bݺu�����y��G�rb��#�����INg�P�@ E��:2Y8҂c���ȅ��ʮLKK[	����A��)S��JOO;]Wx��3p�SR��+Yl��:p�Z0@:t�������Ԕm4�t�TVV��-D�9������z8���Ζ��0[�b)
Wi-���2Yō�!]|�硐��������7�|󑳵xX-��y�WF���q��Fׁ����]8O�r�L��v�����1bϣ�>��b��|��2�q16s�0�"8C����Au>`�\1��IQ�vp�T�#���Ƥ=��l4�D-w�ygCmm�jZ���^�K�ͣ�455�g<0�]�p.�F�Yqhb	L\�����r�ʪ�l�6M�ۺu�c�������1�6�����"��e���h�kp�-�z�񺱱�W]]�,r�R�'��ǐ!C<��r�Nr�����01��,��-�Qo��=]����������a�!���lCKkی�_%��Kٰ�y�z�h��,ܫW�N��ʼ���a�Q/E�d�0#��tx ��[�3Q�J�-&���7ܰ�<��Mjjj�Ņ������5�n&�=]jH��>o�u��(���/�������)..�G�d0��i@��Ɖk{Х��������p��S�ֈ����pLM�QX������}P\\<���̎��4�� Z���7�) � Z�T1�>���?>@�����SW^ye]jj�g洷���PDnB!}��t�\��E��Ld��VT�����R�U�נ���h͚5[233/�s�m0�tu��%��CR�S�gpq���-�'G�u��F���ڳ�m�՜���-�9GeÆ�Rw��_]Y�@��K2��:L�Fk7/�b!Wڏ97��2p�}\\\�^�GEE�=o޼�H�Ι�5�XV�ɲ���<#�혊�rNZ�,,�U��7�q1�2���%a߯��E:��
2 6NgA8�1����.,N�� +�}dp�����W^9�P���D��E��&0�2��8��<��̈́h����4@��@�9mC�[I�..))��?��?_��� JiiiG�����qj���ҩIR�]S�GT]���u�KJJg�����]�E����W���lI��h�0��\&�1��#;X����jmn���m؎TXX(�黸n��!�)/��i��]t��t����sP���ڵזWT�M�G�N���X��x����G��n_q뭷~:w��&���^~��.�k��n31�2��031禙��p�]�+����
l�Z�*�ر�kl6K�@@&�b~	��䨍����ڀ$��f-}��/�����h�ɷ"�v�J_�bŲ���D�c�A�����s
0�YRs�D����j�N�W�W[���f̘�X�~}
��+h���8�Q�@���,���������C�o 7�ٳgW���JKK��y'�q���0X���r�J��"k�����sd�k0c��b���nZ���666�=��[�S4ps�	�}�ᇗ�?F�MiT/�L'��A)�U�z��+��!R�z����+?$`S���a��"555֢��)�!�������?�B�p����)�F�Q�{֬Yd�:l�6�=��ј�r��lH؀����a#�)*tF%$$�WI�l���w��]�c�=&i��&�.�]v���ɓ_lܸq ٯ���"����dn,�X�9�p9r��5��`�׷�]��8�����l۶-���h/�w��h����C�>�;3�+�B�l0���v�0�]�222��4s��y晔E�]K6Ð�؇�i������x�}�9T��)���8�J�E�r��'�99����lcOm���9$H��b;�x��_����tC�pCC�ƃ#\,�sH�ȭ��P�)�蛮��wo�����=�),,����O�i��\7�cB`NM�g��,V_��/'�nWW�������yא�	�<��k����� S&�������I�&�K�RMN�(�7���Ջ:4� �,r�,H���Z�H�"�T���$�&��8}T�]�G�b�f����9d'�q͋z��zj8w�"Ov:���~Nrr�:�[�&�g�>�|��}n�w,ِ(�>���^_����4�4h� )77W|��T)�|]#�s�IL�G�M:���E�5psɇ��7=}�/�~�,�Ym�@��
�M���I��c� )��P��ɓ'�����,_�F{���>����mζ��NĨ��Ϩ��1<n�kf�{>�?p|���M�}m��ӟ�47;."�bUS�s�����kl��@'}�uܸq��w��3�&�h���E󉆆�%EEE�i�T4����K�����>�<�U�ݑ��W�ٳg�M��t����~��ɓ�>�w���`�;Bl7�قp�����2���d��P���o��C�qL�2%o���utQlÔ�Kxہ �^D��Bc�ְ��YpޘMV)�IA�B�Q
Z$�}e0��t:���;v�2!6�AǛ��0ܜ#�Ψ-[����o"��u�yQ�5��@4��5��Q��BO3f�K���-�CL���#�@�^�G��]2��aO�'�*�8!�v�@ x�������>t(�J2�c1��W��R�9��t��	����|�*7����iQM4�΂��d�jllAz�+z�3���
�ar?ϥBD��7�^"]�s�ʕ����nq�Ⱦ6�����K��C�FǠ��³�����T][;'r�����xg̘�?%eG��P�"3��}��_%�[��a  Q���>�hB�Z�S�4����U=ٮ�f��$�9d׮q_|��������M�$��1��p0$�ył-��y=�����fV
Y}�y��ѣ߼��v8�ǅ�C�c��?J Ĕ��ʼ6P\\N�A87�t�t����z��A�]�������ݻw�H!�ǠRM���ۗST:)>>A��։@Q=�u���UM�7��kj���?%�F6���x3k�z����ő�S��M			��ݻ�ڿ�����n��B�yIQQ.ٕ^��`�
�a0��L ��-�-��͎���߿��/�+�v###�8))1���\[�VTD���ͼ[��#�(�#{ń~�����h4q�9%=���յ��toINN������@[��CD7g����80����.�Y���s�;����.Q@�v���'�҂짿O�;$})ϲ9"�E***z�ݞ�t],jo��0�p����?pr䘑��ے;|������3�=��(�z0D��Ww>t�@H$^��"	�W���������4�D��'X�sssJKK?~|*��HL�{1@",(ԭ��O��y���{�k���؆V����5��G�ԩ�5%E�:���lҷ��G�������ң�h��fs]p�Ĭ�;w:n�)vu�m�z:9�C�k����H����X�'Jf}kKˀ�����m�VA�:�M�����XP����Ϗ�9�����y-�&�M��oU�}�"�@Hr���L)�^u&&&�ehϟ?�СC�9,Ǌ�%�=�����Ev::�z��/� ���=�ZJKK���ƣ;At_q��ۄ;�������:�/���&�t�`��ꫯ����-�?����I,М.�9K<z"w1	�i"�\]]��_��W���N}wץ�^�ܺukZccõ���Z[[��4���h
K�I� ���'@Է��lҺu뾢O�����x㍌]�v�ѹ���3p�;l�`�Fn����f�s���O�2��Ki)�.�_��769������6�Rmg_O�]�9K̛�V/���� �x���v�����H�_CQ�^_�X�*�<HY�bcc�_s�5�v�p�kRZR�DJܛ�X߹�)$�:x5b��Ń4d
�ht �C�������h�L���p�K�N���R�����;�t��'%��y�7���&�������@ɚ={��![w3�E;��0q&wEvvp~|����皌��+W�L��) ��������$`3ɀne��^��<�O}��)<�vg�EG��#}��L�<��lK���F��ƶ���;wq�z�nq�.$�_�F��t����(���v�ڟ�q2��`��:��n�RټysTڮ��8��見@j���!"B��Q����f��J�V%@����{�����ѣ'�K�j��H:)V�Q܊0���SG������ut�:�����,��9S�fS?@z;t<�[��߂;�`H���9��@�ԩKε5M49�2�������eee���ӯ�=������J� g =~�v��\���;l�ԩS����Uf]C���/����hV�Ų	u�M^.��K^����/:^pS�M۟9sf���C�dee_J�aS��������V�0�VEEEx<�

Vg�����t�O߱=�@��iӦ����9u6�;�]]UU���b4�uPJ�t]�t�����*�B��3�E�K#xi����ÂJ���ēO��+fA�K�YW��g����7��ݻ�R��TRrl`mm��^�"a�������:�S����^"�K����8������o�F�QM4���	����v|��G�l6[����3�L���!����b4�UYYY����r��^�����:t���
�Go�0턪���oG]S	U�USh=80g�wW�'��{���>���UKۍ���9����Q���6�����D���.1�YOσ
�>пO����g��V7g���o�1��X�Ct����?&z�{��F%�������-��x����DF�9|��^��;O"���g{[\��dz����";C��k��rR�O�1��_�I_M���n�ε<�fN#�KF�MX���	S�%M4���ddd���ΞM�z)�xc$f/��h 0h�� ���nݺ�>����[�u�ֲ��9t�i�65�9�N�@����:1�(%	�o��̙�~��G����~�_��I�.W�(�VApm�6�����"�h�8��.����9ٷ�5*��a���!�9�$�L��<x���}z0�B�-�b��L){ ȏڬ���l�`�Ȩ������͛�%11��p8F��K
hPw	�9:�1��F�F���oC���Zyy��ȑ���#�E�k͆Hކ�k�6�9D��	UWW7�L��a�.Ң6�hr�D^�_RR������0�:�Ŵ��_8���SY���/��ͽ��?,���������Eo��0��G]G���UM&����c��s �^�]�(}K��ȑ���VK��뛁�@��S���M �_�F�d~�'�}A� 6�#xp���#��}�������

Vb�tD7g������ص�ζ��{B_�_A�V�M�M ʗ����Qm�N��!C)2�.%&��Vk��d�|��׾9~��;��tHEE��h0ĹB!�h@�G�s��ੈ
��~��>�\@��?~<������b/�=-5q"҂�u���G��-����`[[K�)S̘1��M49_d�̙��k�nY�fͅv{��6��I0��E��EJ:��Q�C=-򽣢�w�\�r7}v���`�����U�,渶�&l��;b�c��6��Kz�]���׭7���a���V�7�`�Ęcƌ>�o߾�?6��(��a�tAeLN0�".f���b��%>KJJ?�d4�E6@��iv{$�� �6;$��&h-�=!��]7����ov�ޝM�(�Ld4ps��l:4���|-���D��#ء�'�B�7Uܬ�h�ǎ+��r1?J�455E��\v��`�t�S�tSR��:9<,R~4�C�#y&1�g���Ԡ�sڋ��
M�����1bD�Nk��D��.'N,����XZZvill�h&��p��\g�7�*��G74�^�dɒR��S��2v��ʴ��c�om����ڜzt�5O6mxyy9��.�8̆^I�G3mC�4GG���0e�]��ۨ<DM��~|���b�p�]t����n�L�F��T�A��2���M�+<~ۦ�TtN���S�9���{�Oޱ�;�����esب5��F�N }%&&��	&|2u��#��B
@�瞋B�Zo4ʍ�B:}'p#�g���A�:����?:��{aZ.�ɹ�X]�ǹm5S4�6 �d��cbb�Ǎwޤ5��L�СC�k׮�W_߰�t{�G�*J�w�����C��t=��p\�y��Tz���ތ=��l@���r�	����br͋.̬�twEXR\\!}3��9��Χ�#A�.VVwMu��X�5A�"7>oG^0D��I6z�!�&���#�kj�g������?vzJ7g�l۶-)3����--�覉ө�(���\6�!���
.�/�BZ2x���7�pC��@�-bp�Zc�7�'}��^2Y�����~�����ϟNK�����󻀔���_j��D~jpP������!C�d0���5�D�O,XP��_�i~~��������zt;��p^�9"΅� ?��&���+>��ҷ��;B��ݯ_�|�'մ�X5�D� qM�Rd$�3���Mu�0�!@@��lN)mw*m��vH��uF�3��!��ac�I&(H|aGݺ��LZ�>�؊ʊ���ec�z��#�nz����W�Z>�����������!|��2�sf�D8�W�^��]O���x�[�S`#�۝��^g�ώ!_�׼Uۤ?22�V�"o�R[[3�b�Z�À;
�3�n�{0 8��<'	t����h�	�ݻw-**�I`e�7� J�[��p��/����7����򌌌��w�<� 98����דy���:|�Sڛ �<��h�~��{���u�����G����:�Z#9z�up�k!G��J�Z��K�-�k�58�z�\��˵;N��B�pqvV�씒��9C��h�nz��ڵmĉ'�p{ܣAo��S̨�=��yp3"�A��tCo�ꪫ��7�I:ODSd"I��J�����f B�z���WUU���2`� #���I�xm:w;p.����HF�E��1bD��}5�D��'�^zi]rr����ȶ�G�0;�������VYZ�Lp���1)))s���!�.�~��5���#�p��Vȩ�S��
::����K]:H�M\\\�ɓ�>L�gL���q2��kMLL��D��1����'<U|��5Z���[QQyˉ���y���i��_|�e˦��|U����:(GDT!x�>a`�ya���G gߔ)S޺�kr��� ��������:Y�ôr�W�.
�Rd��9c�A���k}�`�Eg�ɤ`�:(�q����ZZ��ccc3Ə�8i��&�_@r�iӦ�������������=�7�"��ߒ�cbb�477_�cǎ�����9����QGNOe{�ˇ9P�O��(p����<���j�*�7m�l��\pθa���4zGч�)$���[�v2�|~�=����' �!���*��/Y�)��\N�����z����i��ҏ �顂t���˧544\K7o�$�A%��&��;�/� 7|#*|6z.:t�26�g�-�'HMM
��Շ�T����6F�>�A�����N�,�C�>J��n���1��L��{-�r�j�$M4�������8�%��|��a��H���BO9��if5��W��霺k׮��~�iy����Z,�&ڟ��!��mɩF�+�7hd��ۛ����CF#]ȸq�|���մ�6r�v[$�,w�Ju��A�Gͦ�악�M�s��n_��`M��Sו���ښ�9�D����E7=P �_~��ѕ�e�3����(�d0J~�|C��+党s�HE����fl����p�Wn�ӧ�nW<�^��P�'�~��\/�.��{�7G�>5��WVV�X,f;�6 ����hJ�V���c�D���O�,1bD�L�DM����{6n�x����>��}I�m'�cԴ�h0А�qD�����ʙK�,c����			ި��F���$��̯�H2wK�}�(��H@�?�0wAd�g�i�Z-(K���U�2�#B��ڂ��/Dv�:!!1�~7�l�DF�:����}��3y%�N/�
8v���@������+��كYX��3T7=P0������ֶ�馵�[��(����H�(�MJ��Q)s���h�ԩg|BkO��@A^�#�(�"K-+�)/F����ao���P�p8b轈S���Rs4��ŕ�<d�������D��$�{�n�ׯߺ��������3����T[8Gr����i�@_+���@�!���RQQ��h0O���j0QHA�mmm	�o�>����C��T4�M¶��^�������=��<A6q���4 ���7���q��ksp�=]kkk��b����#��{駻DB7=L�����P]]}yIts���=u{��t�pwP2n�>}���袋>�0aB�N��	��v.$��k�>��	RP���!���lht4ƙ�V��n#����ſr�z�ۃ'$%��f��kwTTT��!C�pM49�2m�4ߊ+����e�N�%�`AJ�if.�U`��DM�0�]���=��S�}S.dǃ���.`v���2:�}����59����-B@�C�i���5�ыsUt��ĸ�Y�f76�]�rY�{�nr��¦!��8$jo���� }��K����v���e�#z�+���nz���O��[\r��x���Ʈ
�:�`�0bNQDDD��n_5gΜ��k��7	����N�ЬZ�p�.�؅���&���yR�-ʨ����kmxМ��))�D��h%�������"S�D��(�:A64������Ⱦ��:�a��ε)Dy��jii�d�i����|$'�o�G5����NMȩ���Tʃ���jnn6I�"�T�9+�"7�ו��S>׹�.Ck��|�ݷ�=zt�kٮ9���ݹu7��q���H�p����k?=|��f�M��4�e��M̎�9p��&G㵾�?���;/�r�/L,�����u{�ϟ�����q���(d�B��|�ý]	+�𢤐��LX_PX����QЧ�m��{�:-��� �Ж���7n�n4��ˌ3<��طo_>��>��cD���H���� �|��G��s���{��@DD��h4���Cݐ��=D��2
�lhh�ִ7ĕQ��wRR�ȶ�y<^��	dee<y�d5�A�Q��i)��`HDjP{�7�$#�G]���q��#08�XQѼݻw��.N5�nz� :��/�w��,�z}}� U��U��L��~��lF
Fo&L����ѣK$M:Hbb"�}t�Bjr���S�O����t��ƃ������;�� (��ٓa��<��)66����D�3,���ٳ�����Y����I�uͣ�pM�Rw��r#�?>2%%���r�(4��䢧ց������^Z3�܀z��۱L��M���b�B#$���O�2}{yy���T'���3�Bʺ�v�d���"�fyp���.��h�<�X�V�^�����M�իW�)(,����^���d�jܸ��d~O�pX(z�SD��>}�|2o޼�Z:��BJ"��NM}CHV|��V�3aKs[[�NU��hz��:��أS�����;�ѿ]S\\�kZM�&�� �9sf�W_}�\^^~��n��֮Ss�ԩԳ���:�M ������=���r��Ln2)��
�>;(.h��TB�}��A/}��6"����;�Bd�p�!����%F����yyy������\.s�1/�Lb}Rϲ��&Ӵ���+7oޜ/}�H׷�nz����X�z�-��W�A�n
����;�5�`2�d�G��ftC�85}֬Y����v!HKYL�����	�A�����Hz�g����7[MF#8s��*n����R�<;nz��Ii��&gJ@�t�Ҝ���c6��/"2j���<VV��@-�V��3!'''�>o��z��oذ��0��ly�\d[l���i�\`���2�+pC�Dͯ D:���!�NuH|G�nowzM&s�?޻lٲ����-~_�^��C�CJ*��ވzC�AdP6��0F��T_s�ĉ���#�iܜa�d�[o�5������3m}<?D,�z��Zo�+�ZO��-9]nɠ3�"bR� =Jƌ��UW]U�;Ϧ}��B�/۫WS0��.FQ�P�m[���dn��O�ZLR[�G���cǍ����t[���bC0{��� (��059ψ�	ɣ���E�L�DMz�L�0��СCi.�k:�����Z18���vHIbh�!����� �����ѩ��'��95E��i6��M&2�2P���� k0��g�ұ�f%e�B�-d4B��OL;J��1U l"�!�����^oK�u�o߾I	�ۚ�/�����$04�_m�Vʀ��"'<�
neq������~�nliY錴����3gv{�A7gX�m�w�d�퍍��3�,�2�~��C����)]7 �0`���/�|X�%M�I���h0��F���9�QykF����������pG�z"�G���i��DM��L�4���/����V�������u7�3;/�5�u%`
{����{�%u����ا ����\������cq�:
���g>Gu�'�9^p��������]YY����u��f���2-��G��v��5Rn�y�nAQy�6:���`k��
�����+�*�A�\��A�Ry���4k�����c�i�6�5J��A:���n1�LW���'ֹ�^��􀅉/))A���	����յ<j~"ޞ�O7Q�'i��&=J�v���(������C&�#����[����2���*����}����]�	��)��!������2�w|�n����֛�E��M���`��B���Q�h���3~�p#�2vH�+�S��t�-�)����崹n�������7�V��_�jo�(�|Cˎ<����g����<x�ƩS���Q�Z�9-V������.��+���>�D�~@uu5:�Z l�P��;�G�#C�NѸ�t0�d��A�DM~\4hP%�}>��O�f�6l0�
7,b!��;h=7����Ko/f���m�"�S�����qچI�iǨMg��v�]�G��E�@~��[����K�e��j�hnn_#�i/�����]�Xɑ#G骔�Q4ps��������3���nv�<��ӊ�����0�J.�[����MJJ�i��[/������O"##�d����s`����F�	�����'���J�8�HWab�Z��b������H]M4ѤG	9���֭�imm�&�}�[�3="��������2�ϾC���p��3��)� ��+p��N�NZW�ǅ�(u��n��]��z��6�z����u��fC��vv9*E6��lw]B`��Uݙ���ܼ-�hPeEŭN����yT�qcc!4���)� Q��4]8f̘5n��D�����{-fs=]_�c��mujJ�X�<�^	҇�7�x��_6��3W���6���nGM4��%0x������
��:�@�x��C�::�B4��H<}ТE�L=��wj@��Ψ��7e�B6�[�fO��"A<ڙC}.9Ru~���9�:t�����.<VYY~�|�!���X�x�^g@�u<���7�k�j�<x-��;��Y4psdϞ=��9�W555]��p�I�s:P����čܫW/1�hG��6N�2e�����G!p㋌���Dn�����s��s�/w;�w"	�&�����=<��SG�X:�ȩ����ݬxjZ�&��A�۶mU�����l��F��r�iv@��.�PoLUU����N��9?$�Ggp�?�F�!�ֲ�Á�饴bwئ,�SR���� �����gnoҽ�Œ��"�^��&��6��nz6����<�d7��e�/�X>��N������ؖm�ɒe�r�n����f��H�⊁9~ƺe��ܹsμ�����\�T���1��ر㻛�����n�Ze8���M<%ڳ�2(����!!'SR&�չG�y�6uV�L����A98���sIOOO)�� 
Ą��js��/.:�9�!.����'�ԋ�/L***���,����(	a��`	p��HY�iz��YD\�9?�����Ԇ����}g�a̐����5$���=t�>J�|T.m-�vVS<�39-#ZZZ��uA�cd/d,�ޜ�I9R������j�>B���� ?0�|>p��=�r���}��شi��^��*�sfD*\l��������Z��Ȥ֎��hD�tD7WY֯_�\�q�ͽ��qt1�4yM����\ox�i��a�1��x�JZ=s��*����Q��~�P�?�,DM��M�>i#.���E}�N��۷Ͼp��z�Ā�f��E�"�*��vr�SB��|>��������� 9��X]�1!G(RPPp���-H��":��j#����B\Z��.�Ϲh����?آ�_�=f��^@���؞@bQ��L"to�@p�I�d�\�
��V��ż_N#a�'ٹ^:�}܇V�Z�p���J:�i?����)*���b.(M�q����njl�O��������*
�R���;����E���ٸ���Nmk!D-��q���LFc(#3c�̹3����/�r�����L����� �F�5mۥ�{aORN�KEmmm)}��~�sHM����m�0�>�m����Ia up��.ט ����8��.���p8,���Nˋa���i����b8�S��4���M#�@%7a:��x������F�E�T�5X=f�C�N�`-D��C���EE�Ϟ�����Ϗ��X�}p�>����h2ά��+O)�.��K7WQ;�N��^����C����e�X�XN��I�zAg��3�.)��I�s#G�zu��9�.%�Ņ^���$�H�I��ښma1���E��J	�%学�Z��E�w�k��Y�s���H��<u�6���nt������^��F��H�Ӄ)�юŽ�kD]�ts�v����V�#�N&��j��u_jE�����$	$�&�/��ؘ�_��� ��u��}�6���$��n����ӻ�Nz�G���ןq8��>ZB�:c�/5տ\�}ɉx|X}c�=�pɌ�:��J��Ͷm�g����� 
��}�B�T9�� ��������ܝ'N�s9��gU�vf�\m�m���\\���I���0
�7�������c���5�GQ�}�A��3���x3H�����2�ꢋ.�����_K6`&=�h����\1��bB�n��i�z�V�<_۷�F�{����$	@�����ʐ!C,���0����i��smzB�#�D����?@3f�w���{��t��i	��ず<k�Ն�/F�&���3��x����O�����ohXB�(���fdlP��.8 �Gg$(
�QNgF���Ĕ)�V�_�Gm.Aʊ�{

�jC���5Vl����N�����~�[>��ș����ch�8�����d��m&��ޝ.��r��@A�@���%�uj@��^�w�kt=e�����j���Ӭ�����>�}��X��<x��Fn���l��
�Y6��(������p8|�j�~��>.���?�w�\c����A�����4����o4�D��	MMMä�@觃��  �{�g����^���ٵ�L����E�( i)�??�`��3v����K����XAa�9:��*o�x�AO�7�o3|�޽222ܲ$�#h���oL6.](�eB�q�}�
K����|h�W]t��RQQ#}m�h �-k�̐�2@=0�7@�G��Y]]]h4������}��>�k��9uꔛ�5��tڹi�#Ԛc��R��E݃>r$e���g�뛪h���;X���%���S�1$����𶎶1[S��.��D7WX@��ꫯ�466.
�B�(J㜦�h����Z$����B�����6m�꒒�nI�K�dAQn��f��oP�@���;�!��k��Q��B��x<Px����h;�=+�]񼷷ঘ��[�E]�9A���ۿ�Tpӯ�@�(������~�{,ل<��Y۵t��>4 �������pΜ9Ci[����g�PK�t�it�4��[�,Y��)S�4��w�X$��l���4p���$p���4W�#��Ӯ]�K������
KUU�g��݋c��P($�7_X��-LOU���Xq3�h
�ׄ�W�zLo��tA�ҦM��322jH��d�d%��9b7*�x,����pg�竭��l�F���}n)s	�㐬���5'��Ha�����F:��F}��MvGGR��A���;�&���z�h���~�L�n�Mm�ٳ����9��V>;��hq�'os@C��-��/(E�v������Vڏ��yv�\�#��{����
���y�r9��:�������M��·�!O$c
�~�=�%#���y2��j�22ܒ�����ܰ� �B���2a��իO��+�:��l F@�n$���Ѱ�o!���ހdKt�h�Z��M1:f�I���RT��C��_��l���� �V��;�l�.#��.��ry�n� ȋ1���xpm�� @�T�����(� �����s}~Q
�V�$i'8]kC�D���I)�?���r�0���'\�~����\���iQLl2��v�V�}�K�6��G``�-..n���UQQ/+v�����f����F�������r�%�řv�q�F#:��tlF�ƒƖ�2:�z��K):����{����=��c1�y`!�PC
!�4�a$�Z̐����t��ѣG��=��'yyyѢ����O� 9�^�#5�x���������_;9D��DB�׍E���c�J���]t��D����Fe��"��,*ȱ�~����"�r[[[n0�Ɛ^��r�^������b�p���D��{6\[[�O���f�S-"�
�1G��)6���664��B���+����p���Dl� K<�����'��m�Z Z9c���vK8�B+:��B������4oG�"6��Y!��!� �6��yT."�]���A�́ɓ����^�����W�X���#��,rȫ0�'�\���Pp2��7��h�\`���[IIɸӧO�׻�]t����2Az�T�t@�pH�vK�G�2)�F#����l�������!��+;;���q~���{Gж��ʠށ��;������������N2�+3��N ��l���]f'F�Z��皜h4����H �I�_4Q�n��lؽ;����݁@`0Ri�ZI͟&U���9 �7)Z:�"Y;f̈Z��w�����=7'wSS�(���tZ�~Lfp�h�j��q���3H]�/�̯st��m���-�ύkhh8!]~]t����QM��ϵ�F$&��m۶�C�Mss���M	x�����6�[BN��;??��|��={��j�O��Z-�F�~/o���wi�{�t�J(�gώ�Z��xKKK/��LL"�r�����5�x�`(<��I=o��:S�\A���u�f�4���cQ�!%�Q����ʏ+	��J)7U�<��r89�M�����@OW\��������KJ}{(�P9�B� 7Pv�AS�[DDϵ��<8��բ��e`�9<2 y#G��x����nt��K�� 6D����d��egϞͪ���a������؁���� �k�{�y�hQo���N��˷���1j�)��u��YYYMS�N�`pg��G���9�@�XH�6s��։D��xo���F�:�����c҇L;?���e�	����9s_0N�Z�#I��ȟ�0�=}�5b=���t:]�����O�<��^kse��k���^:Vy��I��W�,V<Vp N �Nx����a=��1NC꫱�+"�o������v{YY�2p����z�N]��ӃE���huZ+ZZ�)i�
�����1���9J���$�dK��^������ �^���~7���d�,�<�mg�Va����}�k$Q�w����k�X{���;�<D�q<�93�s�ݘ�
����=�;���s0�D�.��F7�Y�ǰV=:�.Թ�==���Ȩt�Ȃ�XJ�x�8P�\��b�6N�3����wʔI(��	����5�~o^���٤P&NA	E˾�w#:�Dt���u�zUZ�a������|����1�>;m׮]{%��O]�g@���M���x �?'[�)@�/~��,�Ԙ�Q/�xhx���٬ :�Ǝ�����j����1tY�"i'�smذ[�qL������P�j̘1�=o~���s�Ir�F�������ޚD��vr8�[�qx�u:���r�̙�����c�*���ۿU�`�F��C��v�֦)77w��)S���͕��������w���w�����' ��.�̂�W�!\�%r�����ц�9���Hͭ�n<t,�y���nt���<_����#�����?Hl'O��A��7KVI?a;��x�5��΢����s~��=�������sgg9N�6��/r��(v�T;����M�TUTT\�s�d���я~Zm�Z��d��T[w����|A &#�P�������(Ptps���޾l��|>��1Z��(%�H�Q6�Z�8����L�Y�u"��������t��6WX�;z�ކ��S�����p���AA"��x����7����� �uDw�Ɔ��g�����M���d-**����>������R��F]�!a%}��Y���Fge�ќ�vCM�������?�A����=~��4����O;����ئ��4�2H*�B�T�dɒ~�#D�������~9p����7N��D�Vy<�jL���sWZZ\w�lM��2�"�u�����~MLn�H8�`�/�/mjoʡ�/j��n.���`��u�uwweq�M:o���9����@�-�t�݀骒.W\;p�@�[{�����3':ٓ�V�C��.�xڠ�7K���7@�º�iefN7�h�e��'`����{�ѣG7�:z�N]�!gC'-�|`
��ׁ���ـ !��կƓB�Z�j���I;F�4��6dC��NMyyy��m����\YY9�l�p�QѶ��mB)��6f�·�vɤ��u�L�sC4F�0kSS#6�z&t'���N_���[7�I:::���=|Kk[�X\���v� ���0��mĨ��HYY9)������5q��=�>��ԩS���m����~?y8L��>.��sDc n�::�5��z��de��,Ɯ�bC!�Mwpz�9-����SO�>=���x��t�E��M�Y�������� �6%���N%э<Bv:��N�ɓ'�{��Bs0[�{�)/��N��II��H$%S=a�Dyw��QRWW7��tdq��v�9+l�w����l`;٦�iӦ]r� //�O砖l����ߍm�8��A,���|��&'ɼ���܋ݷn.���X�e��ֶ�;�F��7?���^XuXXR�k�'jm��ّ#G�7n\���Ut�޼�DՑ#222
}>���#]0�u�Z�H�7���^�n?n��	��,�ޔ�q����!z����E��O�m�f&�,�Ŭ-&f�r�0 I�ͣ�M�OKeee���^&shi��3cp��F�K����rrr�dee��)@���}}f"�Vj��@�|��a����9j��G�~tb`��b�����a������m��1�q���^}���@8\��s1[:������>q|^0�HJ ��]�����<7L��F�E���ࢊ��d�#~@��i].N&��ж%ۮ`�7�@KZ�E�%�����.W2�{��&γ�uDo�0������� ������)�Ν�[UUU-]C�.��riB����D1h"��;�����v����f�f�o�J���o���N è��r��kRvN��I��RZZzv ٵkW�}�n%{RD�70�т&(�Æㅍ�"�������ܹs/���9S�����>�~�������1��K4)��J1�F7�(@�[��:������n1f?.q��H?�@�))=[��v�;)B�M�F�Y_VV֨{�W_JJJ�ƍ�����x<����&������Ey�p;����
PP�����Pd̜���]	2��H���m�Ed�m߾}7]_��׃.�|<���j'�.M���o���ڨ�eq��^�%�n�mۖ�w��Yd#�Ѻ迶EZ��JG��h2y�"�жjժ�6q?���������P����|�,x��������q-{.\����}��Q��~�����d��վ�=�_�d�p8X@��tps��P���p����Q����oh
�����8���qc��_�Z-����wǍ��ֹh^].^�ؕ�����<�� �26�St�V}�E�Qs��)� ����#�~WDr ��V�%E���`�Ñ��5;;{2}��͛7�����r]t�����Mz�G�i��Xq����-�$1Z�����}k'7n�8����sd+\t/�bI�O0�o�#�O�l��>�w������_��^w׮]Z�{� �WF�����1���1(�8�	��e#%��o2;t�x��Ҷ���-����X2e�'�^��(]����(y_eeA}C��tSsd��QtҘ���⸰�tڿMF�����N���A�J7�3�S��c�����Jwm������$R�~�b�V����`
>��.9�nph�z�fc�W����źMMM�Æ�魷��u���m�ڒ��.�\� ��裏"�̄�����2҂~�Qz�F�}^�P[[k����g�-a�)u1 v��遘b{�GhA�Z��LЩ[o�5��P����nrMM�<:'wx�}Ѧո��C�Yu�z����2/g�8777L�����sb�s��xi�C�o2�4�)97b�|�E7� ��ط���@`f(5&�)�l�I�8]�&%�K�%3:o�E��xB����.ވ۝�Μ93wӏ�t�؄�������S5;B��Ho��4���(�m��0�^
HA!�5���vl�8HFN�A���|B�y�ap��jUxs�`����7�	Ń�g���@�����;�Z:���t���IUU����m�/��3�H?SJÒpP!`0�5����ȷ����\�6?��φ��ȕ��m�XF�)�����~Tz	�G �V�WM�8�J[h����~����gƺ�n���d\il��`��;$�Ն?�T!�F �mw�M7�y��'/�y$�=j�[ϚL�(�*;lj��I�\c��(
%�o�k�p$�vGm�_�\�����476�H7��A��˗Rx���F��)���D�o���J���9z��t�$]>vA�fȐ!�跽�~�������ݠ�&''G�~x��L�M���@u7}���Q;$�Ş&�b��\�G���vg�km��,[�ׇ��E��$��w��Ʈe'�6h���B�"4,^��=WM�6|�j��#�o�H�^GSk���'�O�x���7cƌ6�v��׿Nhii���pd����;�ũ��M�#u_a�����7\�.)��={6n��[�y�j�G$\TM�m�B��/Թ���E
��+K_�mo�,r70�z����~1;�(6`��;F��qg��]�''L��7;;[�4�ћ�۷:s��R�")v n��cx>�����
0#a��'�R����.���>������O7Z�6)e�+.fC�;dl�oavvν[�l<�{��s��љ�u��
���/�8���5�t�"� D[L��V*X��{^��o�j�ﰦ��y�E��HC�4<4)M�6����C!19Og���K_�R��_��X�رc������BN��?�\k\��C2�x!���::�p���馛��x��z.Q��v��N�5�2c9_zJ9)t��8'��@�n.RN�:�]}�Ԓ��7(�ʩdLBcTJ��$1�C�ɢ<%
�!���v�(�j��KJJ�:���O��fd޼y����k�������<P�=!-�q -.V:%D��0������h��-�t�R�3X��ˡ���H�2���y��W������������g�Z���&�������ֆp�J�A'SAAA���nڴ)��7߼�ޛc6�,"��h�c@��[K�ZZ9�B�0p{��G�>}�6��d0��r���x���֋�����n?��_�2�����\�8����݇���y 7��Vu~�h2Z	��UUU�d���J
�V�\Y���:#Z㱈�@�E���M"�(R"�#nX�A��L��rf %�����Ul�x<z��x^o���������)���#jox���(�+,,�QA�OD�H4$�TѨQ��x�:0&0"�2vQ(�����G�2��<:^##+�3fB]ݹ�_~��&���C�颋.'����mmmH���ъ���`���7�"�=INH`�g_���*ȑY����K` ��4�v���沆x4� Ҝ����'?����?���.�+V,&[1�l��[���D|a�p� pP+�))Z����I�&��Ru}�� Q���}Fj ��z.L�D�M��;�tpsR]]� �|3���]�F�PE�Tӟ�(wI�FT�'cq�I74]\tF�7n���N�kLfΜٶgϞ5^�w!�2�#%�^"-���Rv�G��z	��HMR�����%2r����v�,tD��@�f��q��Hq�;w.c�С7UU�?�����-�.��rE���~p�Ro#P��|pW��l��uW�:J��nr~�����E���立����g�ܹs9;"i��Ǔ�~L�LȑlWDv�؆(=?8y��*M������f6�ϑ�qq�>������`� p��Tx����>�w��فg�}���Or�c�l��\7i �a��x,�����n.Pp1m޼nTSC��tQXcHG$��b�R��RI�h2�I��	ɐ0����F�Ùr:��Q#W�Ŧ�^�B�ݺu���ƕdP�A�u��0�'"1v�U�x����{Q����Hmm-Rv�G��pâ $��1Dk8��948E�-�0H���=.,--Y�s���ի_���b��.�|V����ݻwO#gd8���)��tGt�>�3�m�^����<���3gθ���o�>w��fs��E;�Ee� �Bڗ"@R������;�l|��g�m�V�r�ʻ��h��cD��bP� ���) l�Ώ�����~�[ߺ�NvQ�K���
�~'��e�2dZ�)�M")'�q�@�":��p1�<Y3���{nT��r�HH5�7*���e��	z_U�l��Ns9�Lguy���H�H�\�2���cǎ�ioo�K�c2�@�b<Rd(�RV�G�{v`� N`��#�r)E�x�#3Pa ���e0��ul�!���:iԨQ�C�Y��s�D	�s��9I]t�lB6�S__��tݥ���)"~�힂N�I1.�
�EV�y��555�� ᡹h/gr>u�/�]��Ǩ�9:mڴ�܁E�5��G?�{������l<�J;�I%Az��FU���Zw�ĉ�hiD"aJ���W���;���Gg��1z�^�\i9~�x��C��'���4��M�`$��������"�������s���`��yy�ZI�kVP�RYY��'V�"�455�e<��� . $�*((H�����46��RRR"����Dx����:NfJtf*���dt�aÆa͗�y�)Ú5k����%]t����W^����<�l��6ܱ����و�qW�;^'���k��Ǐ��m�����'?y��pL&=�����5p6@D6�^UǾ u�����e�7��ͳڲeK��+��}�̿\���q�	��a��~GG��-jD��� 9LG����_Q�5:MI��F�plZ�����_��J6#�}�����=���+Z[����O�_�Bt�1�0Z!"�8�,�}>�bWr�h��t�H��fԨ��t�wK�\�#5k֬76l� b�{�0XP+�`y����"���DG�a y�Gw�Ǌ��t`8�Z�4A )|�Yx����5����u����Y��͗>�����.�\��ne�:uꎮ��b���n�F;В�w%A8�K��F:}t�̙,>|���C�M�|{~~�c�s�۴!�s1�Ne@�6i�
�n���rڴi�.\(",mmmh��;���n����~<<��o<F�A���)/}f�M7��t�ۿJ"a������x ���{.h�57WX�y���{��Cbֈ��D2(�15)�1bQ�FH�d!�M`�bIy�F�h��E�xA~޻��&���5.������VWW/'�w�R,��B� ���Q�����X<"C~2Nq��츤���JO�Z����¡cDq��� A0\��c��744	H�����_L9�$�$]t���81uuu�	4Xy����~���iu�.�m���83u��8�@?��g<x�����|D =�	��mJZ�̠	�#��N!�/^ܺf��u����fҾ���M�L����v��#̽��V�]���q��U����|=�G�(����|'H@銞[�)���>�a�.+��WZ:d󶵏���M0E&��u��,S	��Ź��S��21D76L��9]@Ϣ��l�ȭv{v��i2���4�~��r֓�?+++���C6D�X �{a�����X�� # (�`D������Z@��l�clޗ2�Ӓ.4�"�0��%����G����_y�'[�n�����[��J].\Ξ=�q��ѹ�c#�]��ݍ�<$=�̪��t�t�(館�y��'g�\������Y�XxH.�)���?�M'�p��~��t��vvv�Cz��+_���ڻwo�sy�[�x|��Xq
��@
�(��#��U:�٢v�ٺ��{�j�J���.�g��=���aA!1�+3��o� :�� 	��r*)��dB��d���eLI�P@*�.�J\R~F��{�+d�Nw�Kq�U�M�;�%������;:��b��O��D�������������x<����)pR���!���S�4H��΄���%555 ,Inw� ���{�Ŋ��a������5��X�c=8��$-�n�~��m۾��c�������u:��E��S�NM�������L��Ȥ�7�'�͔$ �Lz���y�|;v�(y��g�O�;����u��s��I�bƓ Rj7&�GmHh&gf��ŋO.[�u?���n����j����\��)-N��	�s@��2��i����óg_��?�A�>x�ϭ�(j�ږw�9ն�k_S�q.8%���HYA~*�'��TJ\�f��g7J��O*�vKC=ْ)�R���ƶɟ$��(�������+��"���ԆfggQ&���E��� :Å� 1L��C�bb���b��?�`��Ɖ'è�;�`�`(��a�Ǐ7͘9��ࡃ��?��G����}�^8��������|ggg�	�n�ֶjk��	' %}=9v��C���G}�n��9���nԍ@W��\�+F����b�sY�%E�jm�c�6��0"����o�nٺ�K�5$�8N>�a�p�`+��B�1��d�+c�m���p��@Q�H�g��LӇ��h�L
�p�}.�8upsb��%��X� ��9YR��$��^��IE��1�H޸l���d�PJ���S��pdz�F�(;@/%]>q2~���믿~�ƍǒ�����)��Pq /06ø�(N�;,`�8A�0�<"m%&�+��-.����<|���S[[+RT#�������W^y������^��	"u����nݺ�'N���@�ū��8C�i�d@'�9 ��s{�O��}�g��}@w����܀�@��� ��r�ل$m����p�����Μ͛7Y�ץ$�)h"�t���BĆ`W8m�}����;{��mK�,�_�s���d
������2 P�@B�b�����������Qu��?f2Hvg2&�����R��.}~)�f�8]���+��:�D*�p��1���Q2EI���}��w���4E� +��2��J��^�k��Fe�����O��pdF�A(<Fʋ����	�U D0l0�X��L�TD���������g	���Ϣ�E�������={�����<
t�� ��J��x�$�!��|4�z���@va�޽{�C�% �M�>��E��A���TБf��)Z/ r�{�wÝw�	�O~��/����E��DW&�:�\�k�&��f'=֥��Wد�������T��cO^�sL�b��m�b����I�o�l.}6�����\����%*F��ط'��s2.g�,Ҩ�R��IN�YJ�"�d��a��j{%�䒲\�R<il�[���v���`A$�0ISS�K0�o0�J].��FB��Q!�C HxN(0N`.L\���1���b tO��Y�	i-�hQ�mE�kf�U,.�3��0X<w&H��LH�����2><�޿{۶�P(���ݻ����u�彂��SO=5���z�SG>��7
�kYL�� '���ᕒ�ӑXNZ�3[�Z�nji6[l�2�V��"s�/��X���`�&���h0K��_8;>������3�ǎ^������Ǐ�������,6s���0�,F�mi�> 8T�u�d}���X9%N2�-;Ə��c���Wu�!��]��������b-�
zRKt����(@���m˭�<:�('��q9��}oK�Y9R]�6��IQ)H�A*,&uwI�-�TR�|.�{��Y�����d>�6ϵk�.���D��e��r��v	�S�O7�ܠ\����"����QG`��8f>f�����\��A�9�"8x������_:p�s��ۿ������+^��]w}�E�n�KZ���7�СC����$=wSN��9t���PW��t�D����D��� �!R[�hZ���q�\*��bQ��x$�*Lz�"���n7+���-�{��g���|����>���d�� _eX�Q#l �yᴙJM6�ڡC����|�Uo8������ą�J�N�7e��U��E�PNN���`s����W^Y�����d�:Z�j�L�Y��8%�L0J�q�H�ڑ풲���T���^��V�w��<z��FI�O��r�-�gϞ}q���IYo# cQj��aP�q�����Q	ӘR��E~�����(15:�����s��� ����RÑ���III��#�鹭�"{�<N����涜7�X[��}����ӦM��pt��KKK�EħO��E:g�x<2���,w:A��T@�ىɰ�8򀈄�����`V:�6B�����!�
Ń���7��wע;�Z��}�k����	��#�w,m�,�m��q��	@ac l8�H0���>:�u7�����]Q6⁲t�R�֭[3����g*p���z���>��zA񕐚���g_xᎺ��*r��ý��:W�g���Mm_4�d�$9s3q��'.�������yc�����ŝ������omm}�������p2T&t?A���6Q_EFk8r�C�MwE�P� �O��ap#F9�,�,��7�	�Ց&�1��Ɩ�����B�����嫫W��ii��������j�t��Z��^|��)G���t1�t���3�uč@:�u6�I����p ��A��r_���H�Rg�������p����<�d9�ʪ��������1ޚ��+�t��3�c_���&`5J#�tx�ؑ{�����^�s=v�X#��\�sN�������Z�C�ŭV���OB�@��͇H��i�^�}��'73c��l0�-���K�T"�l��F#y���ಧrJ����+�o���f�;bܼ�|����l	BO���~�r�o�wT����	f�U�����*S~E�;�Z[���c��ϛ��X8C6h�C2[��>R]!���gBG�sWg�4|�pSIɠ�3g�|q���!oj��ŋ��4�.�5A$�ݻw�#9�	��+�M}?�kX�Wx�0�Ӕ *V�Y��xH�<�y"���bpb��*��;��z�D�n���@`�=��w��\x�_8t�Н��<:,ݗ\4��/t�mv�4�E�7m���h��߾�ݏC�kjjL�]�b�sN��L)>_��b������RQQ����)�c�,����u�vn�������LWf4���8f����E�������H�E)��$e�g�2���C�.�i�FY.�۾?Ų`�������{����_&��CRa`�&%}�5y�6����Q����u��9����в�K�[� �K
�<���۲�mR]ݹt-�G$Gx���t��	iĈ��ɓ3O�<9�С���Y}}��>��T�|����*kժ�-����鑋;��c��(NGTDa   6�S�t��f�Ѡ�N����;&u.GtT�����������΅oZ6c܌د�녛6n�ف���L6ۀ#�uvx�ǈ� �p��C�_�
Һo���W������D߷�������_"�fbm���z���_�~up�>�9#/=�ԔM�7K2Jӌ�5�eMY��'3s�M'/k:����Iť��n$v�����6K0f2u�"���R���ƍ{�ȑ#C��ĭ6�|
Ј���9=$X Di�K 
��bءh� ϭao ���4!���RQ�ں��GD�Y�۩�o��fs��G@�:y��s}z�ҥo]M�]t���,�l�tˑ����3RL�*k�*0�@ �
��]T�,+��W&w�
�f�$�Ǚ���p�ǩ09��E�o4�+ڝkF��b��)'��mܸ�[F�q��e7��8 &�E��Vr��HBԆ����NG�ȑe�n���Ə���@���'�G̈b�.��X�!�!��/�	G7� �W�}v�����)]8l.�S6�Rf��+�m��}�������x��0	���dϰJ�]��ϑL�I�;O����[�'��{2\n2d�;:�vx\ هa�������������!�����=���P=�s1�dưM��"�^uu��}�ν	Fҭ�x��/r�Ep�:q�j��e?�����7�di��2�˧S0I{�ƍ�ߴi�wSRr� ��@&�C���3��o�aD�L Z�rf8�,�Z�? ]�* 	��9TY�_z�������r��5���_}mُ,f�,Z�Ɯ8�ʁ�3�8��a��6O�VSR(ĭ#'��E��;0v�؋"»B�+��7���J�Xߜ��3�8�N��6-�W7�C l^x�1V�������peĤ(f����o=���?9����u�f3�9V��M%�h�J�JO���ڒ��9n���gB,X_�~�a����WF�{
y,f�k* Qڼ�Y566
��؀�d�#z��ia���0aNl��+`���a[��y���ؕ���T��ۙ��Q�QM�h����ױm2����S#h[_۹sۘ����W�\��;�躘0�.�\�Bz`y��f�[��K��Pg�H*,�\��7XD�Ox}�� r�3㸨W�Mc:Ŭ�Ce��Ĥn�]�_�=��a=5��
�"�]��-�c�$�/]�ڷ���f�.�s�A ,�u�8O���P����<x�̙s	��x�?������8N�ݙ�����4�	3�q��s�̋�W���F l��G'�[���N��֢�O$��dhPN�E�����F������޶��P�͖���U2fX�=��f��j�I�|�d���;w�_�l����O3220����*�1��a�HOA��.�F0! 
ovv��Ŏ���E�0l�XX�w�6��1�q��b[�ހ0|��\�C��p̘1&S�t��74����O;|���>>I]>�.���W�oذ����]7����; '���z�(*�8��t�!-�HGf�m�%�{J�1t����=���3g�|��`pj��_��캓t8�7|�p�p*=1��c���ݜ��i/�#���!Ö�����QZٶm���s	�C�7�PL,yF���1������:�ߥh�y�;���]\7؍�B�r*�V�e��.��=t0����C2Z�q�M�x�dvɒ��)ٲ�R�"���O2�����Ϟ̝;�k�ҥ�H7���-������2rA0�n����CX^^.�wR���qy��!��B��\�N�%��l	x=	Z��� KYY�d���5uj�j���#���H\�Æ�;;;mmmm��ڷ��MM-�?���7̝{S�^p��4̈�  �IDAT'U0�qժU׭[����s�#���i	5��|0 �p0r���+�u�K��]L`X�Q��N�������m�ui��?$􌹪��h���^�;�e#�./ֹu��5��~��A�@J�i��t�-��[�הh�c�[Rq������3��%��z�{?n�a�5�d�r4�5冀��mR��\� �銊���?:��T`��#��nZ�]wf����t�;��T4�;b�Н��q����p�,�G7���S���%.[�?��dGD29M�=�Fe)b��,s@��:��gTP�K �͕+W��bѯ8�C0�O� �L����b���{
�S�N��I����Ǟt��.�U S2����R� "8�4!�Ëu��"č	�����E�0�<����VL?q��o+W�ܢ��t��	"�[�n�b������ܜ����z�e0��,� 7���0:�ZDC�0Ew�(Ta�s�E!҃.a]����㓘?G���c�Iұz��7ǌ)o�w��*++g��d��̑����-�S��͜;�+���|����h�o̞={�Ǚ�b!;�
����:T��~39�3p�uS����M�>~�"����_�����zk�?�.Y`�;<-�M)��ܚ_\�yɽw=;���w�	�v��g����t������D���PgFB�[#R�KIo$I7�e�)�+V�����
�3ZŅ^Ó�'�]�n�;4y���X���hB��;I̫�R2�FN����2jz8��#��|0�N�t� CH�y�^3�Bw�XՔ��s3>���ݻ��hv�I]�uI�jm+V�(_�r�O���X��l�˲14P����݂. �C $�?��@S�"q�Y�L��x�i�H,M�	�B)��$ up��!MǪN|����w��� b���`D�-9-�S l_�����f��8E��O:�iҤIK������ߐ>n!��O�6����d����tGs8�M
����t_�?���Nd�s_x���gk������&ey<����d4i]6r�7x�O�'M���
Λ�y�d�����L�|�ٙ��LY2�eIr���R�M-R'��t/�3, ˢk�l8l����[L]]�ȫ+��{L����40� #��,p`@����E��A��Ǔ��2p��xc��1iο���=ODo��Ry5�qb}�ŁQG��:������2ȥ���铛������o�}l�̙>��r-
����_�0g͚���z;n&p��� �|SU�Y�$�U)�ō�Q���N2���S��UI3)���}e� 6�;'��o��)�"����ȴ466���'����t;�D[���9q�Vxa�xMD�z{�_��<��)���������7�p��k���������:oƾyR�`�~S\����Z�|\t��gܬY�����޼���uIɠ��d����(nH���Y���E>z�lU=���ގ�/��ri"�k��P�'���c4g��n2�0]�ɘɔ"p�&..]>>QNK$��L"C�}��!O�#��))*�Ƅ�'e��G1�bP��tw�ȸĘ�A�F�,&�ܪD<&xu$������dH�!%�2i�F�!�����8�#�t�=m���t|C�~{��'�6TUZG�����To���{�Z���u�6�S ���p8\�l�����i����PjӠt �-RTL���S�XW�%t�@��6��*�܁	GU�#&��l��s��'��:N3;;�{Dry�
��|:x਻�+��uP�G�-��s�=�s�̹&hH�y�����q�!-�s��m�Z�b�N	��-��{�����A�����i�_�{���ޛ�)�L��A0Gjg̙���������M왶nx#�����[���f�dsڝ�`0�;d���hv ��N:eݮ��AW}H2ڼ��&.0]>^Q�R��֭[�$�EnU �*N���[L��B�"8pd��--m"}��o�m��[�Μ� )�a�[Y�C
��� �0K�e ��>�xMrܴ��Xt���;�ٳo��/��e�С5�g��]>.�H'yϿ��]{v��f�Kzc�kZf���U�@���dJ��^��%n��� �� ��p�u�G/�\�<8��b�t�7�:$�4��R�/�@ɤK6�~I����l�o�!t�;��m���I��0��l��p��O�~��	�\3�����T:~;����j���c�kSV�@����V����3n�;�z���N]�~�Wmv��Ņɘ4�twG¡����r����濔����Ϥ}ny��l��w8��sҔ
��~��A�s'���=vK��`#�i´W��\�&�L���"q����h��[o��$�t�۝��v�I���!W
~;::�ad0#�(JGG�ʂ:DDWx��bw�0�6�EtT��}A������:t�HQ��w(�?�8r\J4)V���#�����A�0[h��x<�
ǭZ����ܼ5��ջ>\����r��}�JW�\�@��#_��ʬv�E8I�X/P:��v���8�J�@|Ks����%��z
�݌�p+�K��lQ�zʅx4!t/B'��"�Ujcb�0��pf,�����tLv��7���8���{�t�c0����K����y<�gn���(����|�gPo3�������(�+��>����F�b��$�XWQQq�䃟p�u�Vף�>|gSc�9�ٳ�ƑE�YnnnY������?�xÂ���6���ğ�0,�ٶؖ�vۜƞP"�XN;�UkQFe���8��>�`�R�S�5�2X�6up�KZ��f-����}��)�=�+��+3M��\������6L(=F,�6��A�6J�TJ,�XH��qr8������TRRJ��.�M�噃C۪�4������� 3{�=E����Ohii޷gϞ�O=����6��*]����oٲ�+v���O��N[�����f�f�;�@���(545�:7��aCJ��z\@��jb�b�x�R��N� �7�9��i.0X ��N���clH����a�'DQ����h,43� ���t�1o޼�_��W[����I׊��c�����߃����@8J�iy�g�c�#���A�t	��O=����'�_z�{:�ڿf3�F8�P'B��7?k�ۋ���ɳf�����W�Ա�o�U������9�l�]�_�|6smV��K��y-b��Jy�1�C��F�@�f�9i���fu(*�9B��k֬	�A|��A���g����e�I ;����(�'&<R&��v����t�Q�c�ӌQh �i�d���R�Y|.3�#�/�Cȑ���l��������������޵w���Ə�R5s�̀��\n��y��9������;v����ֶ9tS̴��ɀ�<t�FL����-^G�7@w���T\�ڔ�e�I8ݺ�D{�b[x��E���S�y���d.���\�,"3.e^�ٔ�9p��a�@��p�#G��i���,�9sΟ���o�_k)�'N�����H�̍� 7<�灇�B�13�߱:77��޾h��7�O��>��CSO=r,�� /��f5���хw��|�ʻn�g�ԹS����׺�:�޹u���0�v�c��9F�M�D��·F̜�V���ЉG�t�He��)�=I�$]_&CP�t�3]�+j��)�o������}d��oj��e�l�aT�>j`��G��G5 t(���P���m�A��
0$=����S�M6�����b�0����*�,Q��=��}Ho�=E�r{{;�UE��\ү�7n�{ǎ������ۛ6��***��8�����Dk6m�4bݺ�w644~�������ź�p�ߜ'&���P ��Qn�� 1 '\�
���b�!��}�����ǔf	�0{0�����v8��z���沲r�ݐ�>��|T�Q��QPX��lԨ�|���k���y���g��Ϣ�g@����>�������y�����R�ۧ�,]�������6��~�N�₢�d4tx�B�tr��O���+��5�ϳ|g��q�������0��,�S���v�L�,�`l-Nz�?�kJL��K�e��H]tOU��5��@J���˗'|��l)�A�x��О�H���p����Za�����p��n�4K��#�J�D�����j�K�Q��M��d(ɂ������U������t���&>z����|w��!H'ߝ<yr��͚��'WP7��SOL��΁/�47^J�m6���$R}���C�3X�<5�ۑ�?�M3���KR�9��y�����	�(�|�(��� ]�~`]�S�����a�Tn�J�2����yl�#
�U��,))�&�Z1~lşgϾ�Ե��7�xcľ}�n��3G�����S<NB��y��A:ߧ�s��}��]��e/�e���B4�3��(7�����H�%ӝ�kѽ�?y��A��GB�ӯ�j�m�~v25�n4���M�&bM%c��8~椷���v(eN�l��l$,C��'ɀ�U2Ȓ.�|��]T'i��Ν;;N�:�MR�2�FY�v�LN�g�� p�#:�@<���[Z:D x�LȝT�	���҄�0�L�	�f���ž�c#Μ9�	�� ���]nmm5�{9��Yt|S�ގ;*++Onڴa���_;g̘t��`����,*�]V�|����8�l�2��������D<Y�n�x,)stM�=�����@���0G�e	����Z�)X��p4E)썪l�mTE��a`�]@ʼ7;���1�B����;���^�CǙ${М���f�葏����|�El?�������t�.�vq��3�;ošs���8hР×:��SnR����?Q�����{;ۿ��t.����Iʲ�>߹)3f��p�o̘1�0]�4Z���ғ�w�c�,/��N�:r�����A;�V�]-�]��u�Vc�l�%�r@�#�d��$rqup��G��j^�b�32�uuu�b�"�`��l 9�C
ëN�]mmm�-#>���.)��,%	r�m�tk�Rg Т̲B���*��x�v)7�& :?�|�
<�!���h���A����(��6�\]]-Ӿlt�CȞ��{�wv��ر����>}��]�v5]w�u�,6]�#��v���'����G���n�ףN���Q�WK�t��g �qC x@�Ƀ+�!� L��K$,��h�Vtѹ���DR��*�ߟ�;�tqR��d�d0I�*"��֏��z�,
#��[f���ۼy��$�l���yy�����p���\S������9r��tl��s��N��Nz�031�v�C���49J��� 7[�.u��o�=w�v�Y6��t�G��rƒI�tf�����+�s�ʢ"O��8־�ρ��{W,�Ė����E��ʊ�׽\8&�Z����J�qD��)5:�>7�r�E��(w�}w��o��쫯��SUU�=R�2 &��8Np��1�cWW�D��!�ϐ'�s䇽�@ ":CP����~`��}�����
�:�_��| ���Y���xVϴi��B4���Bz�M����c���ٳ�r�m۶��_�'�ӭ��t� 
��C?}����Ͽ��št]��s� X/�X�wr�E��'"������d0���Q@�ԑ)�T���=���/t�P�����FIa)���&��s��(�� l�<G��J�~Fd:��<�@$����=#��Zy��?��]�`�5ǡ�l�2�={й���I�| 
Un�tm��0Q�yqF�n'�wɔ�Xp�Xee�}���S���En�d���N;�&q��`�n��Q����_����d��[��/{�m��Es��_<fK1�|Co$�[գ'��c�Ԓ-r�m��n"H��T$)2
�I�R�\T�k_f͚�z�����H4>|��I�g��v��a�%=LwRq�9�<T����X�5*=��ۼ�a
�*�l�S�:,Lc#�m�̷����� �hi�q\ؗN��yr�D}���L�^_��~ҍ�t3;�cǎݿ���L�<���	&D.vp�.�<�]߰a��ta�o�����.��ib*){�@��[�U�� ��k ���nK�����d|Bw��t���ruEŁpz��	����@@���چ1���&�O �c�Ϻ�b �e����4��sbB�xxȐ�3�{/�?��_����Z��۷��y������8�Ā�gF�|)��t��%�\�������&�!����_��fͺ�::�6�m�99�e�"��/���/�~����n1bD�����gW��r;��_�L�E�8��1oo�v��^̛<a�\~�{��T�F�F�	�X~��.!ӦM@����O��&�R�[z{{=0�ඁ�C8]�.�tP��¨�P�H�}��[�� ]��|��2���~��硝��xU�.n &l�b?��)`�6K|5}��qa%GrP��.t������ˉ��d�� �,@����=zt�o�Y5v�؞��2��X@�˥L5����GC���u0?��$G���9K\-��j.���l ������C�Ƹ�9���\b�ө�y��*����\�ܦ�0+\,��<�����v��z�7y�#ǥ0ӱ����\��ְ�IWZ�0q�ė�_�����t-�֭[mO<���m��91s�3��2����Ӆ���I�w�#;�x9��n�D�ׯ_���3��l��[b��D�'+߀���6����zd�����0wM��ٵy�����w͋��֬�����a��V��K��h���?W6m����ϛ��G��6����knt�h!��>}����<�ڵk}dD�"C�K ��S���p��b�J��2��3J[w�t�d@a����Y��������q� �Ra�kxD��$����f"xr���
��`I��w�T�GMY�ȴ&�[i��0�@ѭt����?E�}l�С[^����ÇwN�4��NWJ��t>�P���/{~������#��st�L�K*��Ck"�2�u��6QTڧs�ӹE{6v.PU�J"J�7�� t`@��1�S�}�t�GIA)�Բa����b{
��7]Ǧ .K����(<���ڇ��J�:�)�� ݈�5MK+*F?�����Z���z��ӻ�q6�3oGm ����1�D�0ӋtQ�8��Zrb�/Ǳ}"���m[W��_��u�N�\D�N�#+ϝGW����@0X7�x�����oL�=�ć���#4�ZV�{���9"��[���V���Ǣ!�p�d��'FΙ��<kV��m���D�`��٨��GF��H��r��֜~�W�����k�z��n�d��?{��ue�ު΍�� � 	�Q3%��HJV�r����Yl�����Y�y�{�g����=Y���e%R9���H
� �t��gW��hQ�d1 ��X��]U]u���}���"5f��89�,# ;�tmsx��(��Ch����[��0S��ض�/�혱O�$������SA�8<�o����rtϜ��a �>�
���	d�:J��?s%�c6ms+}~��ݻۨs�M籕����^{�0��ٳg'�+H@at���k�z���_�����#���eLq���Hw\(��=���M��آw��}�0!A/�yS8�[{�}a� 낲�*��'�����X��@���`-?#�h�d���f$keK)�c��i�Q���	�X��q��'��v�kj��4�������777���
:~O�X��}����\�5�hCj�Tyyy+�ݟ],Sƨ&7����_����r˖��Q�"��V��[��RV���p{�+�Z�­���*1���o��7������n��ɀ�M������8ރ����1m�����G&3DӁL¥ѭof�����!r�R�F�#㳟�lܿ�Ж���Rz9�����2��`�Y�=�LX�~0�"2��	���~+a�Ԍ_o׋*
	�+��b,L�H2	ᬢ�(ҫ���Q�k�h@�9p�9:7t���?~����a�A�㊊*�XA�P�m�t!�~�7�c�����蝨J�}���%%�����-|��is&�%ÚJ8�`�O�|0R��o}����m����պ�ZD�J}]I���F�Rȭ�{���&%�Dz)K��vU	�Ⱦ��F��gE��*�v�u�z-hgNf	���v�m�d����%"�Ù]��&F��1����6���m��ͤ�:RYY�#��r޼+^��׾�C�F�V`|��w�;���
:�Rv�FPvS��C��]�>RX�U�����0�}�iN��1*���_/���~6m�损���x܍��>�[��0i��6c������N�}�n��طv�j�m\�י��Ϗ+.�O�z4��D�d��)�:k�u�����h���p[���=���L	�%>"0�#t�y��c߆�Nc9u������t6L�η�qȈ]U��5�QH�M�8��p4�~���`�0q'�BL�3c�Lv�,�r%ft�L����#H�7�B�{��3f̰�� �*��P���N~���ڀϿh0<8�v��{�֭'|���R?���������U�N�~� m׿|�rt�ʍu����'���*>p�@Ž���44^a��t��}WM��������b튝��4[����8��ɷ���294��Q�?pOY$��ɖ&�~�䢟lK�?���w�:S ݈��s��$��m�B
d�3�~�+��g ׈�+�%�w0�{�Y}�����,x������b4�g����Fj�9�F.�|-�p���Q�x�m�[�ms��	=�g�80��45�֭���Ǣ}��\w���Ƣ����P X==�tD&�����\y��G��r��UUU���|�	W˯~~ف�������UM���m �쏧��Y:��M��yA���%J��x
S:Q�M+��G((�8�q�n�W~��_�~�g�c�u��y��ɴ�&�Y�-6���={Ei��B�ftt��%f�4��ޞ~�5�|�c�ɳJD����pqN5�����.��^v �������D��� �A����#9 ���Uܐ@��M��SiO������i�L$⧢]�����������C����;wn�0aұ�7�р���r%�J x��.�S�N�������ɓ�������B��'�u.����а���ZJf]�и�~�`�[�E���l���9�]�e�-�N̥gC�q�a��c�HH$�"w��X"kY��_�J����A<X�ܛx�4�����,)�c�,��s@٥�J��Ne�"B&���������O�������x�h���}�ߜG��:�2:��91���,r��B���\��P���Z�DnΊfuT�0|z ����ݻg�]�O_��x'UW��ɻv�4��ee�{n����-^�d�i�N�ׄz��з��_�������t�β��2$���Aͻ~�����׿�M����"���#47���ͅ6��QS��قS���A3�4�DDd�~���ڝ|�1�ۄ!OY�l�.�(+��J+�
b�#]���t�*x]]�e��*: �x����m��e<f�Lr8���B����Kdu�vx���L���jll�F�tw���f��4ϴa���o�i����!���#����#^��HA��]UY�ZQ]�wժU����1 �U�?��o_X��H�w���ww�]�F/K��3L�h�Uj���{�zj<��:sAH&#EYk	��}i[t��O�Ł���b��ι�lwQ0k����R��p*��t�"�,�>�j�5���A�����n��Zں7o�eK)�d��;�)YQQv��{�����;Ｙe,�駟<x�Nj�)t�����Fv�3�E۲�	�Z�V�,�:�b���a��-%g��������_��~�OS��o�|d(�D7�I5AbܚU�#K%���@p��+^��%ơ�x/m�����ܶͳ�G��tb����o*�yBb�1�w��W������[��ڨ�hHW�-F2mhi�c�Hь9���Q <Vd�"7
gN���5k���:������YB|����1SJ9�a͉�Ѕ�Έ��t����"Lt@�LR��j}�=V89H�=V�Ʉfdh�-��̣�JjrECOvkJ�}��2���Gi�R��ėL�ؚ�?r�����q[��媳f����$�IXQ��ە�x�2�,=�v�;Nw�}�3��w��ֲP����������ʪ�}�S��Ј8PCSa��b�k�&����D�Ν�*��������K�gCL�����n�VР��	�~m����������\���d��[��bK�e�kԕK]@�=C�5��i@�mא����ʉ}d����:����4�ı�4�`�e����n)��o�/L���@!�B���ж�!R�����ߟ+�
R������d<q�������.���9����ۡ�v�Xb�,g����ٻ|��In�pK��)��w�����gY��,3��)�E��ʊj�n���/ejFW �ݽd��7�[��Y��w�.��"b�Y����ꅧ���z��sK��/�2IƆ�'�Zx�Ϳ�P3y�ߠ���]�ۇ�}�@�WCd���.U�VA�,�fw�����Ϟ\�n�}ԁ�@��x�\ݜ}��۝-D�ɬ���a@���5�
fb���` ��18p�7'�C���qN��.J�a��;>9��]U��]^�-�ir����bk10D�c�&��I�k���bn����45���P���7�km� �_׵��}�H`KUUe7�6�՝D(O�l;L�S�~�Μ&"������6Ϟ=oWW��ԩS�?���;��&���ģ�Yt�����d`)C/�-ٍi�┑%$���A�]8�k7�)8tXάͯ�#C�.g`��si&����f�%m��X89\<��)���Q{ �ؖ5gL�x��c+�l��IT�����.�*))��f���W_}���|�;�cx�x��I�;N�N�<I�1Bc'��Ѷ �r�,5�@�}��
���j���O�~�*|X�WrC'�~����6o޸����U�Dj��������e~�Ū��4��U��.�b�+W��N̞fT���̓�������_+0�%�����1O`0T[�j���~^1i�>m��?�)��1��X���/��B�p5��)�s��o۶m��q�Ɩ���������/u̎䂛��/܎<qg�6�sF��SAr�j8>���O@$�u4r����{���i#:C���u�=���cZ���v8J��KK˳�Q&C����x��zaǖ+�Ω�:�::��_BK�HO�^�]���~����	�J�
i�,,<��?;U^^:\PP��
�����ԩScc����ܴi�?��-8y�����Y��o?2-�O�6���bu�Drb:���s� I���K�bR��=[Z,�j�חC�����ɥ��)�|�?|���p�_���p�Zn(G��!?�Lϒ|���K�,3��{�#�d}�|�r89���������=W�v�-Z�h;��Cؾ}{`�[�����*��\3�a�M@y��v���,�}���k�����՛o���g?�9��𨹹9�s�ۓ���>|�N��f�	W�<�@:u:���/�YR\�c���/.�Ն�W�?*>��i��n�����ߟٵ�����[��)��DO"�S}ٔ�Ӯ��巍;�i3?B4٤�`LdD�t[�ka�)��%B�(VS
�,H��ux���������`KK��Q�0� z�>��F�xst<����	\'3X���²UL���N��������3m˳<;O�k��Z���"?�l��Y?�D�u%'O�@���L��˩d<{���ʅ>�.څ7H��"a��8"p�Wo��f��9���.v�!�~���x]�_����������/�qGEEIXz�E�@�?��y^�'�F�����ٛt~���kcc�����v�,����Pۇ�D�"���"��k!]c?�f0B.!O_w���w_U4�hf��i#]�Ieʈ�TQ�R;\.���=�	�,6לZBْ�`��E�+�[�.�l��Q�}aU�v�3�Q����l+���}va����!�L�a��C��V�O�$�db���C\kM����Ρ�<����t�^����@MM�.z��gh՜9sz>��O�����O��ɽ�=��5^ӬJ�#��|p�=� %b8	(����tR�<s��>���sFn��ٻwo�C=4mǎmK��N�H7��QU���;-� ��T����M�,z}�ܹoN�;��	�~�������+/��ڻ�EiqK���0�J�AC�*���TӲe�,��w>zC�.��d�R^�L�e$3%��OYn�9�?p�رW~���u��}���۩�m�g�C�gg�,jd+
:^���N��<\ˊ$tPp�p�2N��fx�>��}���LR�� ���]V<��;M9w�+��[��x��x���	3v�?�����YIƒi�NXǆ���ck��v����gI�\�)Z/u�x+PR�5Z�q���vZ����;���z�N��v%q�����'x3���4�?�)������(]c�|����M��Em�Uɤ�M|�T� �Δ��5�y��)�.��Nj� �/@���h}7�5H��8�T|-�:��XC��� -ax<��6bA:mK��ҳ�E���c�#���>��ʕ-��A��%H�Z����m��Ǌ�(<;c��t�	��\r���{�ݶ����M"3I��S4Ax������ӷ����?m�b˖-E�o����+�-����=���3ˁpCq&f�"4�ˊ�'&	��N��f���gՊuN������.���.��
�R(������w�,))�p�mKV_s�U[�ꦴ�g��e�����"�r����(J��>��C��=q��e�Uu���C�6u�?�ʸ4�Hr�1�z�LӜQYn�&M���s��>۹jժ殮����g6u���
�gW<˵ɂ9b0�\3���R����6�e��9|���<�g��vC� �$��ښ|�r�+K��E�F����d�#Wi�+�:`��a�Z��V�2��{�14O�S}��κ|�V����A!�께�Dt� �2DH���oC����ണ��&�	���r���I�C�ieP��W'rci���ј�$�?�![/������+|�p:	��3�s"�tjD4�n�.l��-u����r�)��`���˶�f+�C��ӕuA�.��z|�&6|�|�;���9CDj�E��?�}��'`mc�o���p��`�z�?�;�*��b��
�t�e�e5p�� ����&Ԇ=�Ph��ŋ�ig9����<4G�6W����ǻ��rA"��1���Ô>~��ms��[�bŲm4�����_}�����+M��>�7���Q��Ti��?L�r�O�o����5�]���9d&=~|hn��hF��Ȏ�u�p^�<C�7n|��_ܿgϞ�#u��1��`�����aG~�v��1�EG��D�r�a�5��3�e��i�}<ֱ�D���%2<����V�ػ��F�U�u��*Y'�;��XW�Y�Y��Be˅7˞�|y�3]���r�3.�bjg{S>��1L';.o��ODX���]�ϲ�9$7_�˿�6__n3�g�[vXDl�_�l��D6�ߵ#����d����eK�|��X��|?�5���cՑbˋ��փ���"c7�/׃����P|L��gK��C�LX#���;���^��O���{��^�������_~�j��ퟤk�R(�l�h�-OR�ⅉ�%I.�K�+厹s箝:u�Y��0�:����.�4����&9r����t���)�8q�+V\�v�̙�i�٧��z0��Z�ᅫ�V�۷�nc_&J����ᷗ�rメ�״��̶N��_}��q��9�J�F�	��%K�Ĩ#���㏷�Z��epp�3�\�L���<6�43b�-[P�� gf��� �.�A_�  ��������{�<@�>��d��p���3������|7֜�V����X��� �"���
a󉏜љ	�5yY�c�Ȥ�Od��cI&G�3=�(�B���91y`R�V
���k��u"�=[T��9#�����󶉠;��\X���C��8��o+[sK��$��LT�<�R�%��sd��0Qg��G�HY�:�A7L�{������4����Ƥ����?~�{K{zzo�kU�.A����Hn�~�U:���{XH���Mz�a��W_}\;9��������������h���y�ʈ��̈́����������x��mS�L���b�;�N�wY��o��RM���H���M�[p뭿��_�&�
]��'8���$���&˽"BG�

 ���s��������?`�ƍ��A�N�ˠ�@�m2�3H沼f�N�3j,	�61@���kTY��4����u�ۊ������	��L&�9��}%!����F!?
�(��o���z�H^9��u���`,��̕�r�Cy0��Uօ��V�x>�}x��xy[Y�Y'o�8v�`Qg ��#��-;�#�F[��lȚKScڪ%"r� ��c����\��]QrI�`��.�Abb��x�.��v��
{��e]�l�a���r�;�1��4�>�v����/������ݚ6�s#=���;w��8��$:o�	�e��������Y�qM��.�����â��Ύ�(�XrZ=�%w.[�lc}}}�\��MnL+��p�M�D�'�;��)OL��g��N�7n�?�X���ȑc��.���k��fgcc���fh�5���->���@"y=ͳ|�(�q��>����Xv�O�9g$�]�ao_F�|�a�����"QEmtHS��.�g-L��իW�~�g�>q��]��,�Ψ�e�ߝ%,��ٺ<���ekk(xP��A��&��1Xr�u*V%g����<�r�re��it�b��_!��[^xv
0��-"9�Zd���{�q���-BUUﲼȃ5��Sv����Hu�\�6c��vfm��J��Q&����)[�d�G=�r-[��v����I&��b�ߖ� �.v�ʚ
��,������W����ʓ�U#�d&�؎�S֪9��'d***����tz����=��O}�ښo|�b�����E���?����S�X�=�m=�����\5��hK���L�"N�<im�\���D(T��̙3���c���&����@8|�<�1���f���^��
�>_oMո����7��TuL��`mCD"��fe~��e��G��%��^�?X(���VU�f�u��η`i�8�H&+S�?�1�GϸQ��HGJD&��Y((\`8�g���شi��-[�|����wR�^�'�pU�S�Y1GL�E#���#���@h�B3�\����`�A�6��ʝ!���v) ���L?�yQF�ёK9�,|ι�@�2#n&[Td�{�rc�+[d+��~&r�s=�b$�'#�'7��)g��U��o7>�|"%�+�G���K��ɵ�x��N����d�;�T���"�2���G#�a}�в����a��հ�`a"dGt�\Ulqcb*[��7H�U��q�Dj�i�'h�7h?�,Y�d������� "��<k��}QTX���}Op�����|6x�L���^ :>@�>��EM_�pἍ������"7l�!RS}������H,��Dj� ��EE��Ljx��؞������"|N-fK�o�S�M:�jpQJxIS3�#<nG�/Y�+�`a�v��;UT虾N}�0�4=Wn�Li�L,��$�\��(�",]�t���_y啶g�}��رcw��3\j��q�5�x�@ɳh�TȑK<X�bPt|\]�-C��@�É�0X���� &σ�<8����r�7�h�[U�s0���0˖�3�[��[�p�|����/n�Hr��y��)�ұ��[���e� o��ȯ�͟��'C2A�;���L���ͮ˟�����-�Vv��ņ]P|��P���>�O���Ä�	[k`)�s!��xar���p�j�[դ�Dxw7������:u����総��P��e��~�o]���m#G��%��H$�nj$�knnӦM�蚘Ԗ�&LxmΜ9g1���xOr�����L<y�h�7௏F���8�9�N.SR:\YU����j���A|Vu4��V���죷��s��ƛ�BO&�SG4w8�r�8m�_k��U��{cr�0FF��.�O��0�I�q�!�
��ǂ������k�����W_���$=ӓ���3�|�TLr�;���ؗ] ��?���5���'�![p�;lّ�y��i<`ʖ~/Zew��>��L<0���f1���'-��F&)��5"��L�@"9A�ܶ�*o���Ǔ�3�*�-x}�t��#N�{�1���$H������F�;�(�>���H;&��{9�M�`��E��b�^,qB���Y��-����uhk�>��i,���^.����I*i�H�?EǱ�ƻՕ���~���m����5kָ_}����z�""W���}�v(���a��5>z��E
aA�{�������k.���\im�"7 5İ�mmm��T⪮���鱨uyt���Ё�T*�UX\����<)Di�|���Z^�zt�'�;N�]�G��N%��nbXw��U�kg̙���i�O��)��wJ˸��J0��+m&�.Q�,7
�(�@�끅���?�e˖;��Y^TTT><<��:T ��e��<����NtbLj�sT��A����4G��`*ko�(>�����F��O���3�7'�������G��P�E�2!x/1�����\e�vV[x=#����!���t��<�m�5F��l���<��ێ-~6M�ЫȢ`��s٭���d{r=�G������\~%�MU�u?ّa.�te$�����d��+#m�@�"6�������u�����Ϻ�t4������������y����X7'��q�e�t�����~z�w,�äNfbdj>VYY�����{��y��d>�R�ǎ���fq*_lf��2���о���-����b�!
h�����{p�������Y�q]��}�]\�
��.�e�����?;��n�W+��0]��.�n3	Q;�E��.8V�z柾�E;^}���w���).�N��2���̃����$�.2�O�f�����Gg�Y6|����L�<K�-A�eu�)�]�y�/��� c��B�\�Mv�v��[s\ZrT��[�Ɉl9�k���q��E�d7��l��m8��-X����]�<#i�u�L���#�$��Ϥ5��>a��eZ��I�\�kb8�"B���.�f�y�C���>��}��e�,E8F�~B��d]:W������{�^�yΜ9{�򕯀�_���ň��חlڶ鮡������8��Юra[vIM�81���N���sKK��;*B�_s�5�m;w{��y�s`b8<89�L��uW-�����}��YZZ��%O�3��N�k^k*(*�����ɔ�,��d
�Ԍ�E��%o�Ob�����s���&�nP���L�V������((| �1���U�+��Y�i��[��[��\ր��'�ʊ�q,:0���䋑g��S�����9�������d�«3s�z���D%��Z� Tv�Ƀ�l!0�B6G�֑����'#,?.mĀ�_D�L���L&�6r�!ٝ�ߥ�\��l�a]����"ڻ���$�ɇ�Ȫ��D���s���_/Y�-�}�ߕ��yc,�ŏKj���b�ϱ�+�����2�qG��G�?���Bm�v)Zz阚��WTT<?mڴC_���,K�}��'.V�=���+z{��.���pm�bj]K�K$�I���I�+¾a�A�b;D�9mk�uܺp��'�-[x^R��O�l�'�`�����c��E/C}�&�.a�C-B)�;TZ?n�,�Pw���:�����|F�c�]�fw��E~������-He��+�t����H�

c ���Q�v^}���W׬���ڵ�\�E&PD�Lʶx=v"@+�͂ݚ= ,����Zz���2)��"YUx&����5���8Q6֠��G��P}�4!�������bM$aQ��[Rc��Ȋce�k2���V�u�L.�0��	�מ�r��\o	�a�����&ߵ�d���L��&���z�Bd�'郕Z.3�ׇ�r�9rdW"SY�#[i�y~��h��1+�m���A9Sl+MNG����.��I�|��Be���m��Zh�/ѽ�̹���ַ�A߸����Ŏ�omnضcǝ�hD�U�ˁ�x��5B%p��ul�����|��~��>KD<{�l�2�k�v{��}eɒ%��s9}&���Kz�[��E;
|G���na[2�ɟ�v�����t�@uM����xYݤV�߯T��=-��\�c�+�.-ԙ1�I]K�].��z��"i%�;O�f��͎r����EK��zc����9���ֶE�Lf��I��ј��5��hAa�m�%�������n�:Ea[!R�ܼI&<�l��08ꥰ�~���x$�ɑ�;3�R�������pe������[������=���!��+&|l�� !W����3�J������2��B���������l��Z�wr��k��β��� �� ��>�9��50�^.`)�����^9k6���Qy\������Aǐ����wh�����X�p�N"7aT�����-.�_���ч~�93����e��b}d�&�A�.e�g���e�������H�&Im���k�]5cƌ�6�w74L�:0T)�j�TwT������t�{���)	�B���u�v�U�
uu"���23)���߫�4����[$� km={]6lصvݺ����s�鮮��`��&o�x"�|~+↉k#�	{�dr�5��͉j���t�\��&>|��+G���f�#�,��0d���!��X��p;z"���9a�`9��]�3���$'�d0c���8̙-6 [vd�
'X�������!�~�QA�9��L(���e�\{�ޑI�lIa�U~�_[�p��?�6`��$�>�ּ��ӊ��1�E,Y�,k��RC��IP�w����7VVV��>}��o|���%�|�'}t��֓�Ȥӕ�ڰ�κ]#��d�������������aO���>��<o��N�&����Ŧ��{RG���t�\ZQ�ZTV�����E;�QZ�f3�v�?�r���h��{Қ�+�0��\}�����Z�f�;n,���5�X�ʲǃ���g�I�T���!5<h�ˑJ�`�g�l]����L89�	�J�œt�+�Dg��Q�c�����3�u˿��W֐���s�0X���]dwkkXD�v�9�[�d�5���ڿ��(��1yɷP���Z�k�9h���m��k9�w��2��-4qK\�$V���l)������Ӻ��~7�/o���n����?��χ1�~����ݵ�����;v����1�~t���#ϰ���F<��R���wQj�5W_}���γl��<� ����q���_�3�k+�*��K��:_~�M�����t$KM���J��>_=D�K��+\�hҴ�o1[~�r�5��{��]�w}r`phv"���	�=OhV��1�L=������UnV�k"�����F���̛�~�בg���N��ͦ�灟I���)@�Z�.2�/62�w}' �; K�s�]]��0W?+W��������$g鱉S:[ނ�.��Ax��㒬T�^vw1�6/[kda4޳���ܑ�9���5�n�������m�HĲ�O��Ḙ��w�M����c���h�mDz_���ۻdɒ���v[^���[\�صkWɋ/�tG"��>ed�.����\��]�y���h�����}�B��޻'O����˗��:���܀Mvv���v��oS���jk�VTU���]?����j�;�6�����̚��%e�����hP((\DhҚ@rNn3͎yo��y��o/8v���'���fhx����B?
V�i�\g 7�ylF�g ��v�:Wy%G�v�)�:�b����?W�0s�yd�#[N�+��-�~>������u�<�#��������/�p��.�*#[�d���ؖ�3���������d�d������t����5U �f���:�������d�C�1�9A�q���Vmm�Ɖ'����gΜyA�G�m<��o�vM{��Ϲ��*�H�	j޺g���l�>���<ɠ�����ʕ+�j �zT�hl��;Ʒ���m2��)TVv����w_�FME�(D]ݍ�tL{��#v�)*f��'�(

!�.�VzVOoٲe�m�^i>�ε�m��M����9}NTO�f���-cds�p�A|dN�0�39W��9��`�À�� rX���p�<,T�Ů���V�Z��9J"2)ʞ�q�B�m�I.��C�����]�4g����2L��D��KR��.3�\�)d�䂔����ĆCѱ.��g�[W��Y#�km��mMbD��,�t��c�p��8���v� ����n�3���3
�9��G�^�a���ij�E�<L@-m��m��rۼ+���v2A��$�����@���7��\Q���g���|�Hen�(�h����y P�25ܨ�kR8��Eon��y'��h@��.r83�6zn;����֖;ٷ{��mm�W����4��:;��-9KD.��\z�-��`Ɲ'���S�c��I��7� p^+�JOO6�Gvkq�s�j˄G�~ r���.���|��MnF
��m����E��Q����N���D/�.&>r�q@��m������Rp3ɖ-v	�Ƞ9򫦦&�bw;���ȑRL��kϮ����zo���1'��>z=B��}�ĉ'M����+��?~L��	�ٳ�r�k�ZImh��о���rP�w���W���H+�	���>�����ܹs�\(O˨"7���u����j��<*n������E��fb�(.�14�~`��ӝ7���~�PP��t`���8�s蝃>�k׮�\���l|����i� ��3k�G��r�=���(���@�3�N�57l�;e��$�>�B���ph6k_X�*�8���ï�@���ɍ��[�΄kz�왏����욓�a@�`�%[��U&z�o;�%s{c� �U��l9�k�, F���p4�6�{c?�a1[|�b�XG.� G[���$�������)//�Z__�qѢEG�uX���DG���G�mmm���Wa���κ�kJ�g�?IG(�ף�v��{
���n��K�Ƹ?B�P����D*7��˅:�QCn�atDE�<���T2�<TR�YS3��M�&"� �8SG98�Gӆ��>��K�����l�X[[�+{�{��[�����6������#���C���2�#}��	��҉�#yg���ʷi��K ��\%�Lz�]6Lv��Y��Y�kH��2����2�Q^��kw�9�[.�)�&rR=YC��H#&Ol���|ȸmpn /8'~���a=v�9����XL�W���ꒅ�r۲+�-M��Ei��}��Զ�'�#"�άY�:�N����ф��7��ܳ�.j�&j+]ֲ��kf�+���Q���<y�*�p��	k\ST�v
��.����/�\��Fb�
r���GO�?��V�JC;'O�����Wǂ�FFA�����?���S��O((\���|�?u�78p�|ǎ�>|��g�`]'�QI��7�1i��59��=�9B�����Zx�PpΣ#kJ�u�d1�Zs��,���#�k#C�}�\i�u��r;� ga�E� �2���+^�H7�<���!�L:d�M~�XJ�6 HvO��4+�w	���2�}AZ�f��l=b���%�%�'�_�$�]���hG;dܗ=&���~.�}7d�v��s���&L�:}��=�g�$B3��N�7o�~�W����p�:��
L�����bK��91�g��d���^�d%�����g�V��N�7���k7k�\�'7pE���=~䝯P�^,�466�gAAɺ�Fl +!�[?F{��RPVrD"��}���ٺu��������*�"�O�N��?":�	��6�h�|1�&R�Z9C1��$�i ]�GF&%�k�Lb`@��ȳ_��@��Wdf��,A�&t,9LJإ���u?h.���
R�o-b�����[ܞ��-3<�I9bF��aKg��povgqrR=&F.�6v�9m��ߋ�w��]���{���illl�?~7��/� :�������~v�#Gory<%fڰ�#H9�[ppmQ�kڴi���ò�! ���`�(���A�Ϙ1�{[.(��ņ��䞞��q��[<>O礆���yk,�n���ñD���+(H��|9����>~��Z^9|�`���������4р[C����EuiK��hL1h� n�z.�[�
Οɢ[y��g��6�|�)�Iޖ��QF@>�y/ѱid]-#,5���a��bf޷���=�	��ɉ�q�����=v'����uH�8,[�d�|l�K0I��g��p08:��t"n��1:�!�K[��뷌?~#�C��I'����J��訟��'�w���j�Ɉft�����aٲ���C�Yd�ݤ(���rȲܔ��f�84s��?е:9��#7h�ӧO�8u���.�~3��'N��EQQ��Jl���ܗHDƅca
��p8n+<�ǅ������k�@�<xU{{����x��FF1�� n1��h���X��L�d11o���i����9t��1��r�H��u��!�b#kJL#="����dR�,& ��($>/�I�&e�E�-�	gt��$�%D�xem�a�L~�"9i�_��;_�Ġϡ�0����k�ޟ��O1;:nܸ��f��K�$�TWWG���X�zu�Ʒ�ߛ�Ǘ~���UVAҥ�8\�3fX�p��Wp��j�kd騘��+���\s͛�%��������*��}٭��A��he����ޤF��u����ܓI��D�PPP��p�*�����|���u�L������5k�o`V2���>��4ܦ�Ӓ�+ ���O��]�@w�d����kn�Ƀ �m,ב�ǆ���Y��.jd	�P�� �Y�qs�)��>��<xq�m���J�����ے��li�&�F�n&��d���A��tޣ�PhCC�>���r���6\YY�T.���m۶��_�00�������X4-�����n $d�$����BX��E���ŋ�Z�h�y+���pA�M[[[iOOח���ʒ��}�5U�.-�x�b��� ڷo���jH��z�n̴3�8|�/���NK��C-3�;�g��������D"D�\�V�9�j���$w w�2��z�wYv ٵ�/8�39�9ߪ![Lx[& ����n���a��̎��'��� ��ٙ=������e�|����|Q����n||� 8�\"�p3�xE-'�,�뮡��`{QQ���ښ����{fΜ�5y���4�B��QQNg����>��sK�?�%�^���s���vU�$>|���Od����=;*Nd�^;>~��ǉ�M�３j����cI3�ϕ����P��@�x�fW!�(��ܕ�FA�#@z�`���w�ɷv��<q�DQWW�����Y���S�i`�D����._4�p�.�|u{�AWآd�rgy�A����8�����}�Շ�����������xg�H@k��&�%������AEv�q�?�����Z��	����ed��֕�^��&Xe2�����ޟ��(?J��!"0-��2t���Ƹ�`L $�������7���/�Ѕ�A��}�6ҖU�]�~�׉�CT��D�:s��iZ{�`IL[��Mz�����ᦛnz�B�9�+�A⠎���d⦲��S������͎���(((�;8�],H��A������e%�zZ��i���S��p=�0kh�Rꀽ�x�J�n~S4({�i��B�+ ��Ϸp �Ȍ��=�E���X����ي�D#?Kr�o8픝���Iv����]��,�f�?r�?�v�+1���@  7S{UU����ң���?E��'N�WWW�4�j:�X��3%��}��T�Z��A�Rae�u/�D*���@r��Z�P�<�cǎY�m R����n�C���d"I�Ė<�hѢ~1�p�-7��Tf\yE�����������QPP�s��X�4֢s=L�~��!{{{�6KN�:��뻌�o���H�d�K�S.����0< <v�a�4���roy�d�6aq�ɸr��R��E�����ɍL�dKo�<犃�q��"�d�G�䰐7_ă�W0�a��.˵��e@d"�ް��t��]�E��Dĥ����dEEE/�?XRR2<c���%�0ؼys��~���h=y�3D:����v�J�'�1=>o�]�{�����s�l�
z�������� b�B��"��+��y%7԰Qj��J�o`46������U�n�!�n�������ttt�J�=ZC�g|��D"5.�LT���D"Y�ɤ�il/��?@���e3$9����KX�i�L<X��ODdݍ���31�*�2�ב&3�؏-H�@YQw�T��k	���4��x=}��w�w�n���u�B�'�k�O��ֶ���;y��az�766�T>z /�<��ĉ����za��H;+�xX�p_�]��H���Y���JB�r�S:�����Ǯ��׮�����L8�䦦�&B�
�SPP8op�aA'�G}�qzu�>}�}��O8.���,������bhh�&�USGϯe�T��02�4@x=ܺ���]��!�<����#�`59�^��$<��ɢ�� �	�u1�.�Ö�l����aA���=LJӵ$@�=�}�N��🢁�^�%%����q�K���啃�'׆i L�7β�)23z��/N9x����z^N����r ᢕp�qM"J
�a���\P��Ֆ���O =��c�i	P�{˼y�^Z�|���8�bEl.$��,,��~�M�E���۷�Dp|��i0�������Zʨ�/�����b"<��d�"�N����P��M���.�M�a-D�<�A_�$�M������D���~�rƸi�l�(ٟ���ٖ*"2����N��bE���5-�r��t*�v�<I��`������@o�0�QPP��y{KK˺}>�@EEh���x���,^^^�1c��.2D���`�{��{����qC2�,b�X�E�X4�������rU!�4t9����D�{���\�ti�h&��������3x� ή�I8i�Л���D\���.�ٺ�q�'���D"OO�0D��@*+@("C�t:H��T*W��02����dO&�v�������NjXs4�@O0��z�谶X�䊡�%\.w������DVb��'A��Xiii�f�P(4L�'��`�L��!C�SY`."�_�>��g>�D��
�q	d��^��5UUU����a��Q����[��%
�Nxx/�GO�q�oM�4iTG�)r�������������,�����͎����O���АN��,N$b��h.WBK&]DjZ*��<��E��o��":~��N.W(S^�����dL��DX��t��llL�xQ��K ۶m�����_��y�����#\N�,�"�`�`�A%��ޞl>DB�İ��+N����=��E���={v��P�FAAA�,@�R�P ���~0�؉#�J��#�'~䄏x���,�=gن�ٗ�>\X�S:#988�c�ܹ����{���@�EEn�(����o;����'�&R����)�?G�q�,N��8*46����k��i����ꏷ�v��E��1�={�_��[{{{n�z�!�H㢫���l�Ć0-�L,a��@�7¾!���\��I"��F/�X�b��i����"7





c����~�����_�x=u�%�#�F -��pAU�$�H������bRÕ�i�m���ٳ��;N�%�"7





cȭ���tƮ����x��!�6�g@Z@d����X���p"���ʬu����p<f�������o�y?m�c��((((((�1<����[�n�"�����dJ�pk�½\�].��ua���:��p2Xhh�NZ���;^�a�g�"7





co��V�C=�W���'|>�Kj~�(*����WXft������K���L@��̙���ŋO�1En�P7���V�v���!̚d"�YD�!2��a��h)|�e:��p�7 ��a)ZOSSӣ��sϑ���Q��1�7�xi���{���zg(��a�0��	O&���P���OI". -��ư"�@f�va!��)G{c�����Տ�q��ƚ�F�"7





��g���/׼�j՗�.�R���ȈBx=^���*�
�D$����w���uP�V��u\.W/��ԕW^�jڴiCbC��Q����k�\���{cUUUq�4�H,!�^;Q"�`�QAo�����»���Xp8*
���-r�u�@���Z"6��r�-�b�C��Q
Xl}���o~�����_!R��u$��I~���a���`������>y�:���%��֍J��<}����c%��A��Q�5k������_v���O�>�L%'t2��]*��&0a���3s��={�d���a��rcD"�V"E�q��kkk��"�"7





�O<�D�?���=}ݟ�����W�q�*�L����g�k��	�k�2�H��ӧ�}�zd��\�U�vE��m���bŊ����EEnF�~��гO=��hl�ۺ�O7twA�4�h"n寱�P	�=�S\b�������EEE���5�@h ,�z��!J�ٺx��Go����"�"7





��7o.�կ~u[Oo�W3�
".^X\�rJ��H'Xj\n�0������E/a�@pt�ml����.��I�'s��{t�ʕ�N����((((((�@<���`NG[�=��5���#�@b4���5���	�e'��	�0�������-2������`l�ݮ>���+V�XS__�QPPPPP�� �y��'����7�f�GA���5�`�IeҖ{�#��z��)**�փK
�X�)�	bӟH$��0��~���>�QPPPPP�� �ٵk�ķ6���Cᾕ�`aa*�Ҹ�Ծ����}��H$bYt ,������ME��h4:L�����_�r�-�D|2�"�"7





%/�~����֏���r"�G��0������;V���	����(&g)�u�D��{<�_M�:u߂�ly�?En.���^Z�zž�{�%R�H�ą�
 3YR�kB#��u��������\ ����RLx���js*
=6ujӦ/}�K-��QPPPPP�  �oݰa��V�CĦ���-6V��S�[":��ȋ���+�cbN5p��̘1k�����q1C������E[6o��dk�B"4�d,mM���h.���LX,�#lw���'p�b ��*(��9�N&�����cW�"�"7





�DT��>��oo��9��W=8<�!�����~�0�/\Pl���4Z��Ȗ���+��S��'�1L��'6�"7





���ڰaì�_z�s�Tf��pDKeL����zuy,댮�6�9"c��f=��gC���F����x<.�H�,Q1��&d$�(���ȍ������yD{{{���^�\wo�b"A�V 1aR��D*�˺���"c3�Ñ�����7�� �M�6��F���" %�����:x��m�T��H����0)�*�E��b���3��E�2!rB��������aq	@��� ���n�:sㆍw���z���/�!&+dK�"~��˖lK�Ơu;��ݴJ\\P�FAAAAA�<������_�|__��D"�O�Ӗx:��3X@L�.�EN�-6��(ƙ�-�ﭩ��}gŊiq	@��s"!x��ۏ9r���PV�,�aXv#��A�97�L��;�	��~���G������>q�@��s"!�u��-X��ͻ��ĸh4�ЗC��n&. 4���-7L��j#�_ d�Xm]��p������?}IDJ��((((((�C���5����w������� 6�A�!R�و�t�ܰHمe�L�[J�� 2Ir��%��[�P�����K�j(r������p�@$��/~q��#G?�C�Ġ��$����E0�Y���iY+��3X���ٵ�1�'C럠��8q��K�j(r������p w�o�1w���(�I��͚��Xa�.��n+2��95��������7jkk��{ｗD��En�2 >�rrº5k�i=qbF*�@&��hX�vbr#縱H�Cft�`GU���߁4�I�:[�n���������_\jP�FAAAAA�l#���O<x�z"Ű����(�|��l�9S$�����b�WX�`������F�?;o޼��B6�3A����5o�={Æ��E"�q�l������[���n&3�*c��G����a]'I�\<�L&�L�<��{�'|���K��((((((�%�u�����=�%R�CdG0qaK@�K�E/���r爎��������`*�H4���G>����^�V@��������7�|������E��1�d2)8��c]yW�>�a0�a��{e#xƤ��}>��.ܹ`������ȍ������Y ����뗼�f�'��xE*�ғNeo,�XL�Q*���a���Trd�lx= �b�yJ�~ޮ��x������ .e(r�������wԩS�._��ٯ�S�9�n�����t�!���^Z�}f�Chi�����ә�M\�a�lW����墨


�d2�����nѢE{/ewC���$�{��>��~r1?�g�G�+�LĂr���P����#"���bdd w���Wf͚���oN
En>
Ps�ߺ��L$�D6t���D:��ڸ�i������#�Ɍ�h�%v�[����p�DX�F����丱�D��VVV>��/�[Yml(r�������g�ȋ��ĉů���_���N1͌ni���,�b�n��B�9�$y�B�G$�c�v�����z�R���{⪫�:@�B��"7





&b}�qO=����ۯ R��"�H�Dd(.R3�`V��#4��!�шp{=�5�䴡�l=�aZ�5�%L��t�6��6Dn"�t�5䴹��B!En��(��5k�ؼqݭ}���X<��R	��W�rgú�J#�EQQ	�V��D*��q��/+��>f6jJΉ�Xn��P0|�;�8��Q#�ȍ������b�ڶm�C=���=]��XD�x\bʔI���N����â��Ktt����bh�_D�B�xEQq�pytKc��nYj�(��F�l�>��x<>��q���.\����)!F@���}���Ly�ч������S�Lq����X,"&M�(fϞ-�~����X��CQq��I��q��Q�7q��{�N�Io�DMq�����w���+**^�뮻"B�]P�FAAAAA������?޺}��7������F�~�[��f��IDF��/E���r�xDaQPL��$���DS��v�S�صS���"
���"�J�Y�uM�TJ���Τ��!֣[E1�ؤ��_XX��m��vL���En>�=Z�v͛7����ؠ�]��H���L+�����tҎnvHx<����4{�,�l�2q�5K��O�A4�kS� !��aa�:�~%Rc�>={��3g�T9m���((((((|@ �{ÆMW\q�䫮Z�۾}�hk?)��b�����ȍa���-�zQ����03+GMaA���,��α�ϯ��7���KTU�XI�	�̸]����V��'Ni[c�Uw�uW�PxO(r�������100P�N'�]�re]ˁ����7���*��8�"6^�wk�En��I$"O�t��}VR\,��).*�dB\�l�hok?�����U�Spe�����ܢ��oo���w��d��{B�� XmR�TS \����]��QVV*.���rE�*\T\ ���@C�1��@|��C���R���@O�H$�b��bɕ���u�ĐwP��VX"b��a�i3,��~v��y�;�OC�������X,r�if�m޼�
�l�墶����X�""��5�@l�ߦ��<�4TBd(dE<Ň�,-MoO�(Œ%KġC-��o@������O䆾K$�h4�qҤ�g���/�|�K_
�En�L���}+O������͡C��ɓ'���"�}��KcmL4�d��UO*� �cj�^PTVV���r�s{,b���D�֏��`��5c�x��5 Q�8Tf���4>�p�fUb�A����ڄ������ϴ���k�vwA�/j�W��	�E2>�W��(�i8ل�"��{�HJ�(/�e�x]n����^+�q,���jV���D ��T\K̴���{��fΜ��+�B�A���Ga$2pSO��%{w�ģa1c�TQQ^"�a+�A���v[.(!4K�L	��@�W���Z*
�����>�HFD$�DL$3)QTR"*�j��I��;ﴈ`Q1��)�k�++˟��{��^����ȍ������{�4M___ג���/�ٹc��֣���QW?N�<�p�Maj.+BJ�M�E��E&�E�E�4T!��Bڛ.�ɤH$���>*�>�O��.K��g�~$�3LMk�z\��7o�v��pP�FAAAAA�=04�3����G��y��!:���z+����j�^�Gd��0M�.�"0�)


-��[�2	184d%���H$j��z�R�}��q3cd&V755m���Utԇ�"7





g�i��������h�qǎ��{w�#�]����ֽ����f����ǳ0���DD"��M$@(/	R���׼�,)�%a�	2$A(�3�ͳO�L��6�]]�v��ί�G(o{<U���KwOWU?���;�s�j�B��34>>F�Dr@����O�w四�9��M���2�p�1ߚj�`�ju8����7���dP2���LӴR�4�a���(}�k_��&V,��!�   ����U������W�_�|�����LM��dY�Z�x����@������(�0���y_��� �p��t:��P���&Wl��:َ'W��}MS/ۖ��G������  �o��Q�~��vm��k׮}��=��������0��y�STl��x���d�qT�T�/����_��|�^!�r�e2��,9'&Z[[[��'�O���^�q�o	�  �7T*��5?s����ܸq�	_��y��<y}��j[�)��X�о(���.g��e�����uz=����z8��>�q(x�_�V������OO~�C�}�����_'�� �   ��������n��ŋ�����ѥE��?D��b��Η$�\���{l�b�GL��D��8�"��n(7��_�~O�uɴ3��Å�\6�\�{�g���7^~��n�8�w�p  @��^�:ӨV�p���W.]2����I2E�I)��1cp%2��r�E��_���qWm����R\�	��#Ӱe ⾛��j��{e�ַ^xᅛ�>�lD�;A�  �oԶ���Ξ;�z�K��89�MI���r���*��*8�*�'��yY��{=j6[*6��܆�����V�x_q?��������|�ÿ�?�=��O�;C� ����4��T�;/�={f�R�(�?y\Vm8��?��-�����Q����<o���\� �/�l��"�p�MW���-*�uȰ3$B�������lE���م7�����p  ��~�qpkg�s����v�277K���"��){mTyŸo������'dՆ�3�c�3m�(��w�Á��8dێ��$Z�t���|���sSSS6� �  x��@�_�{��7�;w�t��e��6\�15CGɣ(E��N|훛�y�0_��D�X�۾�-��:}p�uj�o��0�ER�t�����?����n  �%��Y��~����s��M7�M����O�ڃ`��^�&��R��r��w�0FI��@�'
y4��V��u��EAG��T�85??_%x�!�  �c�oG5�C+k��_�z��{+��9V&D�1��ĶR����~s0�*�����0���7�W>��`c;���-�?
Tո���`��+���  xL5
�F�Oj՝?z���._󞟟#��ɶuR)�����{m������нl6O��MM�P��Q�ӥZ��`�_�#(S���풪[�3�8U��i�]�PxC�W��%7  ����Q��}�^�~����鴛�SO}�,S%�TD��I�J�@�y;*�)��:w�r�"MO$7�Q"�N��&�d�GV\�	�W��xy�y��b���:)��f�srr�K�A� ��
GU�թv������}릱�0O�BVVj���j$oG1^�������(�.\ȗ�X'M��ލ(�����c^���`��/>�u7�~qqq���]7  �Xi6��f���{�w?s�����gg��f��l
z]rL�e�z>��M�Q"��y!&ߎ�-����<���(8���h�!�+7rD��(�""��+�rU���]�p  �>����������gμ9ǡ�ԇ��l�Adp��0hE�����J�t���˲φoG�A�`��n$��9�)���o��Q��5�G�B����{n  �Q�o���/^�|���7���8J��+����R(����5\�ID��.�K�r)&���AOC�[RQH�>�:�iP�� N�_d=�G���<7  �X����Zm�Oo޼�Ǘ.�ϗƋ49U&�[���ǐ��
��	��\r�Wnl+CA�O���b��;����NV��8R��a�ߌc����  y�a}O��[y���xn�ґ'DhQ��(M��12�p�aX�ʷ�H7-*�'�q��e)�"���;�jS��˹7�x���E��I�����}ϰ��ǎ�q�C�p  #oggm��[��ʝ�O����/���,�$��)�7\�)
�n�FE��95�2�+Ɂ~�z��@���ߤ�#(F�.���]��?l��ɑ#�Z�  ��4��]�t��۷n|���7����b̬g��Dr��(Je�L���}�nO�&O�������nˊ7�o���<�r9ٟ�$I����{i��M���  FV�����[O�[�Ϟ=3��r��4��M���ˊ�t�K���H�����l�^�X��t��^��Z���>Ǖ7�TUO)U��0�A�4}NQ���C� ��$B�����X�W��曯������DyL�c<y8�&�FU�5� �)?s5��lxw[�z]j�[��^r8��lx
q�$����8J_�m������{�  FS�S�ک|quu��\�d�L�.(^���E��n�^Rē&�q������)9�O�h����+6}l|9�/����c����a��UM��ɓO�c
�{�  F���ꝏTv+�=s����!33Sr���$��������{�"���"�X|U�?@ף4�d�M��"��Q���y9>��3���4I_�8�m��-�  )�;�R�X�V��z��['*��v�*��j��},+3�<�Ӈy_T&2�p���r���0�{�9ӦߑUn(��]T*?|����W='����l��=�p  #��Mowwfgg�K�o�|r�����4�r�<�ҹ�8�H��8��q"�`�^.[���*�'����
ro�9�2�%oX�܄LjE�E˰�{�x���� �  %��^�����ϝ�x:�dz�W&���R�$d��¡F�(I)I�I!]3�P(Ry�$���0�.7�P��Q����v���oWi���)��������yE9��Q� �  	|;����g��.�?�DmwGY:<O�lFĐ��XcȞ��X&5�M�F��T��Qs���ˎQ"����n��]��)�"2-W<�x�!�P��@m�^��?>z�h����p  C������T�Z�ʭ�k��|�^���R�Hn&#+5�C�O��(*M#L���}ʘ.yټ\����H)(����hP�ݡn�=��*rw��ɑa��$-���e�E���8�zt �  �(pv:�Oܽ{�gμ��O�r�\��V/4�r�M"�n�E��b�uól����O�>�E�i��ko�����'+��������l6{~nn��!7  0�DP���V?����/^��Vw��~��MC�,̕n"��?Fq"'
��\./������H^��a}�=6l�s�j�S���#R-��W
��)lj��  j���|�Z�ڵ�￷zG������tE�G�̲�#>n�Ex	�P^�Nb���MLL�kߪaP/��Q�8�p�ɸ�:YY�	�$�(=c橅���G�  �4��޾������?y��y�TW/�Q���y���Ã�zj� ���2�#�l&�Sd9��e0X�����&����"�����q�i��r��["8E��  J"xdVW�������ŋf�Qxqqq���8̏�*�$��x�7��%��M�8|�;�v�M�N��"شE����Lۢ���׋@�Y��i�)/��G�  �U��i�j/޼y����*�<q�,��&"n(�d����f0����}P��\����~Wγ�	�~0��0d[ٶ3��D	UM�`�Ω���
�#�  �N��o6[�{�׿�ԝ;w�'����x��)�X�Pu2[�MH��}��o�ˢ��irrR.Ŕ�Qr)f�|ߗ2#�ic۔�
)��a(���5J�Sf�<��G�  �4M�۷/�s_��pb�Ȣ2??O�f�P(P��hcc�՚��0M�HQz�T�����&�A�W,��n�)}�J�ee�Ë1� m���J13����\����p  C��on��o�l�����h��m�*
y�K�ؘ%�{WEp�I��Wq�q��͑�q9�P��2���A���� ˴�g�F��T�$z�5�SsG��0��чp  C��:�O�q��e�f�O�1����Q�ѐ���x���x���
�.���ǆoG"�Dl:Mj��z�ˡ~1��E����&M�DX�U�;�i����� �  n"��^_h�{�VUuB�����E�O�v����)CV���l,��*�&D��Q�rx���5�FS���p����QT�?�����}nn�E0n  `X(��_���ǣ8��W!tZm���V�*��M'>fj�[�yYf�s�L+C�l^��wz����j�j5�)�bl궼��q�8���Κ�sjvvv�`h �  ��0{���(�ƣ8P�B�af�7�
Lw0�O7mY���ܤn�O�G���+�P��ypt���`c�yn�L��$U�4����4�N+܍C�  �B�V���;����?s��[�+��t�}Vxp���Ŀ�2�DQBq�R�Z�;w�P��h|�H���đ�Ǖ�te�Q53�w�u�2,�ο--��vԐA� ���I�p�Q8̤a,Y�c�A�C���+ݝ�\��;.�8&M�hss��/:-,��N�J�N��ǐ�dȰ�tn"�L3sAS�S����7�n  `(
~���� � �D����&�8�lV^��pp	Cn���a>��Uח��nj����q��qrܴ�&��"��������<E0tn  `HL�M}k%����i�$D�L��2�.�i�lnp[�9�8�GSr���f�M!'5�1sق\��I�����k����T*u��  ��+d���J3"��"����*�j*C
Zrr���9�p�f�V�n��u\��dl�(���y��KKKwQ�^7  0x2p�Ѹ���+����%�lH�����$��T��vF�4��}GVp��]��=�.7'���(���B�,vG7�  �\���y���x���D�Ħ.e뤩�P��p÷�xj1We���_�g~8���*]3Tn�Ԇ���eL﵉��6�PC� �������_Lf����:��F'�41�C�J�-|���
ٖ#�WpT%�$�����0��GӌP������`qѿG0�n  `�LMMuvvv~�h�)�����i�8ģ���d��7Wh8�p%��L�҃�U2�Wx"EU������T�C�7n  `���V�V����˝�Ս?���㤨�8���LۑGO"����QUK��CWs<�M�0Z�����E�33�z#�  �R�X��i�^�������nﳶm/��isӰ�^�R{0��麞����v�iY��������%7  0�E�E�9S(�o//_�e���|��O� s0
����&�W5UK�$I�8��tC��d�:N��'�|rW���C�  ��^0��*έ[�.m�n<t��D�yJ�IJ'%%QU�oA�X���m�o��{�رc-���p  #aos��9�ׯ_���������iZ"�=�<���neii)Đ�хp  #eo _k���   ��   )7   0Rn   `� �   �HA�  ���p   #�   F
�   ��   )�z��gApˈ    IEND�B`�PK
     eO�Z��X��&  �&  /   images/9c69fbd4-c376-47ca-8b4c-793dd402431a.png�PNG

   IHDR   d   M   PA��   	pHYs  �  ��+  &�IDATx��|XTW���^�`�4i6P1�]�gEQ� `CEcԈ�%�h�c��(�h�%�XЀ
�� �O��_���o�/��D�,��a�9e�k��]{�3L������������������������������� �.]��Ap�HTTV�B^�,+ 	ll@ ��zw�'9��e��дiS��� �._��7BXx8dfeBYy9h5�&9�Z=�Tj(,z	�%��]��	\�\���������a���'���+�.à�C �o�h4�'�����K��3��)��sK*(TJ���o���[���c$F���Σ7d���|^GG��Ԅ�Q������Zpx�BC�Ӫ�lV���gs8O��v3f%���Kw���79x��΄A�!�c;�l����Jii���tHIY����
/�
F���b1�!'I��}Z�-f���d2�h�z=M&0�f�X(������i@cЁ�d ��6�U��������«_-�� �Wܿ���� '&Bt��ԩ�{��
2�֬�Z�/^��_�11�lllz���+���*���xR�4J�Z��h��C��7�1��j�#�3�j��jBPh#��l19�z��dq�X�<�l6K��rZ�16U��a7�\�A>�wrϞ=�.�ΐ~�,Y��K�!��6�^��� d�w����P�A(+-���Ҧ�X�TF��SUU՞Fc���ժTz�!����kg'y�,u.ܵ{K%bnР�;8�� `1[0�=
[�[ûrᖛR�����d��`��Kp��	��Xt[:@��h
���J����l�lw}��،�}c�((,���1N)���@�.�`����d,�Q@N�<	Ǐ��������!�mk?��iL��GC,&�QI���k���/��� 	�]�~%/0�9�x<x�<���cGF�u��;\,	�\�H�P��j���b���
8��;�Ɛ �\������E�����耹�l��g&p8�	���8;;]�������3�'KZ�n�eU���b�� 4$&&&��1�G 1�����ŀ�b�ê���dm���kjQa���,4��a�m.s؜=���O�K���3HcC�
u�N����O=��d�0br��[c5��Ӏ���+�r�f@�¨����|c1���H'y�J9�'��&��d�ف.3�+cW5	���p��v�ؑ��^����`䨑0���вe�?56; �.\���" �ys�ة���{zx�,++�ǜa��o5W1���b�]����2��C/| m۵��e{��QVV����&�p����� 0���x;�V�3-`�' 9�V��@1[��<���: �����ނ�C�Y�3l�K#�W���#�ˉ
l"�z}���4��b�߶=5�e��P�E��%K`�ܹo=> Z��m;�C���;��;w��{>����I&��I�сN�{��������˗K��{������D�Ojj��a2)�J�F#��>�'��5��ht
�7�����(�0)fs�j:�!����	)�.a���I0�@�Q��oЛ	�%f��m0� *0J�z����u:'[[�q_lÆ>�	�/7.������?��_C�M�o$77�̙ФIc�? ���W�t� ��
J�Z���
�(�����xk��pi�ڙ�a,{�,/�(%�B��2+�ǧ���bfQQ���)@��`0�7�Dj���d��֢�O��=�$#�����+����$j��	:B'L��KKt���#(Z�h��\giUu�Vo�uC����ӛ��f!U�,��1���$uJ(*.�6q�ҥ'z����?�^|�������~m�t��n
;�A梜�G3p ��C���	�W��
�6�~b�7<�]�]�r%U��z���k�L&��X/�cKhJ��#�Ӑ�x8ЦL���{����{���҈����$�	Z����p�@.S��S�c`K1JJ�{�߿��SǮMUJ�p�F'ٺ��j�ѸU*�L��ʚK;}�T_ԏ���H	 �Cr"	�%����n�����&mݸq�Q�`ڴ�o<^���7�,�FĎ 77g���nS(U]�x2��i������о`��|�>
�z{�<��Ѩu�ji]�Fw�&�,[BQ:��n0�
;��Ao�^�(3z K���W�ATT�����&c��Y|2y
���C��Ci���u�BQ;	��S[[��b5olָK��t�H$��_�߱c�o~���<|=�u�I�++�4k֔�*nE�N��'��/I3� ���?��Ȃ��aܸqp��Iprr	�v��~�Q��r��*�c3F&���9\,>z����^���;�JK�T��jͨ���X�
K�3�t!�O�D�S:�n	�ow?��D gϞ��BBB��у��G��~�׮]K�O�:F���q.��G��}�e�<���L&_#	������%.vv������>��dgg�iҤI1b)b	 D�?x�fT]K�Z���r���g�App02�����������/ �op��t��yx�f�8�V���)-�[�x� [�sf&��6G�0D�B?�![�*�J��ѧs�N����C��({@$U�Y��M���q�.hu2 �"-ZQ����Q���kp��� ���;v�dEG��q�ж%����ݐ:����R)+������sߢ��N�� FZ����'O�@�F�@�R�4���������~�����:�9 s�̡$_��p�;|\T��0V�b��b��铞��n����
����Bǎ����[Ԁ�^�Qi�4j�#ch�������L�����!������[7	s���̊+������G�M��|��_�p�XRR2��ӫH�ҬA1����͋x����Mh8��oyhH;?.���Q���0�_:�����*�7���v�v������w�^6t�o����x�W�ł��Q&`��T]UyĨ7ۡ��b�W-�>��.a��+`ذ�0v�Xx�"�74��L&��bѦӭH�>�������|pqv����W&��b!HQÞ=;��Llr�7�{���w�B�v��Ν�k��r�Z��H��j�Noo����rSX�^ u��|��igz�N���5���p�J�l�eeй3g6�(;[~������K�q���������p��q��������Ja!fg���B�hHUU��n�{��؉#�F��ԩ����k�W��O��K�+���ˣǏ-E��Ә����%���J	O�{��iй�2�t�
�������뜉�d����EF�a^۶Ap�����n�L^{��a��d�A���(�����]V^�]o4�����(a��ٿ~��g���:�;��ٳ��e#z�#���eA��`��DM�XZZv<j@<�~q�8�&���EPTR�c�7+/-�H�n�ް�E�@�ʊ�Ta��`g�8:&bz/ �66<X�f���k����0xp4����k�R�/��,.�w1#��Ŗ-������k��*�����O�؀I?Y�3��
�z��v�J�?s�Ӟ����\��#��U��['֡�Gv�� ¿R�tnFFƶ�#GB��\ؾ}���>}z��7�o4!f��`���|���f"�`���cϳg����x�Jm�5��^0��i��'��Ν�H�ì����Pac�7��Nƨm���]�Iſk������	�)�)�����d����>#��߹{g���I�r��6��_����7o.�H����v�Z��n2�Q9Iw�۷����Cee%lڴ	6o��������2���-�<��h*rv������d���k�@ �J�޹�)�ݻ;�޽���B�T�44���|�` �X�H���2����Y��4:��l0����ڿ�4��	2�R%��3�v���ŋ�O�|��)b��%@��[�24kڬwM�,�d�`�4p�$7Wg��k��>���[SSϞ>����d.�T���F�s'�P(�Z�p���C�V��B󟴘�
�NX�����T*U�>�;����'~����N�{q٬�LF2�I�e���Y�f�'�"M�Ģoz������,U�応�/r��ޠ8:J�sr�WP�a�*���N�>�"0))	�����d�������!��E���E� 4�@߉�`�b`�������l��Ũ�!22ҊJr5��HϾ</#����'�Ffޫ�ݥ����uJ.�I����VV�����iz��Ցr�<e�]�L��i@���
��ټyxz��GE�o���<x�y�.<Q�V�~�� {ezr��E|���F�V�&��z�����`	�!�͛S���Xy�8�{��\��#�v���z��d6�$���x�hJR��34pK�{�'���:)埄�����ز�.��)@��ǎ��ԛ7
)))N$����w�ܙB��l$�wF�@��@��.�(�ju¨c�EM�c^������B��,!a,�%w >>^��+t��s�-�ˑ�!��ҁIg��`��c0h�-Ŏ����NJ��/�In�V��s��M��
����I���%� r@�ύz���Zz7\0vl��&I�H@�F$ߐ�l��x����Z�ջ�TVV�mݺ�����Mt�Dܜ�fݐ��f�EȠ3H��+��^��d?��ju�޽���޳�@�T{�۷g�/�,���ր��4$�0>Ď��*/-#�I%i+�/��k�nm�hQ���`ggG�m�o�\���*MF�X�=V�d������M�8�J�8Х���he2��yl���|_��Ն�b�ϾĈ�^������qY�R��}�]�hA�+Ed���(o}|}�k�n���#*���?`�)S!;�*��ot��730��d�?:�o��GE�#7��P�ա�/i��ŋ��!����/���1tBΣǏ�}��|�l2?s��!g�%���Lf�i�P
_B6�CfWUU7C�*��㥷� �>$\�@eu�<H�@do/ٿf���G�b%-zc@�1:�1[�j��J�[�����b�QN�Q��

�'��>���8	fϞ	K�~�a�B����p�i��)��#�ސ88���]I_��h<I�������{,�%���t@@��B�6��E������-�d6���c��:�()ܼ��췺��/�ƍ����yϞOBY(|�$�j�#K�UU�cCBZ�_�p��˗/a֬$��z޷͜9�M''��4����j4EB;۹ s	V:�p�\��-~^~~�%Yb����R��̷���ܹu�� ����s&�2W����
.�^��͟�q��Ih����=*�*!~Tln�F�S17Msu�R�V�� ����`���g8n7m�S�M���bᣏ>�¶l�B�W������֛pFC�@(l�T4��O�Z�=~4 �ik+��=<<�?F@���Z�.5�>t��)dr���oȝ7`���`�(�����.Xb���q#���s�7��[�\�ƍ�����������k���|��BP*d���AQQ�	��~���5v�l}�|t�6�N���0iR"*,@��i�	�.��H2��ec�0(ʓX�̕H����ee%�6H[���@j��huݒ4�{u��o���k6�g7W�
a��~6(���b7-��wl�����o7��S7I�zI%^VV^���2���䤗�� ���� a�7�UT\tNlg?���`����cʔɰh��Z{�v��MHN^CM�c�����X`1�������H�A�X�`~�N3��~}H�������`Ϟؾ�8�>TWWp�W�@CZ��g��E�������U5�^��w�����v6�§D���S���
h��o�U۲e˨)�%K�����H����h��%�%�G��i����WVV�C0z�T^8p`T!Y.%`L�6��6m:��02?���oI��0 r�� 86|����BIIi6*B���[o{{{2�z�u%/��ς��c��ի$2�x?b�a2YYW���ܸq6nX�*��l|�"5U�.�D�C4�=8�02%FUÏx0�.�����nx֬Y������/ظq�ʮ]��X�#�]S#���R��B�|��v$�����qW�ZI����)..�C��Q-��F�ӧ�+z�kv��QH?zJ�J��<2�+�? r��`D�X68�:R$��K�"W羮�.đ�Fa����t�de�j���Ҝ�dR0bd<!��999�	��.�m۶�����`�h]4V�Q(\?B���l#��^Q��4f@מ��]��M�R!66RS7�3�^���()\VV��[;�[j0�!O@��op_z�Qp��9��q��X�m
�٘
M����:�7�m�&8v�(�J8q�{���lw�ڵ:���q�,):��b�y/1:J0�]xyz@UuU5�y�F�z��� #�3���v�ޝ���O��PH$�,"bX� B֎��1kV�9��.����d%0Yl�گi⧹7�h����='Y���Ԍ&���:v�H=1Ecܸؿ��v�ڗb1���dqU*%�J:1��+I�"�+�E7�e�?����{u��l��uf��,X�%��� �|�ͭ��6T�iE%�d)�<�PZZB}��G�B`���d� �T�Fs�\��B�X�!X*(,,����졢���3X��ܼu�.�#F����жS{8r��D���XD���_�n 0�$S%�/aE�*h�*2�e��l����{�m8��%yBs�	z;��:�z�]���4�X4x�M�َ��LX�|9�Ǐ$�f���4���v+��𫭭���M�NI5@��416����j4[v�qv��Bs�N6��.��t��5�s���H��VTb�j�&Qx���0f�H1�m?<f��}z!=u ���B=$�d��l��TR�o_�K������꧷n݆�c�)E�A�{�'�*U�$r>�XL��&L�`y�D�|��dd���*��͚�7i'�RRRfm�jm"O׫��yKV$��Y�@�32�i��Y�E���y�����S�����c�c�6j��1/��
 �p9R�B)�f�I�KV�0�(/%�(	|��V���x��h2�5�ڊ��J�2�^�~T��Gj3�s��r�NĞ.8�^������^�X����h4��E���uT���ԉ�1�Y��!����M@
� ��6�@`��m��OG'n@����l�f��^O�21���L����o���j��M���+W����qP�}/4��0,���[?�B�n��/f���*���j5?��`~~~�C餆,V�_�r%��	��-�Z|� An����
��Z���"��a� ��d9"@�L�1	j���Y���jukKֺG��ePF�)���'�`��α�ѣGW�c�5%r2�:�O�h���s+�J=��㢢�#�8�]nҤ)�5nu�0����1r�\�%'J�1F��54Z;Fw���9���U�˼\���QH3�\�=�O��o�y���t�^��>��B���)52�xL�����XPґx,y��yHG��L�L��B�"�E6R��Q)��tГ~ ��C�K��Rό�hu�t:��yM�p���1Vc�O�ׯ���	��4T�Kl҄D �v����+W/�3h<�l���K�
9�]�r�ܽ{��ظ��A�@@C_�(%'l������d�u �ʡ㸩�D�4�6d��\�F�����,I�FYY%漒��¢ym�t�\����\�V��� �"@����F:婁$#K��zd��<�N�nq��	��Jy?������	-��l6�����x�mG����2f�����@{��6b˾Z
3gςN:��5)��.<��:0-kP@d:#\+W��d��) �+���22n��pH�2��� ��19Y�B��Q#<�fx��	o�}Wg�{��¿˖/O�� �g̈́��ATt�K����wŃY��>�k4�Z��S��P��
���r�+�T�%{��a�!��{&�U�y@�O�cI����o�ii$u]$HGʙ3g~��Ǐ��5k����(��Z+՚�\TUt k�D⸌����L�C�1]\�~�#��0��\�)

>��,s<����5��%@ŏY�t�����e5Z��ơ�T�q�э���X��ɕJ���<<~�D��Or�*Ek�N�)( �+z���j��y�����y� ��f�h42��R|7����������v��ʮ]�����ɓ���B�ܹ3�iO~��9ސA�T���m���6!U�m�D��"�Ӱ�T�^R��
��z {LHdٱ����@����h�y!PRa����J��?a͚5��K��v��?�p�鐕�#��L&�ZPP@�f�o��#�L���HB�)n]~��0j����fW����={�LJ�`lF�
X��+�x���ѝ�I&c���>I�@����i�C��k��v�b�yEt�U/^��ҥ3���[+��<;�f�H��d����T����C���Q�� ��N�IO�� k�qq�f�+�d��/UX�T'���3�U���J�ċ/�xT��gM��嫨M$612@�ⷌ�{h���!;�YU�����hj<�"o�'£���Ra�n�������k���O��맜jkk '�	5?f��(N'�q���$���r��+����Ml͊��64�\�b�f��k���ku&�:'�ɓ'"H�����o���2�nބжm!�gJoa$R��>��NL=����YYYE�w���j���-�?��4}��'@��ѤO��QN�&��l�4j���HMݴu��ϩh#���Y= ��V'��ZjgϛK2h�Z����d�0g0_Ik浘�X�r0̈́y���������q��[BX��;"w�B���D�>Xk�c����7d�󏨳��`�*��x, �Фq����$k#\���aa�  sjjj�IO�����VRR��	ļ��w���U�
�1�o����[���7yr"U$�I�x= �5,Z0���rc۴m�����?��{�F���c�X�)])))�D�Y= ����	:w�N��;?]NrqS� �R7l w2���=}���G����O�˂<��!&���?d�H��!S�Ri(.� _��Ӓ�n�<�u�F-ᾩ�򖦐����:4!�Fӌ�����7�&c�s~��9<a��m�T���૯ެ�'V�[ڭ��@ǎ]@ �8���Z��f�+���^]#�s���P۬Yc���3��&oc����=}�E-`%MC�v��x��"ptt�~����4ꔏ�j�-M�D��V��LV��z�����!,�)^�烻��Y�`r�d�>�%�]$����s�����=|�cF�������Ub[!H�=�L�*����]>k�&e�	�[���z@���BՀ���k�\]��|�*'���|��Me>y̛4ʽ�o,����F~c1���vV�)"�u�!T/��?���ԮF͢��&�KA�<�����g)�4}��V���+|�2�4Q�4o�:��ae������z@��|�Z���>f2�Q.nv��A@��g<}�]�fq����,���VT��������s��Ud:q�0�3�����y�yCk׮3ܺ}����7~�2�t����E��F���<��-B��҃B    IEND�B`�PK
     eO�Z�Lz��L �L /   images/256658b1-ffe9-46c3-9f0b-70052a8fe00d.png�PNG

   IHDR  �  �   �X�   	pHYs  �  ��+  ��IDATx��|V������E� ����)aADp�m��[q��:�UQk[�u��l�(Sd�����7����wr�Ҿo�Jk�����<��9�9�ߵ��V1� � F4$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A1�!�'� ��=AA�pH�	� b�CbOA#{� ���A��Ğ � F8$�A�(�~������c��AMuՁ5�u�������p�.�Gɘ�i�
����1�ϫԨF���6*,�!��3i�TKbX�%66����I��gqBbO�Y����KK���yUʱ���VVV����o�Z�].W�R�Ԩ�j�]��z�q��o��
���w���|�>ӧ�c�b�S��s'�O-=^V_=%5���dqAbO�Y	x��j�jKx��g��::SO��O�X�ƹݞP��v����
���3��� �\ܙ�}b/���o:�Ri�)��.�jL~^��ܜ�W��
k3fLQBBB��/�_�3j*/�`V�رcI��a�=Ag����O������<�ő����&��i�A�\�%���T*s:���t0�n�_�:���~&�|I��{��UJ�w��O��'��>ߛi4����5����q��9��F��dj߽s����ɦ����322�ASH�	��444���?e�Y~�������Y�b6�j�d��g~��!Y�V)��3����V�x��q+�)�������ʹj~'����S*�\�5L��3~ߟ�:�ꍈH.�G�U^����a���Hy�ݿ\�eK̮�>ڸ*""�&6vzSF��b1� �'bX��+o%�~�=ל�89G�5��ydxX����
���tZ5c���|\��Vs�\�a��нZ�f*�{���p�|\�}ܣ��B�����~�F�t������+z��|U``��a�s�`���,<:��t:f�;YO_?;�ޥ����z���ʓ��^���7TTTl;vl#�a�=A�
����j���F��>|���*�d�ޠ5����
��ûf�w���v&)���px=n�G�V�Mƶ� S�A����u��ڮT*�*���+S��*�����v+�����(��q�ݧ�z��S�Z-[RGk����q�4�B����RxX���::�Y__��j�&�tv%lްyv~N���[w�;s���H�*~⇆Ğ �az�{o�7f�g.lom�B����tڠ@�Ya6<y��Qd���˺;Zw�J�tH~_o�(s��`(�<qr�ĉ�'L�Rb4Z�CBܡ��.����yH���������Һ�{Lojj�T]Y1�QU�a���f\�xi�̩��c���T*+���;:���{�����ܴ)z�5�������=A�����̏?Z���d��E>��r+#�BY��,��m����b���hsi���QW�=)q��Y�g6dL��:+,�ʒ�]�գ<�9����{����e�ڸ]���b��'+$6=�X�ľ��q�2��Ա,)>�e9����͊���ݶg�NӾ}�o̟Ny���=A?(����7�xg�����٭�MxҤIL�R���f�ZYuu%�.�[�P��v{��ys?���+����T7{�}����ڵ��s�����|16n���z����6,ٻo��ͧ��5*, c�d�5�^�j���75�Ym��������;�|C����8����=A?�������'�O����7Q�����pQ��9������YG{����u�����Ą싖.�~��%��9��CGW�v.�k^{��%[�ܺ����Ç�����Ξ��,;�kl�W��5��v?`\�nk��,� �����_���B�jժsy��7775_8*(؜�<V���,*�!�]����sK�E�V���[�r����͌uGL�h!qL�炟w��o)߿��M_~���?_ñc��&O͔n��uҞ={ّ�9���3U��>QW��=�W��'�����_��������B���*���Xrr��d���ɸ��:�.{���3>����0c��SW6�4:�|+��\�ȯ�jhl�%�+cΜyA��%�>���U���$*��w����_���X��G�W �'�ƚ5k��{�}�dgg����	ܣW���2���lLac���n��Y�|酯L�2�Ȭ��+"##��, ..�^S�gMi��-_m���]��<k�ܠ�.\�fa奬��-�d2���;vgMMͺ��D#��0$��#dpe8������i�)kkk�*�Jr8���dx���U�0NYYY��v�o�v��Z�6��2�Neaaa����UWW{��z;<o������g����?�:�%&.�x�m߸��ŗ^�eg��3B��@���)�lo��Z[R�v�&d��}�3��CbO#�I����an�#�鵛^y�-cWg���t��>I`2�bc��~��#%%�388HYVV�����^o@]mmLO_�J�R��jGL\tSld\�}��
E�ܹs�������[�j�9�o�|���R�ә&N��ƏKg>���46���}'�͙������{�M�l���%�_޶뺕�Von8YV|��i��5{�t�X.++)P�NH�8�߃G��85}��J�{}� �C���⚕U�?�Sg���[o�ڛ=���2�n������n��`2i�
��U�����9Ǐ��u�\m6�e~�/,,4\k0�L�ؘXM�QL�R�~��wwvU�U7��v:t�=���?U��NZ��3����L�G�fS�G�N4�'�YscS��l�t�+޿���=������n�.<���mDUuŭ3��2���b�֭cN�M}��=��1��w?��?�=A�����UA'N�*�OElڰv��~q�
�j��	�+J*�w���fSPP�&**�EEEI(�s8̨3K6����*6*8į��bw�ޙn�e�,66V2����L��0�����G��pF�w8�W��~�a��1cJ�@�گ;xpm�[o���V���iu2Ʊ	&���.T�{{��*����,[��}�4��$M���嗟>��㍊��㿈��0:���ٸ�Ө7��v������r8 #{�8K�{��k�E>�x��ڪ�s��	.�=���.%���]{�0��1���X�7�V�*��YYI	���c������.��Rv��!�xn.��4Ҽy粔�6~�xQ_͏���e�--��+�qBB?���0U@@P��q�+���s�n�fSNN~�'�!��>��`�ω��ԢINzZ�02�?�kjj*_~���y���o��F6R���v��~��<��T*�OOWUTְ��zI��E�:|��"�k#�� $�q����~��?$�[���ްX���Z�[T�\�L�����{�2��ʢ##Yr�6.5����`{s����o�����d�'N`[�����v͒�$���˂��Xqa+//g%�eb���.*��N�r��o���QoB�z�ԩS�UX�&�ޱ��hNN(w�c�v��s��cǲ��:���ҟ��U�_�e$���jӨ�Ĥ�UՕ�q��)&�^ji�e�N�R���;v,惘��Waq�!�'������/�������*�F��fWO���;�ط��r�a�ys��1cX���{�]�o�C~��z�q�م_�R�$���Ē����l�l޼y,/�۶}++**b�M�X[g�Z���(�w��»��|b�w�R�Z��Aդ��fL�v�sY�)���ň�Amm�����a�ٳ{�_�=��7���ǯ٧O=��d��W�+jOq�oc)i�����GGG��fq�!�'��.�?>��	k�o����8O��K~�u�ٜY3��Ø�]ΔK���������m�^����-m->�^'�vE|\���v���|���6s�46g�L�P_�8�*++E4����=�����
o�ǅ^�T3�Z�=�����o�XXhX+1��&9�F�b"G����?�|=a����,\X�~�`�=n�lz��WH�S����RIY%Cӝ���(��=��~?H`b�BbOg��v�yYG�V*�����j�o{�ܹȷ���J�ƍKe�kdk>Y���~�������=s�f.��QQQ���Ϙ��"
�,Y*���Y~~>۴y���b�j�z���J�ZB؞��l|���Zč�ѣø��Xk{+���#Υ���9�v�)v����*lu��=���̞=���\�ƯsO|b��꺴��pstd(k;��j�k:������,.�G$Z!�8����0k��s�=v�	��e*�JU\lkmme-[��l�����Zzٴ���ŗ]�v���>�0{���)��{���o�.--�ӫ��-))�����F�Դt65s�X]�P�a�?c����M�4a���7R�IĨT:��鄇h6���ec{v�.��r�w9]����j�X1.j,4|����2wڬY�3gN��߽{���>���N53�lT��7r�M�=!'��'�&�;�w��z��Ğ �1\�������;���j����� �ȣ�\HH���رcǘ�a^t"����3��cOJ���7_�s)Nq��ں�膆&��ϙ�.<����6m�Ċ�����
uO�<e�k��V�އ�e����4����"8$P�!��u�؋/�����7�1���
57zYaa>	f���Δ���+V�vⷿ}�貗���W�u��;Ƅ�Eu��������l�ږ<����$#�3�=Ac��zo�u��Å{6z*���#|?c��m��_\\�5k�&��_����$����w�yd�̙b��-[�dnX�neUeU�b�h�"x��o�9zL�CU~l�hӡC��|��5K�/)����������{{{�>��z٤I����/��zN���v�v;�N�c*�f:u�����ʷ�w�2�ӳL�TJ���y�[ZSS�bn�UP(�8S��|1Lپ}���z�j�Z}��fӠ��f�1.�lΜ9B�Q����❕u��5ulʆW^�)Y豤��?x���SS
�Mr�ϟ����?~���c,�av�=!-�-���h���������=\�c��
��m;�馛؉'��ÇŪu:��V�G�7D�\�3v���O�����Ԧ��r���f�nZ���ȑ����s�.:��4<�@bOÔ��zgjC]��\�#���$x��c�;D���yX&ğ{�黹pT�|����/+*���޶���W��O���cݺu~.�L�VKN�������c*m�F~�mŊm�7o����g��o�=&Y̗/_�.��B1�h��-*�}>&���,+W���M������c�q��{�+�o7�Lq�]�a��"rKg?��2Fg {��p��{ﯮ�@)<n��፟<yR�V�T��s�eG��<v[LtL�O�����o���w�!����兾���ɽ���G���Ν+��#G�����FnT���|��ϥ���T����i�9]r�%-۶��ێ�_O���t:%��&
�0��������` �x�����$����iC�w,=��#G���ޫf�����uw	�][U3�߿J�Z�g {�f����9���p��Wh�������eӦMc�ׯ�����"w�j�*?�����x��<��3b,.��7_��¢��'.�=Z�~�駶-_���7^���-['lٺe:7.��{�w_TT4*<r�KT��*�m۶լ�dU�A��ō��X�|Ǯ���³G�Y��c���>V[]gLJJ�΍�����m�L^���֭;8��l6���k#�_CcsC㤎������A|OH�	b��}�������\(c�NC�]��Qq_VV&������gG�������舆��jkk-**8���\?R\tYww��� ���%�޺��s������c��W��S���p�xK�,����Ƿl�ꊏ�WA�!����cS�LFHVV�8G|�������ɳ�����09�`�=;v�?p��ew�*�J�/�^��j�LV���Ğ8���0S��9m˹h��Å�C  �b����0�m�Ν�cǎ5��������O�>^iai��fOs��*��ŋ����?p�.#=����z}'�g���x\>�l�: 4�ie[{�߅�w|�#���t�J��#'��PB�1�Q�`�O=) �?���3��[�ܷ��^y}Cʘ�����:n���Xz��3�M�X1.=�@QA�T�ק������}S\\�:�F�{�^�����q;�?Ey^�=<hL���c��������{��{�<������{Ϭ�ݥ*�2c�3�!%����ݱ}{�/�{�B�}]6�(�����x��w9�>�F�w�⊺�1�UU3������c: ��w�ƍ�n'��A��q�
LP*3��-iM��M�]���Ą����3��kn�_3OhHh�Z�v[lv���`N���d��1�8���0�ĉ����).�K��=����Eg �(�Êu�G�fǏ��;;�~�O_-���{pISc�e���:�-r�))�"Wo�Z�'MJ��Wu���fx�>
�d���
��\�zs�sO=~���o�N���{z�C��=���۷��	C$� �;>>�%�+��A��%�{�fn�$�v�/,/-.8|���_}��7˖]Pο��~\�L�~��߄���`������E3�8���0���(���X�թ�]Cxe��#���zܛg�������i�gW�>Κ5k"gg�����pq���z��c}YYY�7�r�'vc���r}S]�.�J0$�so�+elr��C{��p�܅?/=Yv�Z����߃���xD]*�Q�9�x�6s�`[]����G{a��&��Ǆ�sZ`��qú����e?"P�����ڜN������G�o@��ɳ'�$�1����O�|8D�ox���C8�Z�\o޷���A�!9����+��>�?���"ae:c��0�9s���7�pC�O>)�-..kio��jDc�$&&���'��\�}������r~j��`<��f�<yDpNH`v@zz�0Np�G���xm���|+�lK��ܸᢟ<%s���[�z��/df��ƒ��ǂ�9|>�W��p��%�/ay�L��@bOÄ���<0�{�>�_(�!r�1�!|�+B�\�}-�-�-_�k��C��0u�C[�0���-����3�pv�}w��%ڵ��744�Y,��N+��@A����1u����>o�.G�^�W�\)0��B��&��'O����҄QR[[+�򵶶���:�ýz���>�1���Qp�W��J***F����
>�⦦�]m���S��~$;������Y��@ms���=A���}}}�c�W�G�����v��9//�ŵa�ҥK����޻wop����J)��!���*OUu�%*1�G�B�r��@�Fm��"���/))�Z�VUT�I���o^P\T�4( Ȁ�;l8/DFǋ9�)i�����:���OOO�/B�1QX������5����|���4eҘ�)5�7���3fL/���i��5p����)
%��n1{�{AbOÄ���p.�q��!x��Dq�}9��Ű;#}¾�/����q���EFYi��|-��gφ����=��D@o��!Uaa�h�=d谗�����i��+���oY���cbb$D	P7 oy}L��5g����"�)w�9�(�F�9��ʏ�t�%^��˖���)Z�z�%���Wqv\ww�v�qP3�靌���͛�/㢷��05O��!����1!a`�#�N�Q0�8���0 pO=�T�#.�hӯ ����l��%d����z}��Y���oݺU��K�]`��֦e��!���.+;Y}�]w펛���7~�1����z} ��x:V�[�hQ��/��?���R*�����bw���"�PYyR��s�9�&���E���������o�j��܅6�n��O�x�;׭���ͱ�1F��I�ȩ���e˖��_�F8j�ѥP+<>���}�לi�*�U���K� �'$�1<���0.�F9�P�/��#�����xJ��˖���wO�o߾����y���a�!4_UU՜��s٥ˎ=���b_�:�r�,���ӹ1 �υ����q��w�������)��֑N�~hы�{���[�����`0 B���5��$S�ө�vI�-�#e���ʕ+�{��k��w�Z������H��ϟ?�Hv����^s�Q� �9y����^r�'�7$�1())Qp�8�?��b����s<G���Z�[<\C�333ݧ�����t�F��!�΅�SZZV�dђ]C!�7N�R[[�������,�h��]�;���s@��I�&	1/,,a{�i�0H��������{@�P��40���Ï������SO�����[��8ݞd�f�@������z2��۱ԫ��`�V�����p� j-�y=>{�@bOÀ�� %�̯������Ã��56mas�]~��f>}T��r�-�N���� c�{]]]uMuŇ}������=1��rM��i�]9z�C�l�5k�J�qC�-X�@̫G��oi���
Q=>o�<Q�___/<z�h��l�:����	��أ��;�s`��S(�c��.��r�G��	�����>K":�R��5SkT�Q��@�8���0�j���p���)�W��	�G�^��"4υ��_�]�������wL�O��1��˽oGk���}���-7�6�������h16�u�PU�1�BF�P=��fΜ)�
�����v�m67Wj=��%�?}�tq�0 ��E�!?g.Z�eF���|JJJwl\���S���s2"z���#)�RtN�D<����h��W��p��&�t9�?�� {�pAWq�3Ωf^��!t�",��Gę�;!)���i@Q����O�//-��X�{��t�ݻw;F'�>RTV$﫼����_��ף�c�y��x��n?B�s������j��;\��;233������0�L4�A� !~,�3�	�/V�������F���/�.t�q�Y~�Q�N�3"�!�ɵ�GU���e���T�.����)��?�l�$<{��ސ��0��=�:5�Ȟ�>D��x������3>>�����b���ZMIQ�L�R��v����p��jjl����o�ݺm��w�c���s� Ӹ�*�*��F8�>y����t	��t�>�Ç��vuvy�w����}~N!�@!`tD$�(+g5�UL�|=�R���=N���_]�3f4��o���s�垽0z�o6���ų���Wb��-�|�_A�{�@bO� .�7<Z����G�!�t��[#C�:�}�m�?��T�\.����T���c��1Q{�?~���;y�r��MF} ���0M� |R�O��Ԣ{�ѣG-III�<�̳��SP�� /���X �urQ_B\�h�s��qGLtTim�ߵ��;�q�4�N�ǫ�hD�Ke��E���W-\8r+��5Wp+Oc���E�O�`�?
�=A�e���P�`)���C�\��Փ��:�)�9���x' B �@��\��]x���S��¸�����1�Iŀ���=����x#����ͣ�.??�u�ĉ�_�x�/��xç��uuuE�5JVh��΂C��޾n�ѪXrrS*%OCC]۝w��<t��g���{$I٩R��
I��z=����2��V�X���ܸQ�e�}\.���+�`q �'�aDW�v���"3�N���iY\��z���u�|l[Gg�@�xʠxs1v�]��33�n�Ey�����}��3���@>��<�q��q����G������h��O?���B���@][GۨQ!��_UU����8D
0U��6����暺�+W����t�U�w3�B���d�+�O�gl���G~�H��n�.1��}oo__r��ZFg {����XE^U����" D�vgg��`4vpA�3�ө�1O[^�{{{��j����ڱ���6O\�f��|�p��E��C\�����ɽ�QUc�(� S�zo���Oy��C���с����Q�r8��;���zV��]p�,=-�:tȲt��iii���=�t��?*  @���XJ��SkU����#�P-77W�_P���5M�P�S�B�:��@bO� �	{�X:��	qǆ�����6fS�zEl?++K���/��l6����(**懺M.�����3.���( &�PT�9� �"W�����c�]yy����;.}��	n}C����z���� g4�Ae�^�U��Jtw���u�U��^ii���1���q�8N�N_�w��`�EYYYf_�T&eA��Į�����u0�0{ap��������H�	b�E������'�է{�{x�r���/!!��{�B<O�81�TK�,>���S������Kԋ">n��ǅ���~	�����v��Gm��	yz��Q̱wG�G՛�7�}��]����{zzB�㙵�"�#ִ�r�ǏwY,}�,���kPZP�t��ʁ|~?��\������曓>�����T��at8\������7��z��Mz��Ğ �^.�X��'�Ň�A�e����y�X���t�mwfp����g�V��WUV�_t����~œ�?y>7&b��-.�^��#GDQr��L�:�r"��қr��_v�e�����@�����$�?�(�C�������M{�ۼz�	Xt���ܓ5�w ��q�5�NNN�l��5k֌�ꫭ���o�)X��_	��6̌���O�4)�a��1�8���0�{�{T̋p��fV.�?��1�>00o����M�u����F�ё��T9�۝NG�-��R��˯]���o����N�u��C��=m�q

r��H��ʟ^YϷ�s}��ק<��C�
I�Ӫ��iw��Vװ�s��+���mٲ����s�����|�g���߿~����9�f��}8G��['L���F ����7]��а�_k#���jc����v��~;j'�����"����^~o�rc���{@bOÀ��t?�C�$5ڣ������B=X=/�Z���GtvvMP�����7�8p@�������1��^}KP`И���G��`�:�u��="a}�;vL4��b�z�u�o�{`��y"�p����h��� ����|?7V�E�EM,�0o޼o����Ծ���сB�pN��Z,�������_�p.�3���#��Q�C�Q�)�� �;��)>a����fAqA���o�� �#$�1<�r��6�v�Zh�;���������G���D��߻w�8�Z����^/����h4s�lW_���~�beyy�L�J�			��@�X�f͚u����itj��	6�|a$�;G֬Y�իW;R2RjO?�>�`̎ۖi�Z�"ŀi�2X������ؔ4����6o��������/���/8��=��c�^m2�Y���J.����4q�s��I/�����Ɔ4�+p]N;7j���#���
g�a"������w�����<��R���8D}��
�=A�G���_oV�U}�[���{���:��A�9����z
�p��%!�?�7�b�?o�;w���p��B��u��O���K�«/))��Ǎ��ϡ���l�o�p9���<0���At ^iVVV��ٳw�7��}]]]���Ӄ��|L	
nL���τ	
��{֋}^^^Tuu͵��"���w������������ q���b@�^��Z�jkk����kA�0���0atLL�J��ȋeN���v@^�V���\ҕ�N�F�f�:�<>>^BX��O?U!" /��g�f۶mS� !}tAA�h�s������տ}���̙c����C�z(��r�z����xH�۷O,��*�M�6Y����-�sA�������?�0/�X�Ұ�PMgg���\���=�E�^z�o+����^^X[[�i6����?�R�������%�Y��:�,��BE�9#���=AbB��$��U΅�X�.7��#���FOXd������5-��r�\���'�~k׮=�!���c\��ܕ/2:B��Q���;�`����Դ���.����ac��9;;{�Ag0@���z,��<�M7���ν��믿���q��z�{��	���k�p:X�F���u__�%2"j�UW]U��_���͔���***Z�����h�������3�����QB�-���\>��g���.�FL���=A"�.�J�ƅT�s;8�|h<�*������F�1����y���!������q!�G�9y�O����X� �����k��{>K�?��6~�n��cG��q��'@�?*��`�ϻ��}�`�[���7^~��W�x�}�V�^��ٙ��]��7~^>��^{�]������Y�!�6lJk;�:���(���A�����9�������ǆH�������NEGG���6 �Ğ �	Q�����{��V�o�ix\�z���@����;��`_�5�a|.�C�va@8���<yr����G#l˖-cd-�-�믿:��s��	����?���!�s�
��:t�SVVv�wO>����.///��n8�?5"R уa����p�y��v[�����f*+�����sZ[O�r1��V�r�j1���=]��R�`}�}b?���6]YDDp%�+2������0A��t?�䓅�v.�f��!AY �EEG7pﷵ��8�fwDc*���z{���
�����Qe�p>B�xD�������~�M����#=]\����uu��h5Z-�G�v��>/7
�B��\R����~k~~��W߸����r.�*�"�|}�7�$��~$��mn>2����B�FgF�{�N�s��G��p��%&&��0��Z
��a �G��;M��.F�{�FD��Wp����,/V����6�R�ʊD��C �^t����T�C���=��!��Ə/t��r�<�$W�ᬖ՟�~q���X�fHlsrr���/�)ƅq�q��������������v��c�����Þ��ӗo�rӃ&s�	�z+]]]}
������z033����ٳGUY^<�0i\̕0�p�`(���=�OL��{ ����Lkk;"m�>�?ۋ�{�F�DE�p���B�� @�e��أYG'+U�4.�:�=r���Q�./�q��$��00^Ûĸ������������9g�7�2�322��K�^s�5J�Rc!{� A���F^ّs�����x�.�����_Q~m�q����Sk����8W�V|��>���ȍ�>v��T��N���:�i��`4Gj�zq��kjŔ:�?�z	�O��F�10�ĊJ~i|�~o[A|OH�	bߧ�jQ�?�q9�"�>������8�zwO�V�T�PԆ<�r�B!/�����IMM�dII	B��ŋW756u����=��cor�
s�\{�O�9�w�
�R�p3Z�����}����.,(8z���t��k���&߽��?���/4�L�� 	.���Ғ���)���+y|cgeee�윜��{��_x�6�-�[[F��l䏡�����nJ��qo��q���,�����ǟkE����Z��q�PkU��8�e�=!�'�aD�:֮P)��w��v�!���!��r��Z�����8��Nrr2�I�����vq,���b=��}�����ƥ�����tY��W�~>{��ٺe�e\��X	=��!������1�~���������?���Ʀ��8OD$`��,����f�8s��}��p����e̋/�|eQq�r��6&$8ج����:+��4X,Ex����""E������!&
�$�X"��LLL��TQaq& �'�a�;��c>�E��� �d����y�X��$���A �G�a|x����r�^#|��o�������[���ުU��SSS�&�%�]n��g���f�d
P��M�&�n��P��4Ԯ޻o�f>�\�u�������55�W��5��1"�w9:��w���G���'����&++K���_/۹s�]��3zzz�����G@��O7��op��S"�"�O����߮����x�C��,~�X�W�V72�8���0"66��c�6���-q+������д-�A�~�r';���}�	B�8b��(��^�/==]��_R~��w�=���M�*��ޓ����g)$�����!е�����YTP��G��رc���s/���K�޸i��5ZM4��\,�����x�ҥ�>��'�س�����G�k�{nh%���)q����y�9��Eő֡h���d���,V!���x��`\7�Ԣ�!�����AA!>��u)�NFg {�^���P���!x�"ޓ�!|x�p�'�`��{��F���v�m���`͑#���^r����?���w�����y�%�{�5��p;ЁH�ر��r97���/ݼ�溕+W������,_�f����8_�!�\��⯭�m����˭��x�l�j���XXXxm[[[bgg���0^pO �E�xËG'<��!{�yuu�@�@��A�"�czc�R��&݈Xޗ��!�'���l2�wj�|r��� �P �o2�~�o����@4 �V��?�'��������4wGGgyyY�SO=�.##C|YNNI��o��?&�����5�1]��/7'�yނ���r�-�|��?�bk�����-[�n��F��Q؇���
�{�z?���o�Y�d���ttt���9����#�@n������;�v.�3p�����(����>��%0���1X�������O���A|OH�	bx�lT5��n��yyy]{�����x*��Eoz��0��x��# ��1�i���{�����
&N�X�\t]U݌�V�|=�?��g��IM�4z�����'pT𺫯�z�_?��?��ѿ�񕟬[��	~|rll���?�"������M��|��7~��?��ݻw�jnn���X�Ψ75; y꣜FA�$�L��	���b<�l|U\���O��9�hYYes@�!�loL��������=�.N9t/��!�w�P/�OJJ`��ڵ�������9�J���ap������q�E|��u�u����zl���`��K=\�]ee�o���}>_��Tp2�������Grs�{���/����G���_����?�' 0 	��"��Da����98N������s�}������l�ԩ��Y6�C���;�c���[�<ܫGټ�������=L���@)����bj~�"����W*a(���f�F\7U��u�����d0���/��.F�{�fp�ݪ���\ܱ��p��CD���z�#7�f,�h�2T$�R^w�mq���M���FC��]�
,V�=&"*���Է��ֽN�s�������8�`�C�u���n��H������u~e`���?����1  0�{��
p�4���a����7�|���
ϖie(��ꫯfq#kߔ��i���\y�B<J�n7��6;0�tZ��ao5:���'�P�%�X��V��w��gKKOz�x_J#��0�߇Ğ ��u�����r�b��`�\=r���C8 ��c�6�m���ȅ{�aa�5���I磌�b��-�w�V^p�y����̙S'�+1)%1!Q��s?38(��KMc���e����:t����Γs��He����?���훥��M�s���=�p�>�����{͕W?�«/Hg�����\Syy����͡|��{��"�*Γ�;��
�Y��>�.�#�"�=9e0
�V��6��I��JU(�G$�����;}�a���@bOÌ���ns@@��a�s�^���!
ȿ#��GU�躆��w��e�#�� ,�q�޺������:v��|��_��~Lxx�()�Ȅ���1�^=ml��X�pN�?�/���ܲ3���o^���}1edd��cq~mmm���l{{{��;n���/��ⱳM�:::¸A�ɽz��H��Z�,����2 �����z�퐯��&�=����K6p����,ǔ��;&^��!���3��7 �'�a��,���j��J��A<ރ�8O�T���b.J."Z���N;��$!�V��M�8�A�/����8n�����--i����8�d�If6�E�?���?~�Dgsc���ѫ����H�ǚ�ڥ�A�11�QJx��q����!RTT�mw8�?��o~�r�c%/��;��1��{���}<��«�Go�����E���|��
��Z������d6�˨�3b/G p��\�߇�������1�qC*�Q�>�oBbO��۹�p���������@�[��"=�!6��!B� ��*��9b�>C<_XXhh=u*�{����k5ڡ
r.������%���>]��>v�Xد{⮆������.@j��r��������/y��W���2.��l�_SGG����UqMY�z�G/�C�{�@=��[ʹz<�:c,x�96����3���tC�X,�����H�F��7 �'�aFpp�#$$����O�!,����1���q!Z��""���������9���Od�w�F�<��ʠ��+>��*��d1�3g�X�~�ڵ�ή�c��/�f/>+ί��B{߽^�Ŧͷ�7�L�8~��w-Z$�瓛��mjj:����Gz㪫�j���<s^^qBmmmf}}�Rn�+O��W��������{�CkQFa�aI[T�L��3�܁r��ܞ��	�g�z*�fW��4z����߄Ğ �\��z�������"��bE4 �}��v����tZ�yn=s�B�)�v��k34,L��|�i���R���[�VKKs��K.^�����/>x�`����s�=�0����u���b5���lgQqa�Y�>��}<&s�Y�j[MM�n��o67����@�e _�fJ�J\KY��>U����e�s�>H\ٳ�+�a��Qy�B���y!�~�Z����{�fp��k5Z��C���I�D=l	x�(�Bu�B����C��c��9x�r�544�G�{��ttt0����Z3/�͝;Wtq+,*lY����o���{��펟?��G�9|xQ���IIIRRb�X���-[X}C�������o���s/�:��p�%���u֩S-\[�Y��":���;���x���r�6�}�S�Yxx���ܳ���`��? G������r3��#��ew� �ϷNn�uR��w!�'��dw�Uv�vu��½��!�T�C �yx���0�[]x�UUU� ������k���>D���>lT�-�PA_RR������ㅹ�������u6�Ƙ?4~t�z�ر��ŋ�����A�=p�@�Π����~��{�-	�����Ӛ��2;;;U�� �-�E�IFN��@�q�po`|̫׉��={|����x-"-J���z	��>�3��7!�'�aFWW����%�{�Jx�)))C��x�F7(�۹s�7)��!2z̭�s��!�#*�=t���G_�޾>1}���KD��*))�^z�G��ܾ��/�����uQDDhTb|���������������h(���+ޛ5#s�Zi�G�ʕϞ��nx�D<B��˞���dn�s����_|>��E}ܣ��7Z�F�9�/���N�ch!y<D�}uk��2���Ŀ	�=A3���M�M��\��x�:�9���Ѝ��- <w�tx�XUǔ���\:��P����b�^vv�( s{=����"��9
1W���q?��,sG��OKK�_�H��g�D
l\L�r�;=��V)#�u�Y����@#����9����\�˞��؍<�^L�\bX~��&V���6�x�o*`���0`Lx��*���{��A�����0���6�{�)\$��Bo!v;
���� �F��"a-W'L�����Ŭg�cd_�5��uuup1qr�11�m`����1,<"��{R����(w��fBȨ@aL�r�4}z��T��
0�����*q̘͗]|�>�T�4���q�֮];���ijKK�B�GO)�(O����v�ϓk��Zů���%?3��C�p]���p��pq��e�>s
�
!�����u�#�$�1�@�?��O�v�-���G��.w���=�vx�X�^^�Nn�aF.�fTݣo�̙��ޱV��10 <^�0��G�V�����>�1�%K����L�V*Ĝ~x�|\�F�>��.{�׏?�s�ر}���5��6�W�///_����h	�C�i��j���N}�
xH��mq�	��N?�t�E|
�S���MKK;��{�^HEEE��S/���{��! �N��x?����A��9<T�cqL��x=����1a�D77(�C� ���ԩS���3Ez���$;z�������p�·�硇HcǎȐruuu7�洵�	U,��b���!~�{�,�9�����"�EopM兊N�����D�c�$w��
�8���0�����0���Vͷ�J�B�9��l�EV�w�H�.���s�=��A\f͚%��|��!0�o�����׳޾^�V�ED �&
�0�^?턍
���C��1R�%�\�+\��-��||�I�t��'l$��f���s;;;'�K	Cx�
|���,�2C��=z�v�0�LF��
ꞇ��|ށ�u���Y�V�ɫ�)*���h4�������w�Ğ �\�%�9�-��ur�T���k��=x��@Vi`n=��x�j.Z�0^"��h��ֈ�$%�3����rs��{���I" �A��ȱ\WMMM��hػt��y��4��F0�����{{����q���sys����j�0מ?�<���۩�=�u��$.�A�L9hd�>^=V�s{��`b��fw��>*������;�W�P�����)�{F�{�F���)���2&J������� �����^+C�a ���U�V���Qb
B����S��@����葫�>��#z���C����޾�}�/~oŊ��͛��c(��wtow���&���^^�Nε˞����)���%��J�bA�!⾠�3%�X������!{n b #��>�&�	�������`#���=A�w��ի�r���r��w̉G���!(��������8v�7}�t���!L��=��>B��T�C��G]� �(���ʲ��ח�U���������C5��؏~�&v�t'���+��p�E�{���t*�p�>w�o��s��FBP@ 3Mre����J�"//�˔
>�R���1����N`XF�{�|��WIO?��%\��onn%�B 7^�[����0<�sT�˅y۶m�� l�رbl4�c��L�֋><~��zx�?;;ۗ�����y�z���?�<��'?�I{�c!''ǰaÆ%�mmA�i B����ˋ� ��eч���1�5�hh�;���G�P�Q^���y��{�j��x��x����"��>���̎;�7n���9.����(P`�?���� � Wi#�����~#G��W\!D
b�c�:�xD�����Ǵ2n(��98m6{�V�]{��{�SB\~�~T�q�kNCC�J6��!���@L��`��4�@��~�թ�"((�����7a�9�C���y�L)�-(8h7{�rG|/H�	�$++K��_����_^UUe@!���>�.j��[!����y��� zx� ���c_���ahx���Qe� 7��{t:�W�-_��mw�]�u��q�cK�~����r(
�O���AxO_�NΩC�e�?�}y
����f!�*5*�]n�c�F�<w�F�N����qkDE�yH�	�E��d�M�����!ҡ�%���A���c9[�b����X�.77Wx�W^y%[�t���C�e��#������T�ѣG���J�F�_����͝;�����f?V��4�B"��>�F���l�#{��llP�}C���准�m����%ϯ���3=���8T�����j4�ɔ��U��{���"n�ꫯ" �r�<�}:���nx�͋��ށ5�������v�[�h�"!�X��{K]]����;EO}|��{�6�sm��ޒ��;É�����B)�R�(�P�9�sh�i{J����BKiKPv I d�Ď۱;�۲���}=�nE�������\�T�ҫW���u������߿�c֬Yk
G������������+��A���$���x�L��G"'kZ�R�.>�F��w���j�$��*~�=��圽���6�m3sj~�����>GA�� ��a���'�WYVV&	�����C�jI��8 ���� q�-����q��G�^#r����f�����۝���҃=�ˉ��׭['F:***L����ȳϧ���9��<���e�dL�xN�Ώi�yш��ɕ���o�Ez8'4|ހ��!O>%f�s4��+J�9���O��>'@��GI�����<����s�������AOJJ���͕Ev�^{���O*6m�$~��/�w��b�ҥ� �7o�<�u0 @:t��P0���~�Є	��	2�2i���W�D��C�0�4!�h�v��?��w2�����FM�8#3]�����>y�x�=�������GB6�u[fff�PP���^A�s�����nҹ瞛�\�˃�}�A)rs�E���/1��# �>��@ ȯ����g�u�l�{��d��w�!+���"o������x��+V4
�80�رc�[ZZL�#q��z#Z���>�t\P'�ɍⵘ�W���r�2�#�!�hH�1���M&{ 9��7��i��Ǝ�#>(�WP���s�α'N�8/''ǁ�;Z����e(�9�9n�8@( r�¼�_]���a���׾-�/[.��y�^"�؎;���3^��v��U�ˉ��A�Z8ݔ.Īy,x����HX���U����xD_Ph	�Wυy1�)�l�%�`��fSMNN���t>%(�WP���/8���o�� �� �A�B�Pɛ0~����HB ���@ЮG��s(Г��k5\�ׇ6>B�h�z��%��>���'"!%����3�(Z���kBK�7K��>{�L�ɡz�٥R���n�pP�;f�8s�O����0�~��F�###�t:v���7)!�O��>466Κ?�۷ow ���8T҃@�����5kD��Z1w�\MU�<FTԣh�����ܥ�΀�u�^!H���E�����0І���뮽捯\����@NU�O=��$"�b�����6��� ���O���y�
z>7x�hjyZ@袧��W��N<_O����)�9Ft��§E�

������ם
��b��;wJo��^�v�$z�� ��h�"����?�	y[I[��x��|��P�!QTX$󺻻DzV�_(�2��3�h򠐑����Y"���\d����N!kܰ�(���F����9���̣lq��,fa0�Z�Δ�0tH��A����i<I"�it�����1�~�ʕR@*x��B(��F(�z���Ç!��իWK��cx�rn4"'�AL}�dP��E��s�ٹ�d��Y�f��P����������e��P�>n��#��yv��N��5#!5-E������Ee?�,���2��5�a$���!�ް��v���)B����i�[o������q��Y�+��F��y�u�G��d�-['EU�aI�0 @�x<g��m��曒(�g("`�6��fs���&�3���eU+���V���D��n�녂��7�yrVW{׌��>}8����D�N�[ 
��"<M�8$��^=��Q"h�1�pBa#����.�C�yR��䑣�Gt�o !�����|��c�hOFj�{ӧO�

�"�+(�F<��Cc[;:/��O�C��;��1C�\/����#��@�=nx��_�Ey����^Bhdd6YD*�=�� ��E:=N_k{KkgggD(H�!do��[��ޞ���.c��~g-���� �H+.k���h^���a|��s�C����b�s��p,�?�p:�2s2��§E�

��iY(lkhh�!L��,Ё(P�b.�q�7
�@���ݻWz�����Ϲ�xݗ<���8_zzz���!�W�����ߛ={��ǁ]�:���z�^+:��5c�#O.���D�>M�����1R1�#�Oh�k�?HƗ?1&���t�����RTTT%>e(�WP8������_y���۷�@{�Ƀ8Ǝ+�Cj�Q��U� ��o�!��._�\����dp�8�]�i*m�&�q��i3}衇�	��z�&�áQ���ҫ�z��A�ɹz^g&z����(��i\����[�����[��H��>t̀�f9@�Tk�§E�

�999���rO��Ly�
���5��b���<q��G�=�� =�������5&"����;j���~��m��=��BAC]]���_=2���?��L� j�E�Y�D��O���(���
��]�U��Ď�A�ܯ���k�K���as���)}Q�ԡ�^A�4aW\v��ǏO_�l����xӾ>�p�B)���y����ϖ��?�Y�Q���Q�a�<ue���7
?]^Y� �ğ��7�p�������ZBkn�h{��Y��n�{&e ,~CT/�7̉����@��1�1 F�ܱ������1��v���(����N�r���0���m]���&1��/}�K� �
E���eH@ށ$�#o�#D���f�M��A4D(>�Q�*��v�2m޼uv4� d�
��	�T�~��- ���0���"3;[���	��&���ȫ��}y{zO��zb:q��F��#;~�ӵ�9�W�L��^A�4���9�λﾹ����zTȃ�'M�$�����ر�� ��`T-���AJ�=��D�秣қI(.�*ϯ7�T8�cp�ĉ���ʳ����M��	˵�Ѩ6��s���o�ox��j����,�&���@89e���yv=�Jz�VkS�˽���X	)|&Pd�����������ݻ�ʼ�<ǘ1c�����D:����+d�8;;W��#���{L�CX}0Ddd0qն$�L����&"-�.����#G�L�,&R7#���i���[�~��-?���`�%z�^�}0�5R�Ez�|=0.���С}���9+��F((|FPd����������w.�}NII����I����~�x�c���_,���ң�\{�g1�p�����y�1�'�W:����;�ED�K��򈲠@�ə�������(�L�އj
'����\|>��'��k���rr�������*|fPd���c˖-����雑F�~���2G�ryy�rn=����G�>u0�.�H������dV���DhXJ���.����)8x𠧽�c1����z�!��x��s�G��dX_;� Eyd��yk�s���z�~}x���zͣ�>�W��o�L�D�g��A����g�m6��?�ޱc�r�9�w<g~ڴ��x��g�۶m2O/IF��'tn	���f��Yk�B[ˠ�@0`
��bE�������.#�	�FD�C�XC<���<���[i~M��E|�/��'�1�a;Q�^WaqXjU��g	E�

���}���~���f�ܹs�,�!z����.��@���_��� ��G�}x�<O�=Ȝ{�?^��fD*���&��@yy�������<)x���Ë�&��>ޫ?�7�SA��{�EVN���x`!h�sz �߸���h�

�!�+(|Fؽ{�����ǎ�>}�t���L�3g�+V��-t��ݴi�,ă! �t��*���IORhÞ��+vŧ��,�v;�p8�
	466�7�h<���Ϝ<q�Gق��b��Z�c p��FD����D[x��q��O3�x�}���
_�3�"{�� ��Ֆ���̜9{Vq�h<z\�1�f������ϗ��ꫫŻ�+��<	�d4I�7�̧tq>����2�0�#�v:��� �a�������m&��°�� ]����f�{����ǯK�����*���0C7D8"I�`4�P$,����	h�Q�:d���0�owNN��W����^A�3��O>9�H�ksf�N{뭷t xy�行�|1=/��pH��h%r0�5���Ɯ`,��"Gz?	�!&t6� A�����e-W
�6p��4K ����'�������&������;6�,c"W�) ��������ϒ��~���C���§�g�y&}��7͘6s�K/�"�C^m���/�)w���ٳG@I�HH��.I
]�]D�����
�vù^9v5����`��FT ��;=N�� K(H��Օ45�X��y-}}=D��D�6�����b��zM��Eq�=��9ߎ�=��].a6����C��6�(DF�`P�Q,�(�`����l6k娒q{�8[��E�

�"�����K�Z[ZϪ����b(�8o֬Yr�| '�!܎���f�B:(̳YmZ5=><|x�ɞ=�X��D�����^k(0:�	�ƍ�����q�.��:������Σmٻ�
ſ��Z��F��3��!��v�p$�����{ �Ͻ���C6�AI+�(�WP�� ����~f�o�^U�� �%K��!7��E��{�79��x �m�$� y�n-'O��ܱ^�'��*�qC�v�FJ��&��Cح���Bo�d��~�ߞ��%�.�H� �����y[ D��vڴ�S�mٻ�1ZZ_�V�gНT8�sr����l���


�BA�4@���§�7�xc��O?���L���Ўo~ڴiRB:l2�W��`T~CD�h0&Tِ�7H�$Β���}��s��p4��`�Z�:�����4���`�����[�ږ�A�Xw)cF��c��|��XK�%�{�I�&��e� �E�.�p":�5ԡϦ�鎦���j���i�"{��%�}��?�a�c���N"��Dব1�b��Ų����u�DUU�(..�Ă�<�D���-���z�\p��� -̼߽{w�Tp��j�����V1�A�n߷{�}}}�H�`��5�֒���K��	X� ��5��!��Bg4�(������v0L&����jU��p���^A��|䬗^z�?�����!3do���j9e�ƍ2?�7n��UEa.� z�7A��	�^>HG���h��*�=�_��Wŭ��'�����N����ܜFo?!F(����ݷ����3O�(nXG��s��V��������������Cn��)v	q�6� �����x\Ə��tN�+(�?�����u�)>��{�(fgdd�[��u����!���6���7��=t�S��<���нޠ���'�� ��m`8��Eb� �t��b��xL���.M�P�������q}}���V0�@�-�Z��	��2��I���߸1ٳ�!�5<&W����F[�3����o�s���i�"{���������E7nZE��9t��r�h��g�� z�AH�����{�Խ��a���w $���#g���tzA�PD�����N�4�ǣ���g�����?�x����MF�D�P�.ޢ�u3�,�5��G�:XS�%�� Hσ�Q���@��±����=��O(�sDS9}�N��p��^A��MMM��^{m�ڵ�l�YKɳ3N�0A΢ǅ���B�ض];vLND�����{/���,���=�!�٣�n��g�6�˰��%��AT >9OBb)ج�L]{[{��hll4������0��Y5d�����>��#���
{�ח(|Ě�r!"(h��>��dּxn�������q�]�Ǎ	��n� ++KU�+�V(�WP��@yy�sժU_�����d2��m��,����w�֭[E��:Y����@
�������A҆��SM<'�_�J���	p��+����=����	'��qLNN�a��=N1BA�p�G7n�8@�uԨQ:�P�>�汞3f̐��A��q�"ʶ�QYY)�Y��1 o&�@П���z ����O&�:'���dl

�����@���ǅ��kn5�ӌ�iYq����}�$A T2FA�q<(=px�L  yx�����ω����ٜ7��| ����28��),,$�1������֭۶~�{�>����tD�r?��"#=C�%<x�U�<,�v!����%��0�ൃ�x��D(�]v�0��F����^2� ��Z(?.�1���RSS�
��E�

�l�Pg��.��X}�O��K�m���D^~���#?��w"?~��Ǐ���{N�Cc�$q.�C�����Oa�d�V�����9A2���ڌ��8\�\���n�S��zoX�0�����|gOG�/*�T?@�;���E��>���Q"b�#��XO�=�)tL�":Y��h�3�Mرc��V㬳Β��o�D���M��J�K������x�j��i�"{��@���Ń��j��ڬ�����{�|�߾}��Ӄ����⎊|T�c�]]]�$} �y]L��ų�J�g�{���1��@��!�H���Xǃ��v��<T�׈��4iRpa�{�}���JiM��A�${J\�����h�i�o{z{�A�װ�_~���W^~U�޳[D�M�/*��ė��%i���={9�0fТ.Z;_}fv�v�w

����@��ꫯ������H42��t�EI�[x�6R���+��R�x�����͛�Ԭ�6F5�y� j�'B�1��ᡳz[�.;�˕ݲG�}��كXXl!c&���̴G�WD�P��e:Ru$F�ѣGeX�n�	�.�����_�����Dh���5(#^u�U�k�յ��׿��܋'�|R���O�.��iU��'1�Ӿ� '�J	�(|Pd���	 r0}�۷]RQQ��` TL�`�:u�,��I��C�m\��#���w�5��� �K�i��q���8?h�m�1˷&�鰷��G�4�]J����}�IOMO����buO<���斖E�^FBXKDV@�H�ȼ|����Hb��(+m��<��>�~饗d Q�.���80�9gp�x>=z��Q�\��^A�c �����:kϞݷ����Y�9&x�йG�ҷ���X��*Ty��[�l�3f�ذa�|�a�@���y�r�,��ЋlǋK�&
�D��7�����x`d ����\�g	�.�)��G�ș�7n�l߲}�i.�kC�s��a�"(H� ]����k�� t��aTa`��z�)Ҡ
��r���~<tP~�-[d�������o5�k�W��yA����G@���W�������8'���8��T�u�
�߳w���G� x�<��5o�S������N!�iH����MRY-F�i=�B����1���mq� ��r$��o�?Lf������	TS��U}��<�1CnSST���{����~ЄIv�����g�#��AZK+���0�@�F9w�s�HT*�� H�Ȕ��7��?@ ��`@tt�	��&�>g�4�P��DS��������6���$>'(�WPHB]]���G�C^���yO�x<f���у�Ql��:w�\����J�ҥKe��ڵk%���~x��іĄ�xa{� ��8 ���z%q�9�+���<D\p<Ρ�U�%<z.���cDJ�"����ό&�h��� ��"�(h���\��uXc<�>�t���djE�_��@� �V�555��GF�*�[TT�%>'(�WP�\W^y��U�F�9�.�����KR�^Zyy����������Q���E���\�#�� I3Q |�|1��^9�>ފ�~L�9d.�c�T;��!!���.ԃA�E]��V�{�ba����ڣ�i-r��uXs��#�k�'O�"= 댽�2e�ܳ`\���뜦a�|� �.p��ر�[TT�'777 >'(�WPژ��{�����]ta��葧-))�Ev���C��y �˂�����x�7� "����:�P�9�A� ��A+ �}�G[�3��\��'�y{�=��'�����=V�M���:�ȞH8}�����>x���hD8΄1��x�2!+�s0���O.��������� {�׿��/�w��@�'�o�n��!c�͈�P����^a�^��w�=�w���H$:�ݼb�
�䎪z�c�?./�h���

�@�K�,��*k֬o��v�R�%T��j:ق�cUy�9�,����q����L��Hdb��j�勃��!��03>���K�imnM'0���m߾{|{{�|��ԯ�k���"!9�EU8t�<�����z6����9)@� �#�OF�����r9�̙�*/^���w�Y���H((|^Pd�0�nݺQo�������&�BY}� ���o^4.���m������G(�x `xy,��cpCN!|��W���kgA#���a~z���蹭���wx��B2��Ȧ߅p��i�۰a��'~�BDE6�d	d������D�-��ɳ�9_�G�Oϰ�mxF�4�Pi���o~��}Ng�֬�^2�w�u�PP�<��^aDc�ڵY����q0���4����!t�q�F�w�#���W$Q@<e���Rv����A���A*��>���s�$��{��q�>���7�>Jd��3���
�@b���KD@�=�ga鉨�:�w���#���ȑ#�---�#ak	č��Q�@6�8�V�Tw���H��s��4 �~�����!:��i�&o��W�P#l�((�W� O�����J�o�"�Ԝ�� ��jm�Au��ɭ\�R���K�$�
|L���=-�X��k!xm:�#n�VK�qΞ���d.�c�X�n�{�?l�DB_�s��=0(`���ۏ<����F�=1����Z��A�\	�k��ȱ�±S֚�����>�B�!��F��c}��A����p�A���w�y��Ç3
��Z�q���#d�ۆ��DH=��P�O�{\p�UX$}�Q9Ҷ�<�X$J>�z����l4	��*<.������~""o�7h�RpN�	#��8	�b�h�sѢ��͚5}ǪUߛ����I�nĴ6xz������kD\��������S�Ayy������D3�}#���Dd���z����,����RT���e���[�p�p8�7x�Q�
��8�j#��+�H<��#��y���7	���Cv����&��A��ʡu�P=��8-V(�C�{� n�<�<Q���w/�xq�0/9�Ϲ�DH�nt��k�����;��M��&�1�}�R���=j �#��Ym6gK����kjj2��:���pJF��� R�r�x40�9�����sQ ��9��d��1�ɸ#//�W8��^a��O�S���Է"���`�P�5o�<yA߹s��9���Gn^!���=g�Id0H��r������0O��ki!w��>ѣ���0���h���E�|ii�")��j��}Zn��91�����" �њZ�@g��é���h��乨\3��ɂ���z��t@��M�9}n���=<�Z	2���
�-\��[((��Pd�0� �뮻�⦦�/џ��R޻w�l�CXy{\��ţcly��̙3e ����3�b{{ \��㼈
�.�0����er;�ϳ'ʕ�DZ�/~��0���������Ԟ�^�a`��`R@� ���"����Gٯ[�ζ��si
е��=��Y�`��q-�h��������L� W�'��K�^�3f�f�[�W8#��^a� �9��s�܊���`3� uh�C�}��PLC�0{�l�b=7<h�rq�G�>���P?��0*�A� x�L4<܆��8�ϯ���&�c��\�7����l�͛�Q^���f�ǘ� �E͘����/..�y�zMb`ǎEd��Mkj�����}@>�)HF�N�Ox�X�`((2�� d��C�L�ɡ}����������BA��"{���`��7n��\�`됗E�<�S�s��zx� 	T���>�@�9��'J��y(���ʖ��)�#dY\9΅�ǫ�eX�ivL>,��ae�zmw��۔	����~��]����~�ȇg��9<���o ���f�8v�q<��Da�۱0������̹��.D{X�=x>�����0�l�SSS�ӿ%��p�B�� ���?��s��|qss�sT׃ȋ�9r�{ҤI���6'��@Ax8b,8�y y��Y9d�-Z <�g�Z��e%=��s�����0r\��>*o !��GD@M\pA0������=1L��L�>�����9���zbt�]������b������^e���{"��ρ�1���dy\����.4�=iD�Vˑ���BA��"{�����g��?v5���t�0�}�'N��ѭfժU�x��/>���@��!�Cˋ>��!�;u���/�-�?�a��#	�Z��Fx7��%�B9x�f����=�>o��	�ߣK Q�O����T�,t2,BD�^z�d>?���I�|:������۶m�iii�F��[&��,t��hE������ᝢ��D/=�S�5�|ra��Zmf����B�ꅂ�E�
��W�v=��_Cg�׮G���ɓe����>�ǽaŊ��o���q<.�.G*�D���r8E��bI�}�b��]"=%U��hJ�����e^�{��@a�8	����$�P�����&���<D��U��M�����?������1�y� �K��J�{�.QP�'220��i���������61�y��_���119��7T"��ޘ�W`4�d�C+��P8$�����T��!���ǡPP�8jB=����}�ܹsG�:��Є"{�a�\�ryvW�� � �lmݺ����~����3���p/µ�����e���Q�����$�9�g�_zIV�]zը@�$Ώ>�cx��p}��v���WT��M��#ŀ��
|��!�������>q��SȄ���1��;|�nHE$��RS�-��7�׷g�ܹ�<Z�4���#�Y�ׄ2�o0&�Ӣ�O�ɟ�0�=g��+�q~�ö��zTᇅ��E�
��w����C�Y��եÀ\��\�{��9����x񂣿�ݓ�t!7��Q����$��8(..��:G��jzhwc%5 �5��L�A�����#j�6�uvv^��d��Dx�{��^(�'l���g̘�Ͽ��S�>���k8=UkD�  �63<#Ozj�����APC8����x6�v#�,�Gt���>&K��5��n��@j���?��Q����x��+����777Wy�
g<�+[����꫗�]Do�C����������<�߭Y��Yh����Ё��G����Mk� 0���_]�1�?�Q��9z��<{��A2�v�Wz�1�3g����u[�(�L/^����&�|��^����]�hQb&.}~��������O�q��@�R�-.�˟���lN��n���0�t.��+3�7��CTk��9�5+rQ{�R�(n����"L�8�G�r>���h���YO�PP8á�^a��駟.����voo�h�x�@�(�>��s�7�xS'y�5k^��.�鸈��j�޾^���.�z�8ހnI 蹇��mnт��P �@o>�d/� ������+�m�׋�3Ӹ �G��=qv��uyǎ{�~N�k433����%c#�#<����xx���p��ub�����ݵ���Ʌt�}�^�*_������<����`��u���g^O�+bQz�pNNz�PPPd�0,�6�o����F����pG�=H��^�3f�sW\q���~&����Q���e[���D>w�\���5y��H�'�xB#�8h$nJ�A��i󔻈֦���s_��k���ߗ��.$�p2�� ��H���0�-����뮻���~&/�gϞɌ[Ȝ.�ŉbb�Νٽ�=e�F�W`<����8E��&� ��{���ϣ�Ye/)��6��! E�
�555Y�����>Eёg��+�Y�s?�裏�n��ɭ?��/�K�w!<u\�!������4i W)\����߲��H�W�Cr�l0�d@���A�F��w_qŗ��9�_��Nz���&��@ 0\���^RR���ºq����H�\�Ć���������:�OX��a5~U�/���J�w ����X&{���Z'
����p���	"##��<��G�wWH��Ac~~�eeeJWaH@��°Dee��P(8�.��dnAț7�z�U_{��.kX�~�����Et1���4.������������A��W��}���Q��v��ᱨ8OWw��;1�˗-[ր��}�����qN�t�8/���322�%'L �O �!i�a�}|_��K�8��L���0b�d��C������w�#g�)Yޖ%p���`�Oj�y�4<&z��c?i�C��[&L[>\���+;TWW[n�m�e>�`��@~PE�|t׮�o~��C���?���<�Ѹ�O�6-Q���ϗ䏰:f؟ι�Bi\ֲ�A�(�����B�$�<a�j��<O#+%U���x���<s��qb��������a������9���¹`|�\��D�[===�*g�¼o�q��4�n�$f�B�'� �b6Ya{.��6<��c/�������n
�OOO��r�:����"{�a����Gg.�h�)WUU�:�;==�D���O���t[].�ԼG_=���ox{a�?�0�DΤn$2�*z�<i��p(X���B�a�1c�v:���7/Z��F��s;����b��n"$�G#���!U����y��d�	�b5��P�F��;ڏ��� b�;+	X{��������}�� .�c�c~�N�5��zv�;vX�1*O(�WVصk�����%t�ϣ��9[��#��������Ǽy�꺺�<{���Dm��=zT���'fw�y2�{��!Y���1��9���|����a�6�xcD���Ν��+۶ms����1�%,I�V��xxpz!����YZZ����
ٛ����xx��p8�z�.Q1�@�-���s&�>�o�����a��N��_{�X����D�Gv V��	�&}����ә[�B�
C	��������⿈��#ú E�\�\x�[��~��e9�%��®��M�B���P���8���H��˹�@� �����p%��DN�dff�7n���{�������Bz����%B˜�����N������_�>777D�ޏ�x�u�,v�L5Ģ�.�d�v����~4������r�`ر���-#��)ޏ�Ev�&�ēy-�8&z����rrr���:�����"{�a����"�qmm��@ƸH�'����}�s��m�qZN��"GF֢�|;y�2$��<�7���;njj��B� c�Ճ�9d��ZǏek��П�����zQC���p
����#ud�~�?�+��K��Ii)//�|�O������K��mw��Ϗ� �`�x�/������q!��|Z++b��w0�x$����Y��G����{B�Hb0M��V��SY-v�T=ztњI�&���"{�a��>���h�J��;&�^����۷���n��c�����<L�����GqH�:��#_���+/� �Ǳ��8.�����Rp'%�vٲ���gD�o�=���Y )&h���~���\���Y�W\qſ��B^�b�`_O_,�q&D`�]bxy��,�{;�*<���O^-ooH�=��W���!�1�~���*|�G�VCt�=;���Z����"{�a���Gkk�z�ƅ��������e8|���K~��eD�T�[�.!�)\L�{����4@��omj�ab��A
�!G��d���'�܇ƌ������������غu�l�,Y<��@6��� ��c}�����D�a-�!k�\��z�` ð���L�e�w�͖q��� ���wh&���m2iy\��^=������Rsq��
辻��`�)ST_a�A��°Accc��A+��A�ĉ����9r�Ͼp��ϛ��.�6H�2Q��A������p�)[�� �����E[x:����O�V���;��4d����&�2p���Y^�dOx��>���~/�>9Ϗ6�=� 6��+b�0~Y�ڔ��\�R��<F�
<ϳ1�\��������h����O��á� #ڛ(���˯�J+(	(�W6ػko�@�ot,޾~��Ţ�X��������?��g�?7�\��U�(�7�PT�&���.�sDg{�cH �=H�o�+��:=n���.s��P�h��sΜs�qc#�������;�x����mfE�P,��F��"I@��	
χB�62H>Q�.ә�X�q�����8�������t���x���F�A/��B�F@�K��7��2���A���Dl8����f�1�b���eGC{���m�����
_a(B��°AOw�2OJjZ���4-�������{��ܲe�SO�~�y�g��:}4,�����:.�ܶ�V.x�ȣ��A����H���~�+���x8��l��7/���F���_Wf��g���) 4y�Q:߉iӦ�?���wDS�.�N���w��?�70��a\��@]���O'�ͦ��/:�xRő؛`@
����(Dbm�7"6��9��
\�ǅ�:}L�-2m�������
5�VaHB��° ��푇��v��9�����m���ZXX����7��!9� 1k}�~��� 3�;;�E0�}���sT루���³��t�Y���M~~��e+��>����:��j`$�߅Ea�x�?6k֬�%h�,\�8mg�j{��x�[�y.���YZZ:�G�~������Ydyx� O���fx���=k�LB�`#I����<<�V�l4��~nQU�
C������q�M�|��B���?''G��=���ǈ|P�V ��t�A8#���2H!�.�'H�.#s��yg����S��CA�F�|��0�`�3	��TO�'��;::,��}9�t���=U����>_[��C~h˾}����[J�n����a_A��A�oբ:�S<v �6�.h��<�V렽�����@�u�qO{�����&��0D��^aX�����.�I \�"������F��� vx� ��� �Ç'�� �- ���v���钄�gу0p>2
�3�s�̞=;A����楋��X-V�?�O(�aZH�QK�e ?T��477{{{�6�-!̃4��y� ���z{����!]���o�y1���d��A�}}=�#�}��5��ܥ ϞC�h��M�7=����uQ��-�F�~��z�PP�Pd�0,�Jl6���J��h�'B��E���-��������Z�2��牐�1 n�N��AL� wL��={�,����11"����ª��nݺ����,"{��ᔡg�����N&�{��O���n��6�ɒ�A� ��=�x�A�+���:��׿�������Ѕ5�;4�� X&nV%�J|.ZD��卹=�+��X�Q��X5jTA�PP�Pd�0,���ta6q8��r$.��^��j}� �!���~NN�4��:�����Y��|^"����^+�C��_����w���gʔ�W��ﴬZ�*�7���R�ɜ� ����2�td(���h).���~���w(���=΁����d/ d��7��GCCK	�mi4���1�p��oliѪ�9Z��b���	B�\�g0�N��z�@��1�v{���|b���P�"{�!�w��_��Bg��2�]wO'��11c�I�0&N,�>�|����gAqOA�����9a̺G���E�$i���������tãFm��׿��֯_�����6ł���{����y���DA}~x`��N��mw��5���4������o�9��H�M����Oa`�џ���E>�`6���{��b�":�Sf�'�q+"֊�f� �F<r���[[VV�����O��� E�
�(��s�.�^�1c�l�+�8$.��� !����h}K\]��eO{`�_�����/_.I�p��&��t�� ����oڴ����2��������ɳ7p� �����#GL�!rss?V����Q	d�Y<��\������E������[�������$z(�`d��AZ����i��X�����VE-�oL�<p�s��'�U��g�cZ�PP�Pd�0@\�7#��Xi![\��������F�-[��|;��R/�)ρ0�<�>x�\���?&��A�{�����[T�c@
������=��ɓ&W�7.�_^��߸ 7q��=N-ݒ(�w�Ϗ555�ô���߽{�yǎ�9DPf�>?~�4XP���Z�[�������r1$#�(���_C�����@r����oX� ����}9EQ��" ���6�6I� L�6��7�!E�
��b����m�\|��;̢G�~����
z�1o��r�8ρ�A������<=��A��y���x���퐤��8j�Z�f�V&9��f9xh����$B��(�{�r ���L������G?���(q����\c�~3R�p�}X���;�-/?Աd����׋����
Ӟ=��o+v:�:4,����&��v�S[� ���<�H"�r��m|�ۉ���w��ʆ|����"{�� y�z�u'�bR��s��&M�9mH���+� RS=���E�;�؁�a  � D��=�d<�x�b���'ı�u2r�9^z_����:�x�#�߬�F�~��������k�����@��O��cɞ����6JӃ24�߀N"������s�;;��]<�U<&�$6nܘ��־�$�
{�;[&���m�:���t��v��q�{�ТA��d5=:�����1c�&�^((U(�W�E"1��*|G�G�|��-V�$Cxy<Z��h���^��5# }�x/޷m�6q�M7���<�_�J�v�g-��߿pᒍ+V�8%�Ku19��Pl�<3�����s�|���蘏%����2
���V����;%�y!"�="�@zz�>2v����={&�i�6�}(�ľuww�ܜ�IӁ�OII����s�$����w^����)Sz���0�"{�aV���=�=Bܗ^z�ػ{��z��}OWbh,��}ܒ/�}��b�̙3�ڵk��_,&N�(s�K�,"�:_�^��O�����N�g����|��W|%���_�� ��3x�-���5��;�s�=z����|7���K��2�ш.��@F-�5PUU%SH��ǹ�-�_UVV6$��6l�`��o�\J{�	k�5����A�6w^[*��'�.�cOk/���ȡ|�?����P�n�陙{����E�
��X$ƅX�߱D_5<�ˮ�B9\N����xSS2$��|�FFF��j��R@���/�8(N�$V��<��S��w���}����!�7W��|�Ё��- Cɨ!@��	��}����z�>"�f�1���򗿌߶m��۽ހ�:u���q�w�qbC��~W�����˿T1TI������7���������Gs��a7I�`/�G�b͹z�g	 8������:T�WT/�	�+y�ڞ�Z�����i��s:����<��L�Mdk�0Dh��́�녗^YY)�F�2*�}���d.��W_}Uz�ȋ���UW]�я~TY:a\��~�@�{���k#��x�;U��"����UZ-�߁�:F����s/h��O��li��tӅߢ�K��Aqq�$@��{��W����c:�;J^�'*�� b���'?YH���6V
�:a��,��S��>FD���.�K��J` �g���޷٬}������6��0L��^aȃ.�:�٠����H,,�VSbj�Ao������[TU���(�9x��,Q�Cq������cnEE�0[�◿��x���C=$~��'!������;=hc/�D}��6o^i6���.�q1��@8붭d�X���O�*,���C�5�_�/�~�_��������7���Am�U�qϟ?_z�����X��DtC������r�رgi0���~��G�(����c�1�9|��d�ҰҌ�݅$�k��"BW�?>�H�q���;v��p�0l��^a����̌�ѣ��d��Z$�y���'f͚%6o�,*�u���<=H^#dp�ՃL��@��?a�x��g�}V\��bժ�Z\�\�p_ߠ!�{���_�F�����B�g�}��7��2���Nt\4=#�Xnn�)R�0"���"��<�[��@����wF����Z�Zc���]7�p�ko�{SE�ڵL�B��f� ���)���PP��O��GC��&F�~�����kCs��z�� �%�r�v��U�S�z�aE�
�Q���%yƋ�ሬN�����/��KJ�w��E��ߖ�q�CN�����<AM�QQZZJD�F�>@�ҹ(��Θ>K�:,�o���;0p��<����S!�\��k�e4S����&���3sJJJt�=��d�@0 R<)2�Od���8B�=���{���g�y�n:&��kʔ)�|;w��0L�H������Y3�v��W�!��/��+�|�O=�yc�`4q��߁�>c�./|��"	A#D��|?a��qn�����

�"{�� =�z/��>�%�@���	�{�c����i3�	o$�jo��A�𔳲2d΁s!OD-���^|E�r��bӦM�Ç+κ��K+SSӉ�Eh��]eU���q`ùA8�sG����S���E�&����&ϴ'#=�n֬Y���-[��]|�%�FU�tF�8ߜ9s���}�6�}A�h�i�G��*���֬ys��ؽ{����s.�^=���O o.j�
c�x�L�<����>�<�8�Dt8��s�v�;���

C���<���M�Ĳ9�ٺ��va2�7�/�2��j�裏���뢘�sx^#�Y��I:m
�"�w���+��:d����m�v�Βz�w�q���ן���ה��>����*��u{JJJ:�����@gGg�/��mm햮���z��;����1cc��g/=� ��!{�E_��-.,,� z�A< 0�m q!t�����}����~�k��FE���M^�<�mf3��� brN���=�3b�XHG���" ��w�^H��:ݮ���f��0̠�^aȃ� s�-��.��=Z��oEVf�,�{���Env�$l��dIj�<��z��9� )���x�qI ���z��ݍ#B�t:�mW^ye�_>4�Dc��D"����C:�n�ׯ�ڋ/����գ�L��A�&�q���eZ~�����{�}�8p�2>\c#-C��{�񝠖��s2@�����˖���!��o���>��(�S��{���,�Q!@��K�^�hiD��z�-/��J�A݉W�w�gf�=묳���°�"{�!�h6o�8����d	��1�!Y.�����F�cZ����@a@9���aQ]]+C��s/۷\.���/��ؽ{���ν^o����w�������i�n�m���q!�����W9�x����~�y����&��f�0��a�Z���[[/��B��}�m�v���"�RH�3`޼y�C��¸��G0 `�lݺ5x�%���o\����q��x��]55��BA�Y�D�|=�!�oֶO�c����iam�Z�����tD�m<�!c�b��ҝ*��0��^a������<}��EyK�,�a�,�;�D �mTA���EmZ6�#����`H#��C?�BF����+lV�سgy�ex����o��C������i۶m�:}�?�_]]>����կu���.0��!�gB/��:��#�H�H���/������fw̥�a �!� ��{����(<$c F���r�_��_��oC��]�������9��b`����Է����k��KT�#���?�<��?��7p{\[Ǝ-:*�!�+Y���[�KF,�'��Ē����C�¨���􋜬�q�D�������&r��D8�Uk�([<��a�>Q��( "��A  [�񄴽{�B�NG�@֚��Xo�ז����1YY9���?����;wμ�� �ߵk���뿙F?A��<m��z1!���?��K/�|#��tz΀χ���: 08@p 3�l�qR~�"B�����8CV�֭֊��h1	#���~;�^�A�Sʑ�M����&��>�ɶ�����Ω K�!�3R������ԇ���	���$�mn:V3�����cƌ]�͙��"��ĉ�.��(/� 	�a�k��c�M!MT�'�?��Ri�h��!u�uT�#'��=T�PYB��,�  ��Q䠝��
䂢<y�Q"��߿��������/�477����31 ��mٲ%����˯�^}9}��j5d�3eg ��E�50 �]�=[ZZ"۶m���/?~������dDyZ[[����Z�{�����<����8���އ��0>�����8[�N�ٖw,%���PP�Pd�0$��6y�)taw�������uww^���5.�p�q:�v��������%��A�i��ĉ�(��;�� ��yh�[,&IzA__�$T�����c�}k�Q�uu���>��@2 o�#�N�=2g���9��g�������윀�<�|������42"d~�����I�^"*�6D`H���9Ry�E���~����o���+���A�ӄ=�aF<0�ɜ�ay4-?��	�{�[� ��S�(O�b5XTT�$�)�+������f����5��{R\�ğyD춘�����ȼAj�c���o	�X����$�B>hȳL.<u����ɕ�������AVNKK���b:y.ǁG�ss�<����������7N�<�|ӦMW�]�L�,�*x=�w�� ����xF
��Et�>��wp�ƍ�s��}���{S7
˶o�6�8��ZtF����:&|��sZ�}Th0�`�����R���Tϋvfddn�:u�PP�Pd�pƣ��elwg��F�
��h"g]o������H�1�i�Y��Har�$���Nz�ȉ{��RZOo��h!ވ���%2�&�<O��$�}����H;U������Y��4ѽW�ґ*��1{�0�Ճ�A̘�N��|����z���h$ZH����| �d�^�=<�D��T��2<bt�A��]�����O<�fb�c��ծG}�bz��<Ĝ���d/�x����/Ya����� C,b6��KK'U|tb���p�"{�3���YN�� %�m���2�
sxhG��dO<���pӽEd�d�E��V����x�W�Л�&I� d�(����"�ǃ�iiG�{�2��T�xR��Ճ�qz����-�����UjR����Y:�����ލ�;�$_�y�����e '�.S�}r�-��=z^~����!�喛���A��P�-W�Z5gp�?��Հ5�n
<<��1��Cl�.�CąC���{p\ M��c/阾�TϚ���BAaC�����;�B>�b2�bD�XLz� W�G^x�̭�\��zT\�
��ȃD�Z,6"��Eb2<O��dtBg�B�w�����,�~���|�ŗW���|���C^����+�I��.z��$�cr�<r��5U��$��f�7�#<�� }�0�"3�<"x��@�xm���Q"�n"�mii���{���7��Ad/�֬�m��o<�b����W������X+�'<������aH�:{��O��Ţ�HKAQayYY�*�S�Pd�pF���3��(sX-&�REj�k�Ǐ�I�wh�#L�כe�E\~�e2w��Ҧy���:�����Ga�Y�ۃ'�^v"�O������o]�xeݹg�x���_��ko���dB˻Y9�3�g�����QF�;9˸r�G4�3����B>_�رc12x|���ʱc�>��q���r�1��o��1\������u��� B��<�ֈ�ϳ@��l��Ғ��U�x����o 狷�E�SUa�*�W�Pd�pFm�U�[Z:;�B}����������Č)SEw�8��$�k��A���q��K�,���D�vI�~�����Z��@X�R�Vze>����XR[_�7�2]����c�),|���k�]�Je0�����ƹA� ~A�t���$w�g��H0.��-|2$M�!��M�<9@�n߾�X0�6���9g�<�@��ٳC��z�N�
�#�<2��b���Q�`�/ג=w�O����J��8x.--C� ��j5p���ǚ��J{�7!��~��4t�aE�
g4rsK:|��_zn�ٻvo3ۉ\}D�Շ��8�b�¹�P�;&'�բ(O�������d�m���0v��J�<x�N�C R��:<m<7zt���O������}G�T��D�����Z�$p���(�h@���A> �� ��6MM�  L����Hb�*�����B����o�}Ϟ=؝�������:������+V��y�1q��+�&�����.�K^' ����NN6�<R)��~Ќ�D�u����:u��Q�Pd�pfc`����Y���}ͺp�\����4��y����6���+&L(��M� EƁdNH�	i�]�Ñ�0�uR/��w]��ܬLǳ���N"�hOO�A��ܬG�<�E m$��B/�B����X2��ֶi@D"��w��h�ڲ�<f���( A��q���.gE_o������l\龥g-�����_�|yd(��Oq���Q���g�ڹ��5}�_����9&{`��x\Ҁ�Ϧ�{�jy,��=D��j�(-�]���F �+�����Ni车�D�]����>�{��"FČa0�hL�E=?�P�wv˰m��M��Ou�ǅ�o@�,j��N�������B
�ȃ3Py��$@��<aH��Y��}�Q��r劷
�F�{{{ct�X8��A���ys�wF��yD>z��=zt���ޅ���UWl��?�`���'F
P�������)���cM9\�^=�}��y�G�A�S�+�Y�7 n4x�
׺\�;����"{�3D����7�C�����<� �и���x�ͷE(����lq�X�x��e�}A^�8V� �{�|�"RS��e����>a6DsS��O�O�= C� ���\9�.�a9P�@& ��ɓ�����o4�t��w=v�M7��B���j��{�.��~(�o���m�h2�y�����0sD
�����N2�.���P�~ъu�,�0�su��W�c�`�q�=֚[�p�.��k~��q���=[

# ���8�b]��V߭�H�{�>�\x���'��TMl�k]=�"#=S��o߾�܉�S$�VUUˋ?��A�	�X[F�M�A��|B��yDMM01/sxT�L�P|�J�+�c�'����nw�ߙ2y��w�s�s_��|7�|���������w��;0��x"�q�����X���4�+F(ȸ*&�~:�d�5pꓥn?�8q��AG4NKt9pk#�U��Cz��`NN�q��0B��^�CGkp��7p�ѠˈFB�H4,rs���~� y��r ��E����q�P������˖-����EE�A�M��]D���A��%���G46�":z]L�C�D���"'7K�*�5=��Ύ0�|����ZZ[*�L���o�|�o���Oʫ#����d�O��~d����#Ԍ��4�h:\VVV;���{�%Gye�����43
����"�d�1,ج�ٵ���^��l�&J(�%��(�f49�ι�����р�6�%v��wu�twuUOC����{�?2��w�3���l��P��ԼB�\)���<ʐ�]O�	E)��@�(�RZ�{�s ���- ��`����l9`��x>�yN����hGW{�-^�Pi4RQz���zJKK�","��'���"���AY���9"R*�#�(��gɩ��L�>E�_�~�����2����G�Ϯ/.�GKst�\tG��G�����CtԄ"�y9ٻ���ʽw|����XŽgϞ�g�}�z�N?���*�)�@�u%%c޽��k{p��������W�ԼQ�$ �ޛ'|J�&�����BU;�ׯ�����"z��4���v��hqqq�	8�s��[��-�W��e	1���I9��,fF��܌�1�^WW+��̚5�INߓ5.�޿��2�a�3�S����G�R�ҥK�r��7Џ�t;�G BAa���)�O;�*�
K(�\v���<��G_�	i?��/@����r���=x�����L��6�l���BWwG0������O�?_+��0��'�����[�'4���׍x(s�e�.��JJ�Q@�% ς��9{CAݙ�9��O�����q��uI�U�9s�n��q>��=��	���􏋋�/�j�9�	�I���)>����:��َ�S��=�7n����5�\��]�v-���PYI�p�1򈁺���[Q{괬�Ǎ�@UU
֢��[>܌���g�9r�:��!8\i�jGvV.��[���W����G=�9�[���������`�g0�(�@���J�`�宻��~�ر��^��Ç5���S��h1��+�D�� ��e�<A3���N�'��ɧ���z� :'�*��4Vk�`VV���L��8�s�A�q�X��t� U(F0���=$W���r��:��lݺUN�Θ>/��<�>$��5���{����X�h!v��	�Ɉ�{�� ��O�]�>ڲ����v��n���g?�oi�Ν�^�b��x\j�����j��Ͼ���[o�{<�����O�뫮��p�u�mݶ�>�J;�괫�d�6�l�A�3c�U��^=���)�����h4f���^��U��j{�<����O%B� ��s*�T���)�)���Wj�����|�}��~J ��N��'�vKӂ~�!��
�)RJV���1rږ�ښ����~֬Y��_]�<GmU�@���?�&L�'��^p����@��K�^�e˖�n{�N���Gh��;x˗o����L&sY�S��%���rs�d}qk[[��}�����ʕ+[�4<����E�p��M_���)b��gZ���.�?%��+���Bee��c;v����Mcd�U����+�'��[.�S�Fre��R�#�z"|��n�yt�='���E��X5e��>pp�g�d����A���kM0�/���nw?tZv����tN���:���ӀBC]-��Z�
�.�D��/+-��먠/M.����߾�?�<n��&dg�b܄q�Дe�/Ė�>N���=z��'�g���Z������>P&�XB����==��y�����ڵk�}��7��G�馛r:�;/	BN�2��HFEʒn��g�%�B���v�_�-��s�WЖ͍7�8����6�ݭRAO$��J:c���)�u��*�L9&F,�	)+���c��@d�ۭ����B��8��ɞ�Ԟ���:#.�W�:]R4"d
/C ��?-�T��k���5���TV���o�����>�?���<ٓ������4< '���_�<� �͛'o�l6����D�V��fɊK?�٬��������a�b`�#��d0�O����W�ݻ�"�ZCCk$�ágd,))VA�����CG�r�bD_{��555ن��f���F�������+�b�KPH��OJI�u������d��I��_�4�,`;v>o�p���d��
����y.�DC�L�������_�#A�!�q1���*A���n�4�)4tu�b��ݘ1}:Ɣ�������	��F����5��K����~ʴ����{r�@�t���JKK�
�^;v���n#v��{���G�7�iW�V2��{�>���CV����mj�آ1i-d�CcnS֭T�m���Sf<��^��|�u7����j~��عsg������)S2B�J<=ɑ=�� "��=Tp8�r����W|��@��NP�~�n��3fL388�Cp���_�s{Z���7խ��h7�ٛLde�A�7bh�^�L����Q�{�n̝;"Srm�#�
s�=c*TL�M�6MN���ף�� ��RA_<�@$C4��ي��6���M2-Y��'�T���6��G�������_������#���E�y9[`��10���j�7���S�0=�CL}�W1�g<p��(e�`�#�<��}!���W�9AV�ԺrLI���o9���'���CP���)�׳g�,(�5�|788�Cp��8g`��}�x��L+_��$� ��:'Gd�m�l�����[+4B����[n���	;�������GQQ	J�Ɛ�^z�E9E^9y<jNVc�%Hgľ�㏑�����t�6�2�euG�x��݈;��NLX�Ɛ��!���22s�7��gN���կ~�Ю[�uv�\��ݵD��g���V�G4�Ɇ�/,
fdd$㱸��q���0u���>�`7'����S���yQ,&����Zr[��a+\~	���2���H�0�����2�>m£)�S�z��y`ڴ���y���'{�s����q��ַ��]���EW\�X\T��<|�-i��Ӿ�h�M,+-��>w�l���d�&c���fԟ�Cqq�"��/�z�-�؝r�����߿�"S�6��;p�uס�������˕�ꓧ�uۑ��-��9����)��a����_�o����Xв��W^9���.�y}W�Ñ��[��pD�HK���d2��L�Gع�&���/��ꫯ�����=��C�Her���I>�oS���Ϊ��W
��JG�R�OΆT���&�)�y�{��At8�G��2���8o�ɞ㜀-��7��WǕW̚P9ް��@�����w�)��-��ݭS�Fgn�jLY6��{�U�P��0��>~"�_x֯_���Od�������
�V�+�\��;v���F��{���w��u��eB�<y2jkk!&y�?-]����q�;�v�&�7�W۰�U~suu��[�n�x��O*��P���1���hT"#��Z�`��f����3�<����y:��XLH��M�b�����G��(���'O�%��Rz�O�>���O�a��l������ޘ����9�:�B��پ}��)S�}xݻ�CǏ Q=w�\�֏>���o���nG+S�c�k�^�W�p9K&+�WRZ�#㐛�/�����i���B����D�I=u�+W��xrқ9k��
�`�fyߖLv��;�LH7a���vc�ޙK�~�9R��y��g��{��Gǟ�O���Xt�~e/|����bV��bWnPE���On��{��@٫W0:0�`�IA%�fd����N�g�N���{?�����sg����x�,_�Ύ6���b��%��e+����٢��g��u�\�-[>Duu��3�g��a0�A��.�BV��7l�.��ys�y�f,^� ��{�l����mr����_���,\�GW!�5M�8��i����6_4��ߙG�Y��RLpB'���%�V�?�cfH){e����p�]��.��i�*x
��'{��
��޳gƾ-����Ю�r12�)�7s����'pӍ_Awg+Z���%=-�T9O���M�?i�$����eE�w�^Y�_��rD����������l�2��|R�V�o�� =�ƭ�k�+��O���}�؊������򅡽�����p����I��!��#kq��~t��qkF���	Jk�g+��`���}wq�O�����;����9�.��r�{s��N�~|ie�0��d3���	�ٹGEL�0�}��t�mj��2Gd��L��b�V�c��c���[������l߾��݈o~�<���DSSNT�¼ysPRZ&��-��ǵ�	?~�G�|q��J�'�3�k�bb��������/������kh��ș�s���)�<E�+����n�͑	�O��g�>1R�GYv�M��eecO�>��N�g�6I��o]�q�jօ+��Z��%�Bȇ��<ԝ����DSs;����x�t$��`F����i����w֮��jh����.b�����UW���lD�@?��0#�b0��w�yG&��˗ˊ��nwR ���z?��u
_�mۦy���gF"�
"h�"�N	ڳ'(����M夊����(���F���+�Ur��&����'??�{�s���d�q�P_��Ě��}՚LX���ƬU˱�?GɌ�8��F\T�`=#��q�Qs"��S����I��K��vtYz�1e~ACS�L��ݽ��Č�r��땕�ZP�tm���o3ې��d�A�{��k�\�So6�U^>��/,p3���Ng����@�n�]��P������x�(��p8��L:�A
(HT��*�A� y�3t���(..��8�{p��8+��%���ܽ���g3
C'�pD�"a3�]���[��s`IOCcoZ�[����@6T!�6�>EZ?��@% LI��pJ����x
���#����@R�m��n��رm;Ɩ�ˋ���4p���Lf���%���B��А�Ŧ��~���:���33�(��v:��'eOϕѵJ&��+ǆ�_��uu99�m<����ɞ�,�����=��.3똞�A�"R
C���:�Au-�.� �L�ee�ap�j�zxQO�$�^�	�;.��<���V_�Z��ݶsZ^��;���.F��;a�Dy�A�O���36i���.���p���cG���¡1n�[��j�#Cj0*���F��+�NDOY]O[��GDO�t��LIJ�ع�333�����d��C:tH���%uO��4�Zs���d/�L��$���9K.@�͂H�(t&�ly"����O��䨾k�V��'�v"��#���+@�i^y�Ԟ�����.̞3v�,@A^�������S�O?Q�W�LM�`8�P���?{��X,�A��(�4=�`,.&�d�}t˝������r`@cp�3���F<{��E����>8�s�lx��y���n�`A0 ���u�
���D�Xr�eP�co�If=m�"!$e�.Q��*�N�g��+#}� ��ny�F@Br�rI3�(++�g֓�>��]|�Ÿz�9���ځ[n�
v��ӭ3�_q93����8�P|��%M��K��)S�ݧ�녑��B��uţ{��!Z*�����93	O�������m�ƕ����C'{�Rs���[n��O��I��$���[��zF�Lɹ�ʱ��I��dZ��`d�uj�7zbX�I�{�
#����&	�j?�'/ --is��<q�ܞG�:�+�J�\���|������VpS�/��պ_?�����풧8��w
GG�~��rL9�*�[CI���k��~��<�ō�EE��̙��+98��ɞ�����K���U�'�N�#ЙL�"4Z#�l��(�?�:Zq2�C��}(��Pz#n ���0\C%@.ؓ����]�T:-�X��555�+>��V��b��y�54���.\�$���9}�̗K&�����ngoo������ �q��՚���хy��:FirK���J�>�W�p/9��?<�&�7���򨷞gr88��ɞ��Fh���Ck߽��?X�Tk��
1b�9S�l�����L�;��!Db��u\g0B����@���`v��~��N�2V�PJV&�&���'Ґ�3��j�Zv���U(��G��CT�o�K|����t�f��O�S���;�L�B�D�g��Ϙ�|�@�@
�|h�^5<��@��t�����ᬀ<�^dǏ���.ppp���=��W���ˮ���fJ1����0Z�Q$l�b��;o�'=���!F#@B�kS�*j���lh��T�=[���L�f,蘢��c�PF��HL߱�Ȕ]\�����ǲi����/��Hz���/[sǚ믳����c:{�ҿa��?�j����S~���䀍�9��)�c$��M,̍ F;�Q����H�ç�J~,&ʯ��%��A�V+W����e��)|�O��=�߇�5ى��k3I�6���^�c��uVjC�
s�#$�ň~0�`1��cu<Ĥ��Խ
��\�'S��)g�Gi�4�!1�Q����FRC$����A/��{Ŋ��=z�U�Q��O�j�������_�9}vt|q���C���Μ�9��Ç�}=sC�U�Ǖ]���+��	�$glFϲW�ut�2�f�^��~<�w����z������O�sp|��9�fH������W��=�J!N6�v�<h-�I��@�S�-A�@/��7�:g�2%�f��Lɋ�f�TU�'T$���ר�fO�,p�l�g?� ��z���e��8[����r��ɓ'Q�8r�
���	�Z����"-7����Oݭ2�]t���Y����{�ر����e!#z�o"�Z?��J���%�S��Iœ�흟��OeJ˝V��\�텅�����3�d��7�����ۙ��z�keP��Gധ�
 �S�g��:�c��֝;6�bĜ`DO=����s��W�-zqUR&�$���r�32r���iX�^�8�=�֪d�F�6�	��=�9u
����s�6\0m6�O����`����nn�̙��G�K��~SIՁ�6o~f��wpg�s�7�|S��ƍCAڳ��������1}�D��~{2���[��=�<FW�+A A)̣`��+�����m3gΌ����S�d���m��oݐ�HV����=V���5�ad��q`�ŋ�Q�I�L*&�#"tLz#F�D���O�Q��S��{P�{ME���|� f�I1I�[���@��g Ɨ�`���x�g����X ��~�^pL�K�u�-p�g�tga$��u���Ꞓ�|�p�u<�{���t/Ť�T=)u��G�ᐍq<y�"T��</�h4�-w��=)w�����r������pEEE888���9�6���	�5.��鍶pTN���~d8���1q�b����ڷ�HKg��@�w�w^�Rs��u����*ȣU>A�L���*�u�O��O�E��C��:��}������g�Ñ��1���A�tv!��@���<����A��Z���;��:���-�vl�z�C�c��hgMMM�b\,g$/�)mvr�]�!w9s�E�y�n�#U���1*u�yL�*�|�^��uG���<����p���ܐjwYw���s��"kB��-S�z�� "zq� wȏr�c�����ĈVԨ�*��|#|�G�9r�=��'�i��s*آ�-#����Ħ``xO��� ���O>��CQ������Ѐ��t67ëW�{?�!tY.`h�������sĤ%t�X��(�qV���lx������L"x"d�g*?U�'��E�+�w�IN�E1姐��#���Ϗʽ��ǈ^b��PPPp������98�8�s|.H�6͇w�p��M��R��]
GR�eL�GĘ���q��SV֝���h�,l��h�XfS��\U/�"��*��/I[���V�Ĭc�@�q�84j-S�z#AX��3��p�U���~owT�\,l(r����uj̚;��hRR�׍�]����p]G����sU���А���7���GG3�������N
R�T�G��*U��<{��0����S����������5����H�]t�_rp�yp���\��>��Û
U�<Siq1�ɌHRD1h�/!��,�ۏ�{��lVL@I^.j�C�E���nA �{�ML�",P0kHHt� �>k=��1��0,:-t���c�M�I�=�d(��9:�,��K�� ��Ӎؐ����1��1�T����N�����͋�㬁��cӛ�[f0BV9��NF�vtu��}�Z�}���|~y_^ٛ��=�V72 �������9Ԗa�m�� �p[qe�888�,8�s�U�����͗�'�<M`��)��J@T�"��h�������i0�M@�o�?����\.HYd��@�É��~8Xp�6j��c|�m��-⌌��I��$t0�{�1v�9�����,T,(�aJ�X<����R[3�r�*-��
�$���Hǜ�b�[�Q^���<l9��������3���)^�v�}�v۩�S+X��Rᅅ�2a+�x"���z�T��J�+&:J[���?zBc�'�s�++�~��sp���d��ױ?�V�ޖ-��#
C%����O��/H���*I����d
�����z����"�����%����N����q/�T�F�jW�c�}�)<2�a�{�~�6�A��a˺���u0�i+ S�N��x�X��F|��������a�9އ
k��ڋ���s�?�������_��W���I�wvv�[1f�F�CCC#=�"{%�����B�)�
:�#
_1��¯�=���qp�p�����2=�{�tu�K��-�1F����0.f�:�Ic���n1�֞~�ldk�����(!�����(�Gv�X�XX�Rn�a�S�4�\5<�VE���������qX�z��O��&e���`a�O�$[V=t���ցw��+�b��DK��9c��W��ѧ� MMM3���'{\ڟ��xrϣ��˙&��w�(y�hW<�9��+����s�)(`_��h6�*((����'{����ߟ��]-x}:���9�ŊPԏթ��g�Z��`1�^c�Q��MG~A��Z���1A`�^��5-�ș6	j� +��	�!Ђn���dG=2ۡ����\�p!|�	����0��XbOc����AE��"��q���p����؄���Q�s�Wn�$p������>˃>��������SjTYOi�`8�h�
���ߓR��(���l9��j��۟K�3§�����N����/��=�������/`�]��Թ:D��{ �Mph�SU�4�Fk4˕�RRD��
wk�ͩ��*��=6j�B�y��a��) =��t3ә:�B4�&��x��(W��F*���*	�5����?����*
F��I���73�0R[�����$.%`�X��P����3�.��c��������z{{5���)�Ge�&�N��������◯J���4���z�v�鴺Ccǖ�L�_'{���{�N:���/�q�[b�x%�dp�Qä�c�)i��OI{bQ��Jsm0&t�GDH��*=��_oЋbv]9S�C�����5wCJ ϙ7{�S��Qv��d���5uZ�ю]�����D�]kW1BOƐgʂ��65iEĠ<(�`���f�A�"���oN�;�g��պ�k�.bd^��\y��Fؒ1�R��̰?3�N���{�d3�g��"{ń��ܜ�����1���+�d��g!�Y������egRS�FF�l���P4�|� kbq��GR�����cM�j!2�ՉL���b6 ��4F�1�!���x.�����/�@Ʉ	ظc+z���QT����]Vڻ:��S ��j��G��Y��5B!�d�&�� Ea��b��Ϧ6�Q��vњUo
K��V�s ��Ӛ���Yi_�]q���ϗ�=�u(���S��Iy?e�ٻ�Կ�)�|[�J�J��f::mUIY�>������ɞ�������
5�����S�M�g�Y0"�Ң������ς���>L�6BC+����� S�aP����:�M�A�&z�C����6U�����@o7�i.L�DiE)�l�/tf�矇.���>c��K$���fo��X@ARJ�j���}.�I7d��]��[���K�8���H�x��~o`��l�z�>F�є-�J��������@�A�����Pz"h@������Ke�=����j�muu�v 9�%�ᴾJ�9��ϟ�	��
N������~�k	i�iL��#�fG�٠ż���6�V�q̘��OWcǞ���~���ǔ�VH��!���t,8 %����8��j���?r�j45��qX�T�E��ݡnL�1;�n���q�� �mv��503bW3��	*��г�"�f�6k¯�\��/?�U�9����c� Lu}}}�wL�(}���%�ߩ�^v�Y!�R�r�}B��#P�eZZ�b_I�Sʞ<(�O���){��<��jݙ���_'{�O�))����䂎�ǖ�B!!k�L_}1�ڴf��%�^���VXCa<���`��9��و��|x:{��ur`�j�`՛`�Q�w<	��d�������|=x��8��g+<:������]�]��0��`6��>$�	L�(�,�a�U���� �eD@%�C&���ǝ��:::�n�g��Аa`` �!�<��l5�)|�����<�Q�&���*|]<�G�~�.bo �2�^I��[���ugd�6����s��=ǧ�޸%�z��[��d~qI!�LmG|�șR�.1���}͵(�[p��wBm1"��"���I؍&�),���qh�@��c&�h,��M�̠��#;�ZSu��>{z�A���L!���Ƃ��<���(�O��&-
�f��F사��	y��D�B]�3�7���ԋ�87����
��en�[=88(1畔��U���N�����^�W>R���SE}�<g�4g�YO��Ba�N���4g���9F�Y�/�ϻM�f�u��4�K��LXz�L��[��>fO�D81Ȉ݀�˖`�@[W����B K~�L��ۻy���A\s�W�Hwb��c�H�E_,����@��G���ŁHЋ>������^FN����q";/G�b��	��Z�xL�ۍIhi���5[��N����6N��4���g����������{'%N3�+**�Q��5�������v:

�ј�GǨ
�Η�r�Mt���T�~D~�j����1%k�ϟύt88>'8�s�����	����\s_W;��ۅR�
e���l�����`u2u�`��	X�h�����@���L]k��Ű���x�&X�
��`���>F��	�%�Ȯ���Sh�:�XR���e���ԝ��F��Aw[�B�*����42D���@Cu���$@��"&J�1�0�I�������>�ܡ��.���w���1�����X�UTT�����V9R��§{��e�i�aJ�S��<a��^��'�/ʩ��VM4�{Uiia-888>78�sȐ�3��?�U���ѤE��J��(���7�<#T��ɠFg,�~��[Z:p|�Aح6\�8}�[�Va��8��=#�0[����F2͆��s�Q��Fğ}WO���l�D�TŨ� ���JMM�����S�F�Z���gU�N�e��$S�b�ݘ�j4R{8�b����۸_�9#b��?<�=�L��,q��-f���ٽY��'������zGEy
 ����R�#��ܚG�(ů�j����&L����N�r���~<��P�-%�� �� ;�P9FĞ>�>x�J�J��7�1S'�����S5�`ϧMC�g
~9N?���A��"��Bm0bWc=Ʀ��>v~ߐ3'N��7ބ��Xt�7����b�:��)� cn�T��Խ�hE�N/���%8MVH� 4:"�ӳ�R�C&���}��M����8�hii1755�a$�Ni����8�)�M�N�{�=�V顧牄��ixJ>Aq�S������u�Qppp|np�� ��2������*]���|�-��p�Ɇ�����֏[���t
ƌG~�x���W�c����+��f��QZ���v4>�lW:�����3��׽q�D���3k6��i��ݍ���x�ې�*X���12��$�E���L��XС�@�f��@�����{�&F�XF�>�Vl��̺n�Z>��ܢ��7��ԁ�-��Y��gΜ)��yX H{�{m��_&te�-�Q@�^7n�l�C�S��T��b��l�f����9��������ɞ�ΓS�qq�ZJ����� aa���=�x8�>1� [��-� N� �GN������8r���o1a�8l��#T��E�Ǎ(Si�������?"�t��\H�=�)������ً};w�\2������� �ՅH ,[�j��Qh�$��sM{����4:-��<�'�U��c_���o����q����:�)�2�ۭ����^XX(O��[���z�rP�L�#��Ey����H��ݏ���=�C��~v0�t;
����������<��k�����b$\@��^���:�H9m�}lq�9��ӊt��|���L�(��`AA7�z+�UVⵗ_1ce��+�����xo�n��]8��C��h�p555�058�nDYE%$o ��2\{�Mصn#�-=0	�bլ���h
�-Fxt�����X ����OY�_����㜁��|�ɋ����-�����|�
��~7!@&y*�#b'�V� ���i[&I�U���'�Oj~4��{���J-i5����������o'���j��Vu����,	�7^���߈��&a�r|��z�{��j���/��#G1�r*�}|mu�h����d�H��/���HӚ�n�z�U|��;�^Z�G~���b�[X���p�u�aΤ�8��c��7�=0'#쩫/cA� �������l��0�+4�~z*�X �`�d��0��%��C��kgM�U��G��bD����ƾ7JߓBW����SC�H�������P;&{���H�#!�@��>�y:GI�#�^���m�����j��N��1b[��7��ug�N��^RӘ���Op���W>x��ړ�<�����`z6�z0��%���h-z<�8q�����o` 3'O�ą�_�
�ӎM[?�Vz�z��Hǋ/��1?�n��x婧�I}�4��r<�UG�Iu52�:��p1B-��8T��'�F�D��S�Z5�L勌8�ZU|@�ٿ�꫞n����C����_{�K��x!1ͫ��͕�܉̉����<�H�+�{��)}��*_G�O磻�	�>é{zMJJ�`~~��ٳg������S0U�:��OC��9���+.���U�x��[�UT��>�f�(�b���ـ�s�c߮���-���fX&O�5˗�ԡc��_�D ��x.n�X��\�eW_	#i)�D<��-�R<���짰��(����_��~�^?j�;7�P1c:�w4c~��d5"����T�q���Z��,���̛3�ŉ�=և_��Ξ�����c$b�on����e�N)yJ�S!��Mi����'���b�^ޫ�L ���ޯWz��}Rs��O&.���	8ٟ�oښS}���6���z��� �-^��;v!O[��U�p��	\�d��!h#X�����F8���.�D��{�+�QB�m����Ow�D�>���`�"���b��&��׶����k�b����e{��i�:p�8#�/!1��؏V'7֫9���x@%�X8s/��>��͵k�3��w"tJ�+�xR�}\D"�����%Fz��:R�t�hO^)ʣ���^�[OCrT*}Ҡ����dt���'��RU���~�M����_�<{*r&NBҠ�����~���o���P6�^���]l�N���U���%�k߾��(�&uf���d���7�E$܆ۯ�e���������yyX��Zlٲ�y9�����XW_W7�L���6����r���Ia��~2�($e%(%$DTj���i옷���6p�kh�n�����ⶶ6���YY�:w:�2��+3��\|G�@_o�������qii�����ʜz�*��������+�u��^����w���y�jw���o���j��b�}r�A��O��b�PgZzZP�g��K��0������0Tx��M 㳛�on�L{!�?73[�?�P�т4�f�	[�x�'0�����Ĝo���w���^u)kj1�,l�pfWNFz~�N���ff�����C�Pn��SA��O� 1"����btˢk�	�;O�c�>}:���a�{�cѨ�L��PQ1��m��v�(�n������o���Co4�$y0�	�$/Z�a�'��ק�xD��>�H	xR��(v�)++�U�'8ٟo8y2�cϾU�,�\=S[*[��*4�؋��.l�څ���Xq	
33�t�&�qU��B}}?~�ċ����?BH
�����g�^�k��
'ƣ?�	��p�b�lJG�������t9d�w�m�w�t��@��[�����cժU�� b���FvZ����B�A�R�:�ԃx�o��D�C�> �s�}�Mlio]�ZG�u��N:�ꉔI�S��q�nw�O���L���6����"�{e�!��O�x��k옘���w�ܙ5|���N��H�<����5�;z���� m���0T݈�����U�P>�'��ഥ#&i�*3�;�Ŧ��C+d���ٓ�S�=|~/l��hh�E�`'�ҌX0k�`�!��0��D ߾�<��S��DB~X�b���19];{�,?U�9� �Ȗ�����֋|��d��e��"n3�"ѝ�gL�v_ ���-�����^�7�=�(�:,������S��R>�t�le�B�D�t}��V�]�@!{:gxܭ;/;�I�&�*|� ���#t��V��'��5;,f���BC5�j1�`������S&@ѡ��1��M�Z>�����Q�h�F=MZ��'N`FY�q��Ǟ@��c�2�����^��}�ǞaǓlש`d~��	D0&���9����t%B�A��&�p�0҈S?}�$��3�cq�j�3�pN�\�U�x������\F�3��7����a���#S����	d�C*_��F���\��'(��}z���I�^�:���/��������<���c����K��7;ML�ա L�>iR"�:�lF����(/,Ee^9�=ܭ-w�1�t������/�3����-�^ܺ�2��6���h�sN�	S߷��m8�DٲE���{��r�X�)�)*���߇��&�{�#����Xy�J�@Yz-������дw�� ,j�ܺ��j���IsF���K�^���v�=�
���_�
I�+�m����"{E�S�>��Z�f#&DF�F�/_1�F+R�#�k4��V�=XR��	�����b�-;K���%Y:�Z����OF�=�=�d6�
P�J���;��A$<���"k>��s�cby1�Z��r����E@�#f2Q1ס�i��bHC��jh����a�X���E��=����|Ҽ9h�s@v�[��+�XY&��WX�8�����dd�E`4�JH��e��X;��+_��s� 8�9����������������Փs��O�T�O
����>�B�t]zz���I����J��p�_b���l�*..����'����6.MvtNP��0����z�x��N�D_�&O�-��.9��#����''k�S1v��mMx���a4��'�Do�������NǬq����K��Y#�~�	�5����ݘ66}nDh^��͟���L�6��;�y�Mٱ�fzB	�1b��}�J,�ю��Ϥ�y�]e˗��8�-(Pܽ{wQgg�l�ۭ�=�hf=�Q�='�&�O�}"v�=�������@�7*�@@i��_O�A2)�ߎ��&�;�^�������y���'�������FZL�3-)!���p��^�ńc�>A�� Z��0�s)�O�q���B�_[�n�o��Y\y�W������MX4a".2s������WA��Ę��x�n̞:�FZv�Eq�3�#"����=�
�	���*�`�_+���#b��%�4�GQ�k�ҥ� �h�k����Ocd���<J�ɤM$�8�QQ��O)��ޙ�����4��h?|en=='�1���t����z�����!U�Y����K#�1i��`��*��bf\��������a1��]{b"
��_��р�3g�^X��<��G�`�c���k��bÌ�q�ho��(�eeX6c&6܏����1x�/c܄|���6�_�ߌ۾r,y���">¼���e���GN��ߍ�Ph�tZ�=�ظ�7=��cX��t�՟^�H�^__/+���rdff�dOi{*�#u�<&�'����'~$�I��^I�޳��t��d����SY9���>�Y '�b0��Ş��3"�i����C��j2�PF�1O,+S�#x�Z�*B���iC0�Baa9J��Ǳ��f�^����=l��́��N,[��]hb��Ѯm��8�݊L���dӦL��7�FwW��>�Is+�;6�փ2G>:��P�h���K/ƲK/�{�y
��hUzz�����Y��ma��!p|!h�oɋ�#��n���oI�ggg�*]������2�F�E��v�)�)z�k�=�{�N����ƍ��g	����q�x����>렻$-)A�A'haЛ �pGEY�1Ro�����ȵ-ٚ�e��0��uڏ�������";?�+/����ɝ; t�`�/���3/X���BŢY�~��������Q\��?X�S�w2��=�_�e
.�H<����x�-�o��߾q?tV��%��H�H�QuI�{sy�(~�8�=h��G?��<�ϛ�����Ę�SO���>G�M��j!�L�K*$>��i��T=�<Ai�S�U���	�����g��Y'�RЬ���~�����%���a�TjyQ�3"�ZlLF�a7`�M7�Tu�v�Ĥ�BDݽH�5������C�#� 
C���UR��� �N��)�J`S���?���R�3,hcJ0=���̂(Űs��2qԒs��@$���'|a�v�AҐ��h?z[7��%��èCw8�2��tWz_:::��4��m�<��6){"l"eJ�+xd�C�F�^&~���C$(d����{�5�1�cz}j�����	�W��q�����{�oz��;:���^�H�J��7E�-�A��:.���a�h9渣�s�ux���K��?�Gw$����-_�ӿ�d�Βb@-`����N?����׭��GPs�8�����sp�U��ц��&�X8��YH�����ق��?��Bxs݇�����w܇��0����Z�x����xz�S�����q�@�����%׺��܁��)���*�P�}^^��ꉼ������
��N7e/�������ze��r����G�(}o �Q�������Y'�B�-n�W��7Z&��զX6�����V3�z5Z�>�N��� �p��7�Y�|�_F�ı�)-A��=Luo��f�;����5UL���GIn{�s��p��	fI���م˦�C_� ��Z�w}Q�h3;?��ӽ�����i(�d �]�`�|�nSg'ˡe�޺�+���cǎ��m�6�����p��������˔y�=Wmܸ����񝝝��<�)�*��8�Y�~J��?�w��Q]VV���OOmw�:�Gקz��=~��2ҷ���v���㬁��?!:�z+���A��봈	h1��"�*5�� �qyXx󕀉�I�������L�Y��J�1����aӻhmk`?s�]����۲�X�c/^L��o{7�{z�%̜8	S/a�Ϗ=�B�% ���)CGM;�¨(/D�ۃ�ن�ieк%l��K��7��5X1s.^[�.R4}��S����,����6<��=�q��p4Z��N,��s����Ү�.;)uR�D�d�C�����b<J�����Z����:N�Ai�S��z�H~�b1��0qҎy��qd��N��d [ܷ���[TuM��i�*C�5[K%�gu#~uI�}�8V,����ٚ�4��	����ʟ���
�ܻ��n����]���>��4 �3Db0yp��4SyQ���tL �q���n�Q��@<�̂DX�0�G{U=Ƙ�<؁�r�/����Ħ����l�M�ok;:���7��1p�50�����?��Hz#\��������>Id�HY�T��t������8��RiO=�����{z�L�S\�"ј|�*�)@����y��Iڿ��}��)y���삓�?�z�㵗+���\3Q͚PA�D2��V�[�@�&�q��qх2ы�	�8_p�%(--ƺ^B�ѣ�dz#Al۹�p�K/X���+Ͻ����5Z̾����n�GGWz`wA�;!&$�[���Z���GQ�*��=��?g�sTFHmh؈y���3 �Ӂ�Ύ��.}vQQQ58��w�w��
����~&��ࠟ���_{�e�Y���s�͡n�R�T�J9�
��%���#6c0�IM3�z�a���E�����4o��al��	焓d�V�\JU%U������;��.z�z�V�*��Z�{�'պ���������8l���I��[%��!�!:{����!��㿱��.%�X�ϰ��0�e:���ZX���0�W�ul0�mt��r;�,��ϙ3Gj��#b?�8{֕>v�C�3��4�4���d�)�[��!+C=,����D?�P��vP:�$�h����ӕB����!��?����/P��"7���i�[ۨ���ʂA���k�]E��,�'�C�G�Je���4MM���P?��'��5���Qf`����-�3���y�Fz{i~y�*���Оg��ʊ*�KgR�������'��},K¥Ĺw�����/c�5�����Y�v�|��W��}b;��|OO�q�4�O���F�ά7K���z�����
uҩDa�*�������-��ID���E�x���ñ�R���im�-7%���ӵ��K�UK؛O�����Ѹ2���D,L%��t��R&����'�+��#���l ������*gϝ�׬XES�Az������!�ˤ�W��e�����T�fD�����a�h�b�Zn_?�n�@�	�-�ؔB��r�s�(���Ϗu���_,��@�"Q��vx�e�L����qu���W�8q�P�h��0��s�QZ��N>��[�������p��|��c��g# &�!��}z}�n����w�M��@0� ��  LQIDATsŊ��I�K���$!����_��5�CsB�������S?{QC��/��zZ��������ƀO�٧�y�����)
���G�-]��^�%�fO������ƃT����}���(�?DMQ�/HiJѵ�L5��Ɩ:��+0ClP��4��GӲ�kخHRWo?yY <�E�O%���|����ߋ��o��m8F�E�Һ={��fa�5�n	�BS�;�������ٳ�СCt��	%�p$��TU��"���������0��� �_^fGk<>�2p.^MӮ��!��p=��1R]]�}˖-��ˀ��$ ?�g���6FO7����R��"�}���x.M�,�g�4�y�z�_qJ9�Y*ğN����`L(˥���5{b�l�L6��5t�}�<l9�;z���I�h�k�+�]�ޠ��ar�24�b�Yu5��"���s4���޽���x���IM�C%?Y�,y��%�aQ4&����|��D�u�]w=���^�ԧH����]����%�Y�+X\���
����o$6T�{�G/������N��[@�H��Px��%���W���I�PI��Wv����;���Tv~6��7o�!I��˃��d�ĉ��#Goo����X����)�f�=�6���"�5��|�r�)U}�ٵ'���^~	%Gh4#�iQ����o�1�a>�^W�����_�7z������OZ�y{����m�R��G	��k�8r��}s�>
yC���;&�D�`qIE��J�!ᰔ1��`�}��h�k��Ŗ�|�O���g/�����ֶ<|�ż��oCy��o|��)%����J�1Ŏ��_��WJ���o���̙C/����_?00��v��iǚ{��n����=�RWoH���o���'��վ�h�Ɠ$�eA�~0����]6�EcN�2��i8�\(H͉$�yt��[�f�`O*O.44�)�"��y���N�J�Jes�m�:ڤ8C�_B&�FF�����������l���+�k�(�7���B��)t����T��h"M�N�����)g�u��X�S�9�'��-Y�z��Ĺ[?��w"�Z&����=�����Ͼ����M�FǎS	vH�;x���K�9��a��]�����8���򇱀P<^�eo'�2�����~�z�l��>���H4J��-�I� ��	N�嗫~������'����I�(��R�=�c����{����S�ǷR�ᤜ	���p�L����h0.�?�}~{#p�œ�yK��K')c�(X]�~п���Q�_���O��wSǩfz���<���$������ө�����oQ��O�d�����7	cv1��Ea6z(qΚ�����p�����`Q��[� �pdΣ�-j瑅�	v}��/\�P��Cԯ��5�]��wq��7Sgg����w�믿N۷oW�#C.y0�������������=�C```�Z�x����-C� \rD�'0h���{?sO��㆔a9�^9��=Yy�d�.]���}yׯ%r{	e��0)Ͽ����_�ŉ=�pL�Ϫd�DJyyx������q��}�G�CAʲ1O�����t6=��o�Rt��7�%t7$��?It�Z��f�:���O�\�\�,��>6*���?���E����y�������[�ûH��=t�6���YAv<�� �H�Ú<������_�pA���Ϡ���J���ÇU���Ŵf�jl<BK�.��Y�h۶m��oniQb?{�lu]҇�Ó�T<?.��	@�����l��ۿ����:u��S����'A.)"��e�����i?����b5�=�P2M�l���-�5}�FJ��q�ay�[5[���R�_?A�������v
%���}���X�M��s� �\�M�]�Е�t:):<Hފr
Y����W���C4��EK?{��G��Mǆz�'��),�x���A~+gR�a�p�=<���?_��C'�O��1<<<�_6�߉��!�\x�X�?~��d�<w��9և��[�ѣG�x�-�Ў;�{\�g�Q�"o�ʕ��ׯW��+����x�X.@��1#��*
�$>�27�:����MM�������_~������{/� ���JW����?zGo*v��@���RG'�3��3���9�O���"�=)#ς�!u��W��kQo����=�0A�����̤����w�ʧ��ھ�W]���e���"���)��Q*���y��r�Z������%|L��z{�r�B�v�*z�����|��`P��clL$|�|��s�_���n��"Au{��ث_��gx���_}�U��~��i·�_w�u488�߽F��XC���hT��/_��������vr:���tZ{# �:�p�wܡB��<~tݛ9c�J�;w6W����Q��Bk]���YoY֗�;z��}�_���y�m�� ����W'��vs4�ʬ5�C�UT;��Z#G���o$Wm��اJB�;��2��S�L���d&����>�y�Z�|)���>88@������,��l*�Q�yND
�ȉ��T:�B~r�}��&(���T�������0�z跏>F�/���Z���R����#M��z�B%>vR*^U���~��K�?�L�aϺ�5�e��G�_�d	�8qBy�,�*K���6�}���ݣ�{�޽��7K��a0�:0 8�^���	{h��0��?�i:r�Ha ������x�cru��B�}#����)��g��Ç��i"��p	��`�k�_����t��Y�M?xd�Y���F��v0XE�7>�D/<�,}�O�LXwO籘o(�p��Zy:N������<B��ϥ��7��u��H�Pr�|6�T?�&���,��	U����}i~�c��x=��/��S2�!��K.��S�>I��!�m��OM���J+��/~�v�x�̝�o���z��}�������,�[X�}w���<x�$��²�J�g͚��>^�T� ���1������** 1ǵ����k׮-v�;y���QPYQ��0n�m+=��������EK������2�.Ke�Q1ĆH�w��]����h��U���Cwgۺ�۷����9+K��sӷ-����c�G���iŵ����h��k)P]�����cI���8/Go���l�J�D��}�I��RE��E���p��#3ȞJ/,�R*���Z���x��$KYexY�3�]l8B�g����)�w�m���O�}��x�q���6����K�ϛo�wy���ܹ�$\4��F~����v%�yd�#�%oȜ��#	k�0ZZZ���HЄ1��v$�uu�(��x��?���:���# ��~��G� iɁ���'T���?�9��z?B�3g�P�#�d�f��{aٲe�$�%A�~��3�]����?�ϝZo~��[��_A�h�2����fh��E���9������R������%"�f����Q,����A���4��V�C�c~��7i�S�Ӓe�PiY%�.x�9�����(o�?�d�D��z�d�q�$����G|�{��t���^:�{/mٴ�FF#T?s.ݺ�vji>E#�H��L�}ߟ~�uc�J)�����D���\�����;���3�D>[D�͛���Pbo	uC��08q���UЖ-[�10 `4�S�z��C�V@?��̝;Wu惘#�F"��c���6��DO�J�{��w��+W]�B�����7!��	F_w����ӱn�*��Q�$�%c�A���z�Imn�����~x>��e�^8���R"t�M�/kR�J�N�T�=��E�ۥ��t7:��G�В�+���=�ӭʪ��4���G��q��=�L2A��M���h�|�<�#I���+tӲet��~Z�z5?v�V-[K�dJ5��s�Dls��V��R�K��L���i;�v��%p�⏵y���:=�z��F�^{�J����?�q�M���U���S��'q�������V����7�xC8��=���qH��Ӄ~�n��f�������^on������9���`,Y�������HOOo�ʕ��O�9E�Σtx���Mᦓ����i
%(�P��;�w�E�~|+���/����������C������ZO��A��%E	�UX�������L��.
JiZ�ry=��G�]�W�o�$��8%�#��!��>��G�{����
yN���|����Y�Rqz�׏���5u���/�{�/����-�Ҁ���g�b�~*^���X�;��=xƩB�q��D����[��&7�L�>����q���U%�!L
U��e˖з�����?���jI���F%��\��\|̹���u��믿^=��0�n�q|�X�7�����xꩧ�ŋ�	��Ȃ \4"������}�7_���g;ܞ��]0�q�^�cx���Inv�=C#TOn4B%>��:�����7J��,��x��;L��>��w��6����/Q]i�DGh(���=�l��L���p�������jP����;���#JFh�L3�ycUEbԴ�-jm�G���Jk/����g�~�Zj��7䣷�t���#$\�s�d�z�'W��P��Y���;���ec?�k}d��sSS�||�Z���mW�v|��C)���D��>�|��� A������ܹ�zzz�}����jG�����Z�:�=��c�ә�����?�8	�pш�O0
^����3�-�H���g����_?����P��,9=�]FU�C�l�B�rJf�T�-��H���ұ�MK�Y�S�����4�Y:wp?EK\��?�3j�YO�L���{�q�A��R�C���əs�af��uQ6ɟ1�6�?��m��S��#���R�R���3��~D3gэk���#;<kN�O6}����$\<(�������k�k7�q���|��k�k캄!x$�A��Y�s��"FX��W��#����nR��{��GR���GT �A���X:@�=�G���K�Z?Dp>�e``�.�J�?������� ����b��Q~����ytǶG~���=?���/�9�n�tF�q5���X�D)��Bn'e-���)H{�.���hw�~�M_��FӖ.�]����A��뽪�.O_?O��i'�9�<j6=E�t��Q���32�������g-a����:�K�\�нo��D�H���~�E���؀�C�!���!�h��� ֺf޾nm�����A*,Pr#�r��qm�5���;�nܸQ�cy K������c�y`ƌz�l����.`�����u{�$����I�� \"���M���;5uUg�O������y�����%�J��94J�\�����)��L�)Gy%���ᗲ!O$���-�6�/��G�ɯ|�zs�7L��믣�e��ޡ�T֮����s7_7Of4J��NӮǞ�3��2~<:>/���=<d��a�L��lx�3������)	���썯a!vA�5���$<�-�� �{��#�nѢE��F;]��57�*ϼ��L	9�4���Ã�~=�߫ɉ��D��#�����C�-u)@8���w�0X<OY<��F2 G.�I@!���?��._���)/m{�ɯ�F�+��ndh��磜�I�In�aMb���N�{��=���E�a��#Z���/�N�ۚ���OK�l�T.I������g/�4�d��N%�D�H�η\��om�� ����I{�/E�	ʲ�����}���7� ?ޗd����n�S1�^��^!���!�]��!����GX⌵u��#���������>O����j��{�z� "�`����ذ����m�W�>DQ\y �իW�e<�G� D!��-h� 	��p���O"
���/�=������x[��}m����,WI%f*<L�T^M�˲6����<{�喛v?�"UMo�ֶnJ�wR&ߙ9r�X��9�N59/�tP���4����Ҍ�s����F���}���=�t,���(i�mhd�������Ei�r	ao���q�WϚ�Cf�i��IF'�A�!����e�G�<��^�5vlX�G�[��!�f��q!���x�׎�yܫ��[�K�͛7�ny��_5gb���{�nu�ҥKURD_��{��:	- A�(D�')�����?�?�'������xd�;_���ͫ����ϳp;rgs*�ޠ,=~��ĩ��9��G{{��⨳�<5��ea@�d$N�@������^~,��ڰr�8r�2�M�i���P8��t�"�>2rd����?!�2���,��zx��c?^!�z6�ܱ�������� C��ec��n��Wd��ٳG�GT ������#!%ur>�	<^�����ڸ@� 	z0& ��40�:B��� ?K� \"���BRS7�n����~���_��T���ps�@"QVϘ�L��\��.'�Y�=�
��w�������t��>��_&�/&?��S��0k�Q��s���M�L�Z�3�Q=��r)��D���p����L�����ϐpi�&�9sf3�w=�
�Z��a�w��:�Iy}=nǡ�^Q@����,z���X�����Bo�ٷ���<��o�Y	<��`�H؃��8ϴp�|-���q:��}r�x���W�*}���� �?���ZX��v�x���Oٶ�s���ٜ�v�MJb��;@�X�L�)A?u�Q]����6ү���h�֭���O���s���E��ˣtæ̈́HAogY�~�u��	r���_7MV�����m_���|I:�]Z�,���o��B@�ސP��ا������b��;2�!Ķ?U	9r/�4�s�a ��!�il��Y�z��� ��!� ��q�7������m}���u{��1#A.�}�!=��e���_�u��W̌�n6ñiN��0�)#��7��Xx��,'��hv��O�������ђ�7���*zy�:�����VѪ9�h��Ô���@	��)��|�R�}�k���ύ�����K�(
�ϲ���6��}x�j�J�!���3��c ��GZ�b�s��䧔���wc��x�b���s��/��'�T׃� �F ׁ`# �	��&J� �ol� "���B��,�����l�A�hD�?`B�a޶�w�9iz�g��O75����(�+����4J,7��}�;:B�(�I���㴯m�zM��>�Ij駇��_(�NR0������!��hǌ\2��2�Gl���}�ÿ#����А`��Q�JY0?ς���b���Шk���d��T���-�k.\��]��}�X /���ux��q��<��5���C�`Ŋ����Vw�h�wp��#��(�9j�Ø(�*	r�\�T �k#A.	"�`��sG����z��s�������}g�r-/'���Ȼ{U?�
���dR�2)�pS6��$e����r/�M��!*���XW/����z϶������Lrp��OR{��ŽL��F:;;�^>
=�B�����	�ZO��	sh�OB�p;��!����	/�K� �ا[�8p@	��q-\az܇������Z�Jy���X ��������2*	��a6Qe����!b��X�a�����?���x�®׿���|���{����@I&a�����2�I^G��"ar]�_��]z��)�~�}�֭t����������ٟ�UVW��3j_�������M�Q}aA�g��u__�A�f�y5�"!��B�N��C�ui�}x���Q��o�>\C��!�ړ0 p쐑�ux���l�� D�^q<�A�!�}\�/���YY����p!�D�K����0/��/�<�h��]����ᓻ��}3��kj�|�ᘙ�')ef)���P.M����7��J?�գ,��p�����t�L3��f������}�1Zu��6��8&Y�/��v�3�9�Cxa ��j�!���Gh"�� ���G�g��ޡ�u$�a��"��=B�h�c�z,	�hx�����V�����O��ב�}�� �����hw��gI�K������/�_~��߹u{���w>���k2��~�;�_�STZWC;������J��=���m�~�5�=0�8k�M�I���Ų��w.D]���g�b�"��@��G�>�w�̙�y���ݣ���#�8C�u=�E���k#j�n�:uMx���z�
�#D�\�Ë���t�觼n�!~�$�%C�^�71�n�D���m�.�q�����~����{�\ޙ���7�[i�U����(�?�&�T5w���}�FC�0	W��]�о9*��.�U���Y�A��k���n��b�'�x�[��M��s�*!>t�(������C���wTI�p�ѣG�<����: ��� q�3��П���9á��n6P�H�K�����J���y����[o�\h�tx��{;[�/�ҝwz��Gs׬�)�uQ�U�Gé)��v�'?�:���H�b�,�Z����S�F���^���Go^z6�V�;���u�ػ��m{Z��ܮ��\%�WT�� �h�������Uɞ���}���&;�؇�1v`����y��s���~�ZJ��"b/��E��{������?��k/���S�����s'�Py٠�K����ްn��9s���
¢��=�}�u�Y���W��6S����ִY��w��N���S!z��}�'�_R�j�j�뮻TI����_%��<B��VeU�=sNs��f�"��A'�[�s�f:����n�c�k� \bD��_����~7�Ҳ�O���3���_��K�jk�(ga�2�l���w_z�soK6����500���.`���^=DT7�ѥxz��C`����j��b�0?j�\��P#555QKk�j��5�x�L��O�"�N*�V��ݦ7U,��}a�����1 ���<n�{%%%R�)�{�߅�А�뿊��T?��/ozs�[�tww�͙7������_�B��p�`�=���X��������#�u:�� |x�h���;��{x�lD�>?�x㍴a�Fu�?�񏩲��jjj��Su���a$��Numt��Y� F��l��?�����t:w��(�{��M!���"�ćܶ-=����TtΦu}�}e��b����R~�*̂W�3����";f����uw�C�]OQ���~�ajb��3���o�a�:q����,%wXǇ�q�{���08`T��~;��ϐ�L�']��2 b/\4��z]$\5X`�`Ne��Mtt��;o���#�?�^��X��1ɕ�>������*�qq�>�yjj:��%������$=� QG;^����q�`x�ؐ�k#1�D��{���JKK%�/�{A��`�~ppp)n@��k��C�uB�ڛ���c��ǆV���¨YU�O%��#D�� �CV���a,���,]�T]Kx\���s�v�<R��[?�=!�y�py��	j5�x7<g&�z��02�-h�i���1��"�����%�z.�|�1�^Oj�U�?�)�B���&������q �A������)��A��?:M� \D�a�"j�d�_��i�[�@C���m ���;�!daGb�q;Sj�]'�A��v�C���z�Y����t8�CS���6 "���a�4�x�^)��˄�� Lhz�������"���@`�v���V=UNu���Ľ��!ji9�" ��ܲ�j�_��9.*/�P"��.�3�Q0 p�������1�{br�a���Tr0�H�e:].���}��qo���	�pY��	��`~&k�r�N��!s�,�t����KɄ����;�0��!{�ӣ�At ת��V%v:�����B��Q��G ���0:p~�K�S;}n�_TVU����t$m��V�����^/�{A�� ���ӳ��w1����b�����v[\���>������fW��{�;�Yw�r$桕.�z�ǆ{ٽ��O�Æcp}�_�٢�L���)���7A�������mY�jTȱ�b�^�/�đ����z�3�u/z��������H�{x�:R�kB��Gb�n��t�
ײ�p=8F�æ��ƨ�c������� LPXЧ����֯�m�P���7���W�����(hnnV��;�����ΞGx%yH΃���|y$���CotW<����1����3;H����� LPXL�R��,�
�:�!�@����:޷]n%u���{u,!=-�ډz
��S}����Z����tZ���E��!܏���uo|�w��s<�M�� W{A��tvv�X�7:�r��!ϫ��]ŵ{-��$9���dZ��,��F8�i0n��0��'���g��TQQC��J�ޏ�8�."��fЧ����TR������{�֏nhh�� W{A����>����,�N��'��w��x]v���
����qlGGG1��-�流�*Va�s��v�UT�qz{rB�������"	c��n_��?ǯ;�5I� \D�a��Bj.���YM�s8T(^7�A��Wg���d�ut1&���vd�,�Q�D�1��\���� ��8�QQɷ q=4�щ���Q��p0� �u�p���	F���{%o�c�q �{|��H����a�̠����:��r��WT��SL܃�#_y��|����i{ ��O�ؿU^^.n�*"b/��X,v�['���GV�b�v{U�b�K��}#��H��Q |�Y�0�i��u�]_QY��C��E{\�0pǲs��"�;��|60����Rr'W{A�`�����u>����HC�!޺�]�����=ްN�{��u|x�8������(e�Y���B��%�`Py&��yC?�v�D �[}>'�b��#A�*"��0�`q������o��s6���cG��å<z��F'�AرQޤ�����cϜ(�LQ*�Nz0ܔHإ{0jkk�����A�=Nu=����!69;1^=���@�O>��i���J]]� 	�pU��	�����"��A�\{�hd���A%ԺE�N��z=� ĝ���(��aNII)�>9U5U������H�f3��g�i؆�aŵ~P�M�!99�������'W{A�  ���w%�������=D�v��+z� �`C�^M�Kf�w��7X�G3=��H8��%�ej�M(T��^���������cug>d�Ó�A��	��@(��>��5� W{A� ����X\o�!��^M�c��������V'���G�$Sq����������S�<��z4.&��k��bY�}tb�n�S����`P��a b/ T������R	��=��G"�����M*�F�B�ʇW��w0T-�i)#A�a1��ReE5UUU�~�0�P�8 �D�ޣ������a�¯H�K� W{A�8���r��ZP!��XB��c�;�l&�^��y������v�/�#�abBh��q��w��U��y}o��c���·����(?���q��� L ��p��z�-�b�Fs����bR�m�b�^ͧ���c�٣��ԩS��G4 ����*����*��<�ao��#�o�Y��Hp9\
�(�f<���!��{6FI�q��� L X@XhW��촽m�
�#$�uxL��b���T���{[[�j����t�Q��g��zH��J�g��{;�O�����&>8�}�ٔ��5{~���r��#A�"��0�A>���Y,���c��r��l�=G�����u��9�^},W��N���?8���!�H����d9��N̳,�݋_'��������_�I�q��� �s����X�ob�-�_��Ղ���lѵ��L�������"">{��x�>*++UF@6�&#��C�d�Ϩ����@C��ɥǊ}������ml4�I�q��� �s�^��L&3�E��]��Ycv=�������z0N��:��S:��x,B�m�)�*�������u�iUS_W[C5���{�˳��?ٌ����Q����(�I�5��% ~�c�?��q�rI�q��� �c�)ohhh=��B䵨#��n�k�љ�Z�1��^{������ȠGV>J���qhy[^QF���ʻ�d;��l����fLr�P�,���|������H�q��� �cb�X9��gO٣��XZ$ۡ�^���	x���Y���ǱX��{;d�S�N�Cb��� ��\�^'��8]�χ��������1a\!b/�4�aQ�ϯ� +Og�c��yY��C��N��~x�z~��'��ɓE#�N�S�g�R ��jjjT�=�~���^���(��0�B�;���]��8"�la�!b/�'��Rަ�e��C������t�; ��A 1�#d�u�3g�(�^>�������A%�(������.a���=y�� �������lI޵�����Aw���8�������.e���Zx�r���uz^-����D����-Z��x�|�rjiiQF�C�B󕕕*���)�����ņ=�_{�|,z����$¸C�^�),��,�+��Ch�f�Mt�
4�ƀ���+<���{O��z���ު�=|��jx�zs8mo��8�\��'��w�C���>���g��ɝg��	�0.�����l6[��z�:��l�=�_0�W�=<����b��Qc��#�(O� ��^�;���uFq��^�G2 �^�>��������`Pz��8E�^�!gΜq;��U,�!��T:�7D�����:1O;��}}}�z�`�^�8=����1���5�X����(���Z8��'�!>� ��� �SD�aRWWW�7455�8�����׫�=q���^=���zz����t��Y�F�� �9���@�Qc��zH������z�G$ a~=�~L�>���s�K� �_D�a����###�ǎ�kllD����3��+��?�ʠ��}]R�0=>#��#YO���I~s|���p h��Q�٬�k��A?���׍����ii�޾`0�I� �[D�a��������X��^�&ؑ�>��B�;;;��>w�|%�o���=��z����{x�ix�ا�`�@7��_�||�F/8�!�n �{Ag�jkk��5aF��n��~�]��C�!�t������Z��~��� �(��q�JJ�Ƅ��O�|}�q��?����u/|~�<�s��; �la|#b/���<�lxxx1����{<��y/<qx�}x�x���:#a}9�@��N�J[�lQ��3�<��}ÆT]U���c�;�~�b��y���Y��\	6&�����$¸F�^�^��ױ`��I�F^g��>�C|�L��D��q�y�_��uO��K�����O.\�;vЂ��+Qk����|t�>�}=L���o�d �D�a1222��z���k쑶ɤ=7�9�� ���� �Ç�s𾣣���c������@�㣃����y��U-�Hȳg�ۆ����p�H$�k���\�|�1a�#b/�h4���>%�G�>J�p�Lv�=n��y�L�`0D����y��z>�;�m����Y�!�yJ�P�Sǖ�U�sϽ@˖-�o��꤇u�}���v�������<�:����� N�CEPq��(�#���YRR�E� �{D�a�������"Z�˲��s�D8;|�vy�w����#ń:�<<qx�H΃7�s���s�x�����w�}Wy��Saz��-��:}al�:���_X8���F:�0!��q ��ΌFc[���H$�0���Z=k�v��ϝ;�\.���X��j�ew�d�b�hqp���\��o�]�t	���<��n��Şɲп�F�Q������� ��,��~�<��H76q�z5D޷^��8�:�l�.&ёQ����p�ڽ���=o�ޣc��.�-ίg",�;�u�A����8�Ž�t](T�pc^7�v=�� �0�I����V�s�D��L��lB�H�C�u�:l��཮�Gh����~�V��4��W/{A�7��u�:]'��!�:�N{�y5D�~�DF�X�0�T;��C�a \@�!��h���U�s�a|��1��yݰ�_3|�}|}I��	��� �ؓ_�b[;<<h���cd!�z�-^��L�A�e��M�h�� ���v��\���q9���|�kc�^7����xD ��t�0~N7�	��ﬨ��� {A�������y��ի1����,N��{1ĺ��V%�%�v�^=��c��5x{�v�P� �8"�A��붍����!} ��?G3o1�A�0���U&��⻄�Z���]C��Y��Nw:v����N���#��M.���������ʋci3���ܚ)S��r�k��0"����Լ_fGF�����]l�!A&"��paAu���m��=�/��ա<z�C�!�zP�st��~;
`w�۷�Zs��mn�V�X�j�, p.2�a,�v@�ҫ�=���r;D�u����A���	��� \Eb��J��6���c���wo{�Z��n̝��iӦ)qF Y�k֬���V�d�<g���맫�?y�*��|>����>�<�]-�T���*�RCv`4 ��&�%���?�n��%A&"��p�������E��Z�=}���d����a��{�ֱi�%s�� ��ɓM���E�72��Ѳ�K��矷�,t�˫k�q�0"�< {\��ʇ,|�����" 96N�w�$C�^��L&��aY�Xojj��m�cO\7�A�B��t:C讇jwx��������l(��ʕ���/ӌ�j��o�U�s��lA��c=_w�Ch��{ C	|��?�F���0	�0�����iM*��1���F�P]r��g�u�c>��X�Z=������@7�$��^`���o��✥u�6��z���ud�WWW+Ͼ ����'"x�=��4y$�!9O���D�^�,��i�e����Z���,�x]J�Q.��� ��ɛ&�dhxh�֮Y��ollT��z�)�3g����;�A̵7�ͥ)����m��5.��u�N��/�r9�c�CB��0A��� �뻻�o`����j�ZG�<o����ti�;���Q߀{��ݫ��o���1c�>�D�����R���h@x^g���#j���羮PY�vU� ��d LXD��*���_âzC&���n�h�$��oϡO�أ��ݠ�-�n�ۥ�����y)�����t9%�H�[0�M����!���~6�iw��=<x�.�V!~�6$�mx�)����@8�b/��a#b/W��,�sA��'Nۨ�91�5k�����ىv�b����h\��͟?��ꦲ�ۣm�l���B��y ⸆�a�A4 Q]ۯ��@5��eS.�k_ h#A&,"��p�a��n�`x��Y	-z�g5�(���nw,��l�2�t�|�w(���4�Q�-�v�
קRqU����ӧOS��7ذL��8�����=�ǽ��}�>�M~�� {A��$��:�UH̃Ȟ<y�r�p���X����SCCC��=j�u�\|F9��l��^U��sb�(�㠖�sj��`$@�u�<B�^��fΜ�"v}�Ul�[H��9-g#�?*!|A�؈���y�px)��,�F,��Ǐ��uʫ/��E���1?88`���d��#���R�$���V_���f���s��)�>D`L؝��b��ԩSՆϸ�}���a������$F�^� �A�����[{�F��j��/�W���y��Nvvy�YY��;=��zx�؏D�\"N4P蚧�X�uh���P��Dt. S����������^&>"��pa��eA]���^ho�h<ƞ�=V6
*oay�
����(�C^=��,�r$�l&���UWU��=��N��C��`ƀ��g2���+���!|���i�0��3Hm� LD��
��<�i��ʶ�Z;��!�g�V��t(]��W�W)aƆP�^w_�d�j���t<$��[��S�����[�Y�À�����z�M��r��d��G����0	��+��GGGo��2x�U��w��:s�h2�V�����.%�n��c*a�?�%�h�e�������pR�P�уm �I��{��z�j�5o:�^q_�L�9��l�L�?�L��I��� \!�+�嗕,��"��;x�g=DY'���y�������I��y�:_L�õ���]]]4�az1L�����z%�?>�þ^N���Y���:���I�	��� \XD�H$r-*z���t^{�J��cg��9� C��l{��Z[g6�O�U{���f�!�Z������S�E�i����{-����a�`���A�����|oe��]��e�F�@���Y�_��E8^���8��^�������r ����������PZ���;=��وhv��>E� L
D��
�L&kX`��Z:�����-��u��!�(�+//Ueue�J%�V��
Ǣ*�/��R4�8o%�J������P@��2��M9g�m�R.˱�]����0�����D"���v�i����;�0cB�d<�zl�oo��T=���S�p��t��*Ͼ��\gΜQ��z��3�3錪�G_-Xv���V�׵��ޟ A&"��p�񰠮#���C� B���v����c�M0�W3�9JgϞU ̝�9s��ҽ!7�GF��vRww���Ӈ���z-�0ЬG������?�B�d'A&"��p�aq-c/�Z~�1���N�C=��N��'n)O^��C�[ZZ��W_c�=E��Si�����_��������ww�T�{3g�R������È�>}z�F?�ϑ�{x�l^?O�wte]�$¤B�^.3,�؋F�1v�p:L�OgǧSy
���D�T*C�HD��Me�4��#�᡾�Aj�-:x��֬YC[��H［�%!r��d"a����d�h �Mu�@.]x6t�ͩ�r8��nk;y��� L6D��2��gtttK&�)����� ��u�z�_o������6mM��I}�t���:::�y%�R��t����c�
��J�`M__{�����d�*����5����I|�5��!A&"��pa�ga�������@����y�=�u��I}��t�=�г�>KO>��Z{�'�PS�][_V�-����s��0vN=�m�A�ϖbc����"A&"��p�`Awna!]����s�{�n���ܘy������^J��t���]wݥ��}����=��U[[�"@'�\�R��z��nΣZ���q_�������d���D�^.~�e,�AݩN{�ڻ�r �v(�Th�q4z̭�9o�a@`-����׬R�q���U8���(1_�p�:fddXDV1�?v��;��~+	�0)���D,��⼊��	�Z���7=Rv�Z����C�!̨�8	{���j�Gƾ.�[�j�ʺ�>t�ӹX�]�q��e������Ʉ;A�����e �tXt�V?���Db���C����p>�u�XK�,�DGO��=��;�/��X�M�q�긇kh# Ƃ�絽x���	N~�^p�[�Z�d� L^D�����d2�Y@���NϠ/���)�N�^�^��Ko{�o\���0���BN ������GF?^qm��Y�o������'A&-"��pE�x���3�������y���|���>�Θw�쑴�t�!�,�(���&��L��.Ky��j�-r�k��v���?�n>}�A�����e���$9<<����8��W@���)��̏-�{?��+���[�������cjǾם�������Cp�_��4	�0i���C���Yh������5�����aD=]~���c��$����yfq��h�=v{�n����SA��u�v/|�8���[e�^&7"��p(��)l�����x<�Y����nĨ[����Bnh~�p�^�מ����1��t���s������5���Ǌ}���a�į��I��� \f���GX������l�������
d'D����x�B�<���!#?�B/��z;�/�>���U�>Gw��՟�{� A&="��p(x���؞J$���j������\.3�E��}���ѿ�x���C�}(T��{$��>��� ۡO�I�4����C� LzD��
ShIۊ����h45�����Tj	{��,�{ �UX�7� �N�����&9@��떸��m�Z�9���^RcmA����U��;�/GX�["��,�Y�o��+X���|�^�Gy�o���*�����Wo_����x��&$� �{A��Y����,��K&��D�l6s&���[y>o8Y���g�9�^?V���')���(��#�oYv��4e��$�{A'����}�X����_���U,��x�2�y������=w][�f��xSzS��w�Æ�0	���@�^�),�ht�Ƣ�944���6�N/f߄>��,ޡ�u�@���d>�hgL��q���!A>���8�EYw��G	�i~}edd���/g!���E�5��PƧ������+�/���'�n����"��0�($�!�mn����X,6��o`��Z�����Yd7��H�B�>�����7ī�"��0A)��c�� ���h4�{��xC��[��Sx� ���og����v� (D�aP�����"��_�L&k����G�>����q��"A>P���$���bc�o��b/���{�=�@`�A��!b/�~t��,l� |@�A�I��� � LrD�Aa�#b/� �{AA���� �$G�^A&9"�� �0��A�I��� � LrD�Aa�#b/� �{AA���� �$G�^A&9"�� �0��A�I��� � LrD�Aa��� :ⲍe�m�    IEND�B`�PK
     eO�Z9?B��  �  /   images/d18021d8-4522-4af4-a3c6-358ee97fa8ad.png�PNG

   IHDR   d   a    /�   	pHYs  �  ��+  �IDATx��}xT���;��$�I�!�@M:� �4�E?�>D�+("
*
"��HS)�JH�$!j�I�dz���}���|?3��}�<g�L��9��k�w����� ^��x�ex@���!^��x�ex@���!^��U���v��dRR��H�q�Lzt였7��Wo� )1�~���;�={�l�C��B�Z�����j�\.�Q��{Z��`)�r�bώ]����������G�ʒ���/P]u���0 X�3�����|� ���E�3.&���e�kBb���sK�w�	�3�����r��m��V;��\����DF������aE玉h��r��mC�4�F�Z̗]k��i7[���'E\�
���n����.�]�����KHOO��u�!�̌=={FTD(U��٭�]V���!""g/�@��=q��e�X��Q��Z��&�Q�X���)�7���$�1�L�|���eҀ���r���iZ����>������!cG�CFF/475�`�*�� rS{�'&�$3_����b�r���SxX�*�bl�u����3e���sxj�B�8���G"��RDF�]x���~/�+�����ov}3l�ƭ���s�>�"d۶�1m�TT�Ԁ����J>���p�����/^&�a�����&FDx����i-�4M4�ٟ~}�����ԙ3݄P2(�̙����X����`�)����ܢ�z�n����5�!�}��2���d��ox<��`�~�f����:�9��UӬn�{P����
��f,����~a�K�e0݄L�5�|���q_\�����M|�]R�B�pc{[�߾���mc�O��5�!aaa8�w�A��N��f����k�=B���K�nN�Je�m��;)ݒe�*U��sV��w� ++���W�`%� ����؏>:���8w���;��47�`N����O^�O��܌Ĥyks{_�g����fs�&$X.�С�즆����J'�5ӵ�h�ȸ��N�322n�������+0�ᑔ�����j�.��!���9v��j48]Di3OI$��r�l��u?�J-��E�U�¢B�͒�����D"�TS[5���q�[o����\�
y'N@��:��,�?	�9,&<	�"��p�T�8ď��F��������"�hm[[�;^MMK��d�����m"��PKs�cu��q���_����D�?	�X��T(�@����2�<�"�h
B�l6�E��p8�X�@`-))}��,����Z�J�5*��
{�;�[[# �F*�C(���_}�5 �Jb��[6����������k�)B�B��P[V=q��@���	b������P*�%�~�[�P�~�U���ş��p�Q�c9�F?�~�}���1_Y��V��������������1<55�W/=b����'�<v�>E�H(��h6�-��� e̍7�Z��q�		���p����Ψ��o	
{��,i`�r�N����W~�ƍRL�>Ç_,��ݧKC]����*��C�n�n�� �<v�>E�D*Þ=���{��[,���Ga�j�I�[z�ꕼ�v�Y��-�Wu��å2�R�t�V�k���Crrן�;xp?bbb@ޓp��ݥgG����ۧ1S��ݻ�WVV��z�}���h��.�ܛ����y�V��]���z�Ţ�z��͞8��gƅ��l�r���ͦ��!����:��x.$fNEH����`H"�	�6�����/(,X,�I�k�)B�N��u﯇^��#Q9�P���<G��
�E��^[���1�/ڜ��\6w��lF[��/��y��۷c��%8p��xΜ9���d22$��=b����g+UַmV[����g���FYi)M�PBD4""~��	0P��E�:u2�[��[���b����ׁ����lH$���;w�<������F_b���,6��Cb���Gm�[�O�0�m��}�N�!���j�1��1Iv����@ppJKo"H��B.eZ���N���mokAQ�_~����Aѷo_�[�>�����r:aqX����c���$@�^�f�}ᢅ�N� ��$"""@u��=��7�}��Fǎ!���??�º��g;%&�Assz�鋏6m�����*;�0֬y'`�'����,b�3����A���R��3y<rsOz�Z}��g���g�}/��2}����|U�Af�Q��##"�m6�0.����;�H��p�;�k��{�娩�b�YC8�\�Lf��Ƒ�N��syܸ񅇳��~�V� D�����kx���r���!�"����6���*G�Ѫ+�*0g�ll����$�ζ�}�m�~�n]�=�$���8m�t��	1W|����u뭋_^��k�zB���� �3zQ?0�d4�S��ħԃ�
$&$V��eb	�[>��w�ۼi3����ʒ�!;w��d0IP`v��nݺ�ࠝ:wW@�*��;�����S�zB֭� Ç�)�@�1�[�\�z����H�cgU:z���5�q�ֵ?o�����FS�#H��`��5���L���ù6|��Ϝ9�.]:Ó�jB�xb
���P�/���/--C����M�<�F�QL�s��i�m$��=dee��B>^}m91O)�h��b���b"%5ŝ����6�����/{����k	5r,���V��ǟ�������	��6��$G��H�!>_�7�јN����s�O�:��'&�B�����whi�)���r�:����JBF���
���:52*�s��¹y�&�-fp�<���V*��h��6O���PQY]]MLMǃG	���y�qy��L���!��Ξ9��$���2v�c?�q���v�Ԩ蘭D�|jkk�X������q�III����\��
��N���tz������ʪ*\(�ǐ!��~k����o�_"���U����"�����gP�<>**�s����bb $���!��rҧ�J���555�a��ȑlXL�7��V��L������kո]Y~����$>�,�3�^C����q��5�&��bcc����s�B!tZ��K@��l��]���"3e��h�_�x1�j���^��Ν{q��!l��	:u�<�f��~uHH ��g0t�f�[^^q���Bw*�~�k�<y
�	 ~�߽{�����[�.II�&���qTTT���sMD�mw�I\.7�|������9���E(--ŨQ�;\�v����A�똘ZS���^��ֳ�?�6k������}�7HL�DfI��
�"�DT�ёQ�6T�*��2���^��e�$���r��t�Č	�"�^�Gxx�o������Hk��!�QI3ƴF��hi�����7J�k��/x!�21h��l������v�(jF\l,n�A����*H��$,}������
2�4Ԥ� @J}K6���o�9����ضm�s����[�j!�6��E�MS2=D��Ǹ_�
B�eg�V�ҐaD����*��i#5��'P������
*�k��%/j���XrC�4�jn��:RN�>���bĈG�IT��B�D$$t�A Õ�u�p��)�����	� $6.y��!66f0hJ����AgD{{;"��Qt���-Ӡ�+�R�.aVFG�Ҵ	�B�2��\*���?�t��C�Kf�nss�t��`Ђ���y��7K0g�,�Ox!����T�K�-j���;w�@ ��l.���ۚ�[��Cn���W��>�H�'$�m�5��;��!�Ν�[o���{�ԩS�PSE˵QQ��h�f��GD��������իp?��Ь-5K�<<��t9��k 	hM���P���Y��`��n���m=a\�c��Dҿ'U�p7�C�/Ʀd����ҥK�I8ݕ�\h�Gf%`�=q�eʔ�����;!M֯�ȭz��M�����
W��a��t`Ҥ�g�y���q�:H�u���|�&�QE�;w�/Ɵ2e*�͛KZ�I��p�]���3��?�B�H��+������ע��6F>2����;�I��EjJ2��ݦ���|h�5q��ȓ���I��!��K',����:M^ޑ_���	|��Z���B1�##��۝�r05W$l����8�B�N,�Iހ�J����' �/J�S_�ڣ��&.x�e��(��"7�*�Iy7o��&b͡Ѵ_'�njl��ODd[{�ƚښ�#����[6���_~���9"++�Q��`Jw�/!�3O�>�]��Y��L�7��ko���k���p����pZ�)Q��xxh�)::�ʪ۳��8]#1OS��M����O�^����u���?��!���Ν����8��'���+���@P�ND��A�A8}ʳ����ښJ���M��ň��6H�0�Ӷ�6��tO���7�N;K������8���tM��xs�;����E�z�m���\�Z�
���سg��4h�����H�!��$��|eeR�S����QB�Mټh)��$]��[�FL���N�)��vΜ<	U����oj�QR)NK��)Q��O�:���������xxe��YڊY�f��\���
6ף�U=�h4�0L�	����X̴J��С,� --��rd�h,�댜��ֈ�=ݧM�4�l����3HO�'�qr?�z�̤a��V]]�.�"�N+�O:N��=%㷐����Ǐ7��\])�P(!��O���A^�)x<F��Hh���?�%@5��um���a�XwJ]��>8s�,��\�O�(T���B�_:�v�SgʆJ��Af��#G~�\k׾�}����S��=6��`���0���!�Vь�
v�����xq�s�x���I����M����0�/��D=͚V�f�'v�Fg��h-�����6��3U��u�Ug��	0!7|�ÿ�7�ǎd�p���P���.l�*$�բa/	�_��Z�_n�x��#�8Z��]��H�I���_���rd�!
0���(�hh��ǵ2��^9uZ�&aW�JE���?r��H� ��:�.Y��C�a��n-����6G��R��.�7	o�G�=v%�;��R���P���5UqQ �,l.;�Iȹ|h��		���_˶0��w�v�ʕ(,,��I��rs���2����z�&�Bμ�f��+�Ā��m��	i=����������ዬ}�Z�qe%��
h����E~��w�aPt��x��[[��|�n���w�Gq8\�'�ݦw���!{���O�g�����m��	�"a�S���k�N���6.��W�! �Z�`�a�P�t"�ھ�s9���#�n�ٿ�]�����_{�y�ݒ'H$R�w�(�w��t%n�����)�q��wEX)!g��/�
q�eh�e���D\�����h��䂗y�
)b�L" #��b��\cYBG�����x��?}���{�+nc��Y]

�z�����I��.!đw���I��3����R�� �:�Ln]�d{b$��p
�и��NLW|U��G;O�=��a�ޤ4�w-[�={����XxX����݊J̕��v��tEi�-x+�2B
^y��霼���讯��Ҁ���VTZ-H��C�䉈��0���l������l���W��|�#eӦMx�Ŝ�'�	
B������w�A��٤P��ۮݺ�-���BC����V)cq,Z2]~�| R����D���f+T\��
V	��+j���.���{ ��-���_m݆��,��0��$�IlU��-9��j��'��kxb�̜9ފ���s��x�(��K�s��Ke�&��p���O%��X݈l��r=��a�j�jU�����:������ڶm��ك��F_)F�*hBpp0����]Js'	Ỻt��˗�͸焸���12i\?ȫ*�,���\���as8"�Ƅ�kj��aCTp�ւDy�i�:m/�kEƌC_<Hu���#t�4]�OM�\.�:����cr�3�c��w7�<�{Nȷ_FtZo�	RG�Y�3��Bf��<y>��"�P94�D4���ok�oAn�"�� ��Y��5r2#�N����ҥ�>�<�h�"]$�^��p:3�\�����@��7��J�ú�D<��
[ޙ�Epؒ� �߼��.Ȃ��ED���=}�|c�ڳ����^������s��Ԡ�����Uj4�Ç?]FLR1��jܦ*,<��l����D���?o
���I{�-����a��� �S����|��T�G��OA=�77�@k���f��}�\���$�KQ�cȷ�t�ass�{��2t��К��J�\t������۾�-�)!F��`�ۂ�3���n�2�(׫a���id�(`(�ui9\C��W�UՌڿ�����Q�<t�eB�)TWWO�~b�ȑ���ށ�DWMMM���$$t���_�RDB�
x9�)!��=�I�3mρ��K��jW�����Sш�S`7�pk�68O�-/�]n��ٳ����]��>�o�N
���:�%�ϗ�"��@��j)J^\\��4�wg�帧��'w��k�E߽{�8tT��j���ij^5wt���-=K��dm��M�J�ywA�YQ�En����lIh�����]^@�҄"5kV��e�X
��T��{J�O\�Q�;�-��]���&��8��l���C�+��s�g��>r4"-4�~w��6*IH+�5�̧���FP����&EFL�����͔fx	qe,6���!�v�%�0|�D����?�aovL���S'��'��'B*i��B}�{k1�0��i����`2;�h=����϶����y����lGɡ3�juc���o�%ir��� �1�0�5D�m���O��_oH�� 3g���ˏ;2��t�@���.�DB^��^e�^f@�J�,�X�K���칽���HŰǊ7��������j����w_��]�nu>��q�1�/�ŋ�Jt�С� 00r��V�)7�it�#�	��vx�(:����t#KwO/�d���EL������HI�A�\�a0�T��Mz8.�ޟO͹�����z��Pw�V�S��BTW�����Gl|$	�t]������"���Q��9Bh_�"�j<or?d8Dwg@Zj/(2�'�.�u�
D_�OB3�4  �S�^�w�UB�uA�y2#��|��.�����ʝ
��[��m�)B.]��.�Bz�������������QQK�tS��jʢ��t�/�g����ĺu됚��x]]-f̘�^Cͦ���fter�٥�X�,�X4�z�/�g!n�mz>��>�ro���Vr���q͹T*�+�v��w�%�!:��m~�:�p9)cc�&��nXI7��A{���o7��D�{�#&�%|��=�f#�O��8�j��C��z�&�5q
8�}y� t:�'��*�^�s��'�a.��FAAA��}��*�W��ӝ}Hlq;u�M��aߩյѭ�����>AM�Ӛ�	#�L�,9%�]��qY���bh�`40\�l�m�J幏����	B���d4�tKIq��!�aе�p7�m��|8F��$!��zBh�DkZ�&�Ӌ~���>t�%%Ĝ�?I ���ӹ��`�d5C�����P?@��q,	s�t��ś#��^�wD�p���r���c�9�Ey��9�%��
Z�#>�49�@�F|��~X�|L(���D4�-:�D�.L�*������9��j����l6k��nK2�n�l�^&�᮵�2��*�=�l���h4� ������i�3�v�D
�b�I�o�Z�ex=!�3B(���.%����B�X.�Y.�+���W?�֗������Rm�S/�=t�:>Eȿ�v��'�g	�O�������$9    IEND�B`�PK
     eO�Z���*6 *6 /   images/a1588c66-a70c-44df-b30c-55fdbd854069.png�PNG

   IHDR  M  �   [���   	pHYs  �  ��+  ��IDATx��i���u�w����ֻ��mf��=�YD9�IKeI�l���Dސ/�cdB�I��$D�,�4����}n���pzz����}�yοn���&�83�7,�۷�ޭ���Sgy�K��(��(�DE��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)��(���M��(��(�@E��(��(�)PѤ(��(�r
T4)�됶m-�rr�W_�sĿ׎����s��D��Vn5��Ͳ��EQ�M���7�/�����W7� 
�N��2�.-�	�n�g}����tY�8�n��ڛ����&i>(�6�\�s�N�n�nӒ�{r꺶��;l�j���m��~S�V[���%�M'Ek/,'�n$��mf�$�y�P�;�;�U@��R�����*�S��]-�vՈ������1EQ^�hR���� ��q�f���R@�y,|���֡˥޸�n�P�n�ϒ�ǲa@Ԝ�j�j-�S��׎�4yUU�n�uP�,����~Ȣ&��x,v�D���&���ݲ�Zf9M��Ro�A�nO�q������)p,r�?ê*j�\6�ZN��N[66+��IK�'�*+���Òl�t�p\*}�)l��Y�-Y-��vIv��Z����u��gY��عeQ�_S�rRr���q>�ȟG�n��%Q���x����EQ~�QѤ(? )F.�QD�)�b�i�̓��`��Y�ͨ��aNְm���i�ږ6m���u�cLuy[r���)Y5%�O��zȨ�
�ꂪ�U�������[+�9m��a��R�_��P�KvP�"k�x��izDA���(�*9>yA@ESQ]��[��k��u_ٴV�zVZ�]�蚧5��;���)k����n���6����9?k�����W��vl�����q\�v��v�̥6�mg�z֡��ǁG�=������n��ޘ/���(��(�DT��RE�AE��|4G,���"����l�ͳ�uK��}g�Ԟc�q���������Ϣȵ�iX`���b�a��ˢ���?F�'�w�Z,�M,\��ڪee�PYZ��q::Dv�B�O+��
G���D�G��ōGgΝ'�&t��=�����x�"uz}�Y��I	1�A�̢�1���-���#�N�L:���vl�"jW		699��*�Y�V�UU|�1ǂ�\|�QV��<�/+Un��Ǫ��,#Ǌ!�����3<�(��;/y�w?����N�������VB��(��hR�T|_J͙�8ʲlT�VY՗X\�9N�ԭ�x�Z�-�}׵��u{u�xeUY"xPxd�dȲ�y�)��F-� ��-�u�,2�D~$2��,K�x[���k%5�IL!?���4�[
Yx8o�-Y3񾠼��Tp���yA��M�bFw�ܤx���pDA���.eɂ�F=�+;��*�,/E̐�S�ʬ����UC�|I�2��dB�2��c�"���uZ#�Z���ß����?����+��l���Ǣ�*��z�ucUM���nQ%�{�,⼶�`���g������զQ/���u��6��������5_��+��}k������`�$����Qk픢(�*��74,���)���<{p��T�����ES=J~���G���h[+j�l��<+ X��Vc�Y����q�ФˈD"AT@�,� � �����(��+���*M)��%"=��c Xl��f1�9�qL�k��԰�i�U��Ssi�$r��/h��K*o������JRjx�|>��ҷ*�m��J���Y�5Hӱh˫�IN�(��<r�2��$@��3g��%���sj���ҤQl*D�,�7��q����m�xo��ӊϟŕ#"Z�e��mce[[M�vi^v����>xG6?*��;�|�&g�Qܱ����������{�ng�tn߽{�~����Tk�E�a��IyC�H�d2��v��X��Ǔg��y�n��,t�������~U�~Z�.+��l�b�8B�ʦZ��-�O��TF� �e���JDP��R�%sI*�J�CŚ�fqP�QKd��E�>u����M.�.����}��R��[���F,�n'5�+v����z����sE4��H����!D�\�Z�N�m4�9�Â�����V�oס�g����mZ��ΩiE4��I#B8�|J��󊌷YJ�?�X��(ϰ�y^��*��kӔ�\�$3��@�i=������З4`�׬���F�3
���:���5�ٴ�O�o`���c1wӏ�ݵѷ�]?x>\w����,�*RE�K��Iyݲ*����Eq!����ٻ��]W�y�n��8��؎c[Mc��cy�/E�I��t�F�x>�J���߳ȁ�ZEr�b��J�&�f�E�ϑz%&�"˖��Bı]�.�V�XD��>�w�sX�����1��5�_��,r��,F���W��wD?E�8F����(*˜
q�`a�ؿ�I�?���ő�)�F�X-P�}����㴤��sZ*2�C4������,�}�o��4�H�����]~L#���w�'r�2��)-,ʊ��4��(d{K)�SC��s Jے�ɔ�-�)���ѳ�e��x��E�e�Ֆ�HR$�ڟ�ٝ��w^�{?�wo�d��;���ϝۺv�K��z�.]���抢�BE��b%���b��r�>]��墪�V���-׹�yްnk��N7�����ےR��#�e�p��e{R���P�Ȏ�(U�s�|�֬�H!��\�>"G�FA0!EwR,a#Q*~.���J���V�w"�+'�l��j$�TI6���K��lV��b붑�@���#���" &z�T�vE+�Fz|���C�9�_+�����O!�[��D�$5h�t""N�T��7)�.����3O^,W%BMT�".��r�@y��λ@�	������2�x���H=N*ʌ�;�����O.����9��P-��򪴜 ������ʝOg�׾�¦���n���O>qeq����a׿vv}����������_������v��P��� T4)�P�4���yV��)�w�"��?E��E�I��鸑��M.���(��h�g�m[�%!���.�DY%b i'+[J���qY8��#m�h�w��ǘ(�I-�Xl�f�G�6�Ǣo�f[H�!���B��c1�&�>�CD�N�{��:��^u�5+�os��W-��_8nD�X�ER��3�	��&bK�X��kBtL����NRyHIB�5&�'uX���)�����k
j
X0�h�����t�{�����
`I�HJΣ�|�z1��x��-\��s.�û��|PUԾ�2D��2��%+��e��k
;>�_���KeA��cv�ֽ�R��z�,+�,)�y��I��r��YV~�o�?�V/������^����>ya�uP������I��d����r��K��Gi�S,D>hY�e.}Ǳ���l���o㼜�b��]B�ͱm4ҭ&)iDjԔ�,,�"�[����ػI���C#E��*b�HQ8���0"Ƣ ������D� 
��+#B��՜)�^5š�Bԉh�Ԋ�����W������{�uS����4Vdߑ�E�K',�Ƴ%-�s�v":��A�4")7��H�����s����I)ġ�{!j�����
B�aI�P΂g�bu�b�m�B�*]�]%��L�4�$Uhzc�[l���>�UdB�n�h�hE��6pl���gʼ�b�P"���Ţa�� ������|�=~�QӼ��GA�.���ݣ�/��꽻u���~?p��c��������|���B��(ߏ�&�G
^(�������k� /��i�Ǭ���e��'��֪���l��>�>���}��^(�"i�G�)�n$�$�ܼ�bA=�#�߈ ���u��Kҭ�J�5�[�t���!�5��pO���b-�Hy�>�xa߭I���(,�
��VoD���W�$2���iQS[��;L��H��a��|�,NTBT�G	WB��nܸA��ܧ~/��'�}�E��@Iv�5�1��IR��I�Y+�ym,�Z0��2�6�y��.��V���d�2.�*R�hm0���VjMMJe���+�X�L���3�7�"�K���J�ҩUژh��\3��
�,��<l�_�@D'bn�k�t�BH���,T-*{񨂸J�L�T��-����}����֓/������矿�����/�?��?��+߽���+W�Z��(��&寜�|�./�&�u^7&+�g��:�j��r}4$?D�B�i(A��x��E0���s��M&����C < J
^�%Hâ&˒Uq�$"AuIIZ��\�D�����H����|R��{q���Đ��pJE0�X,��z�.�||!�Br$�V.�K��X��\ݜ:l�)'���2�$�&��*���U�,Q��?�J��lF�GGd7k,
��c P,{7S<�X�H��/�!L�n8���U��1�&Q+����в�(m<ڛ��_z���ۣg��g>�Az��:����,.;�J���li?��CZ�l�8�ԗ�q�qBY��*�2~,�����Y�͗�Ԋ�,��6�:I��"��l곐�X�E�����XJ fc lZ�j�p4�f��}��Oz��w��ݽ��+������S��ξ��#�1)��EE��W�a����������g�ے��u�b1M�bx[`I���L�F��a����"
�#=d�G��]|/�oي��x�PoV�����@F�tX�ث�q�DH�ȖH�I��=H�I h�`Z�����߲"OiooOćw�n�XԦ�	(�#JS���Yuǯ�P�ݜ�wkҍf�Je
�[��_�X<�KD��݈�o�����uBH�Q�dZ)5�$[�]Cȴ"����2BOA�DD�1uZM���Z�|=����2a;���{�51Q�B�D�Te�PV
)M�^�A�ʍ������J�T�"���`��,��_��T�X�Q4�����m�p
���m�zþ /�O�_�V�u{#\?���?�N�v��;{��}����3۟�_~��}~�7�}����+ʛM�Cp���Z������GM���(֋��$���|�x��ql��Hʋ�"E��*\�����r�ˋj.�R�$�a��������I���yfK����j�I��������?��j�W��d�z*l �>��ٴꛨRS�"z�1%���U2ϓ޸�]��1i:�W�7�"i�JE��[�(�t�EgF��:�6��E��
|�b��*��'٫9S����n�_'5��R�$={��x\I(O��~Ki,�5:��cQZ�k2g��`��{"�N�ݑ�D#��E��Z)��C���/U��O�+��8���T��#�����f���f��l���{%�4^P�`��P�ﲈ
�cq��X��R;���M���R���Ʉ�n��βt�ʍ{�q�޳/���G_�������ҿz≧���'�c�S�7*���
��RzWQ���W�O�Yq��l�Dj��\	'"���<G���$�j��Ѻ:q�n�τ��!a!ue�h�Gg�')&�M�HT"+�v+h���a�� ���_��W2C�������/wY��:9������a9��8+����MIa����N����X&��T�DX�M&���u2,wu��)l�ds��)��B�G��DKb�ލ�8����ܠ�\�ȡ+ή$݆a^���Ĺ����ϑ������V��r|���洱֣�Q�z,�l���_ϖE<��6��B�Ƕ�6r��j�:���HP��$�)�y~em�xwv�i��]ڿx���ܳ���s4����1
X$&��Zf)�YPMSQ,��,��	�|��7D���`0����Ή���ߧ��]�O��z��t?����?~�����c���׮]k�?�U��(oxT4)����ޝ?�U���u���j�i$Ǔ�KI�dF4���Q��N6�$6����$��K��J��?a����9�.8K��d:�5�W��`������]�j3^��+iUk���8��q��g��D��˕�)���O�ӡ��_u�5��j�}���v!��^Ti%�Z#��?�1�k�{�4"ca`�X\��VE�(����9ƶ�Q-�c:�Pp7r�`�@p_0�*K���٦���f��2��kE��E
f����೐c�X�#~`=��:_�)��6�t.�
_+�-�?�Ңؿ�V�J�}j�-CP�G�����n2_P{�6m�Y�A??���)
`���N�V�F|��$�N�\����ir��������c�=F[[[���h:Ӕ�S��ɲ|�/��+w��~�������y��z��)��FE��P�E۽?+~n�f��E�[y�t����tf�a�Ð:aW�;�'B tY���S�	B�nۮ�x�+6D�I�6�J���(W��JCd&/Z)̞������t�!�VJ�Tkăc�ͱ�W9��:��HO-r��Ԧ�B�EEe��$�E�4>K'h��i,uB��%����JA,A���7D����o։��)���B��o�q��)זk��x�Y�+Q5��n�,��R&������,�#@=..�;D���"ڄ�,H�)�ײ����^��VE���״�Brc9`��Z�k�� �t6"hZԪ��my;�M:<�Q�ۣ��?���:�ﯦ5VEB: �~dal�زX�v�����ԺeKqPOҒ�gsZf�ɂ׌��+��h�N�Νc�AI����c����o}���C7��}�����������3g�%)��DE��P��i����M��q^v��2"�mr��An7�N'�0p�x��"��Ը@4��&�}i�����KNĒ)Ҧ�H2&����͏�Q�5B�#<<���(_y'����b����Z)�F�K�#�������&1����8�,��n�B���;MF���}҉g��QlnF�H��� ���d�"3�k�m��ý,.<2F��rM1�O%� �ء�ώ6h^4���5uMR���NU�GR��Bxd1~Px����(e81\���1��,�
�w�<��I�5�Zm))Q��I��cg�+����E�t��:t��UX��IAQg��ٞMs4����)����%��HG"�s����)%�8�!e�פ���ĎYH/$���Ⴗ�\�Ģ���P�\D�a�.\�`���s'��ٗ^��7�ˏ?��;�����o?s��G����PѤ<r�׋�|��j_�RV����@Z�=�Dl^��ܤ�l��M;>�~�|�^ENj�8��&AG��M)��[b;�*s2n�0���Q�?�^w$.ܰ3�L���G����q�.E8�V|�DIQ�IJ��Vs�LwY��~ו�D�e!��~��p`��ʘo��ZꢈR>�ZF���ɔ��)\��[v���	|��6u�U)z+���7���Pp5߾y@GiM�����[B,y�1�2o�����{���h��K-T��"b��๘����Q��(-��,|:=���J����4���~
��e�S���Լ-?q�G
qԔf.���|��D� ~�����B�_o�̲���Z��Z�C�M�Pٞ���{l��1Z@�y]�>b1�йs��<O3Z��Z�}�<\���ll���>�G�ӷ�ӟ�GY������?y�ɭ)��BE��P����U��c�i�.�����Ն
�!�x��X(Q N�A���8]d����~$���0VOf��*�$�>�>�'VG��eCE#K�&�a�&�jH��qTi)�x�u"�PH�ȑ�X��X�t�/ܞ�3aΝ�r$�<g�]K�)��J#_%��D�@Ә��N8�1t8��`���E���#+k91�si�&��.	��������)p[��q��JRfR�Q��	��q����=��2���hɪ,���:�`��o�`򈞸�E�y�2 \YHG=kbuX���	�}c8��8Zߤ��ޥ�Œ��t]�H3�a��KM��@�ִ��ǂ���Ad����Te	��-�W;��@�w��\�\ҁ�.��|�Z�Y�9|̑�ɹ�2h��t����$��&�����^D˄����{�o~�&�	���鱋�i�X�1����&�1�Fk4���#���&ݺuә�Ɨ��g���G��k_m�O��B�KQ�7
*���B@���9Q�����%Up��Eʅ�d�H��7�lKt&p%�m��5I7���y(ڮJ�\��ߠ�
⩱V)9�A��96����beܶM�Xk�1w�WWKj�L��F�5"� Z�)Lw����a$����i��+Gk+E���6x�!&o�e��yvH�I̤������b��G����ʌR��X}��� ]�
��wali�U2'�Eh`�n<�`�9"R�-KKā���sJ��9�%~j�,u�ŔHCy`��C	�qV��VS�H�G!;R�,.S�'����N���;�i^�,�BjY�5��3�[��߆�C?��z���:H�j�Xf�AX�XlOX�N2�g�S��"��X4�>�zCt.��{5�!�*����iY��4�!�Y@���)X(0u��v��oݤG����B~��1��>��ٔ���T�s�!Z�Е�\��l;}���^z����_���}�կ��y��U8)�M�C��식N���e���O8a�O(�\6�IY���I�D(���㣉��ц�k R,�$]�67�8����d{�V��ޚ4�D\�Z
�1�Æ%���"�����0[�þg�(Q&�2��	��&��R�p�����V���I��Y���-<椛�Z	={eU�s'F�(>N�yv$��G6�;�F��Ll��5�g�ᕹtˡUNR��I�aL/J�a���~9���Œ��H�/b��^@���uNn���$������s�aښ�.�̒EU�y��o�Geˌ�|��Jg�C%5K��c[�#�^c1�b�*!��Cj���C�G4����Z*�ݻ�G;�5�v^O��X�e�����B����!9,*C4 w�	וN<$TS��mB�J}� ��hH�?���R���E*#\ tע�O7i�ץ���'{�',�豋�h��r���w���K��G?�s���`Q�7*����I9����w��%>��.9�@�=-��
�J�>р�	0Hy٭��������DCp�h�W�&�h�[��vR�M� Ja���"�P���P�->HU#�a=�e:f^\��R")8��vc�su��4^�Q[��Wk\˥�]~2�Ε�����ӓc�*�϶M^��R�a���T��@� Z�1O�B1:�Z� d�r�F�")�B�lpLe[�bo����?��k0��<�p�X\�b�Qds��"B%��Ř5
����̫[*Ft&eq[�u/��"Q��-o�-m�$V_7Ȝ���P��ū!cQ������Ļ�%o�U��}��©	z�̐� dA�KJNC#~.ml����v~L9�b>�"��z&R���)(1�O�$�(<O�1ᩫO�tm@k���&����Z���7�QH��E:����pB�]~Y*�]y���s���_��~����2� EQ^��hR^s��|4^�����I1�E��Ȫ����2�)�\k� 2S�1�I��.��g��Ɛ��׬U*-�DZlS��"D�3��Dkj�"
�>�������*����b�|����%͇���0+1>�xe�(�օI?�U��8�u|jx����xO�I�8���E!ͅN�͍y~(i57������$����*2M!_S���
����>��Z�9�<+gt;b\/�3, 
3�,1��'Dbp-�_��K=���I���������8��m�
V 9k%��-�?�F�_��!T���;�q��J���X�Z�'ʤ�G��1�]�͂���ߔ�5+RJP�����bBz�EVEM�҅3t��E�6�d�(���͗	��xD����8�2y�O�У͵!�>��k��K�[ͯi�����>���Ǉ4[,i|�K��1mllXg7�Dd��ws?���^�o�{��R�u��&����2Y,a�#F�X�jV��<VK�D��� *���ot-�ENߌ�#/rY&�`��[[��m�'�B�3�hB�Q\�V�i$x*�f���$�ī����z��d`�Iљ�I4�]_!Ѡ�.Ă-�N�c��MD�<��5#^PkWl)To��i�7�	�O8��d'��j��8f�Yf;X;ާ(�k�y���hNS���y�13�jn
�!Q腔��.�b�A\��r� ^�߇RX-�ْ2d8G�2�J��U��D@D%�<��6:4l�6sX�ՔI���s�C�ۣ����\�iY3�J���m��,`�n-3�0�i\��x? =ɯ-҄.�Ǐ��tt<!��)dQ6��t���}��>:^�����ծ�u'�R>8l'�/i6��Zǣ��e�혱5��#jW�x|L6��n4��ut)I2*���^D�0
�����^}�s7o���˗/g�(��M�C����h!$\I���|F���_Z�Q�CF��&	!,��xjk���\��LK|+f��8�cJZ�A<�]�fU�BIm�+
�tq�P����y�=Vk���Q$]����_��_�3O̔���.jnx�'��f���5�`<��j1w�<��zI#:���d��(D=��wRծ"@����wz� ��E�i��P��#;v��DA8���H��UW�笺�m��M����/�b�]����/�'©X�������c�,�|�n=�xImp;G����$;N ]���,��\D�+����!�n�pN��1�ID
�5��\�v���z��{��ƥ��hg"nas���t:����#xM��E��ɢ%ߋX�w)�� ��ʽ*�X�ш�R}>��x<>���	�|�||�4-8�ta�5�.�=��H�����~�4t�bJ:�0�6���_x�����?�C���nQѤ<,�(�C-	����0��݌G�P�G�WV&�#�^�2���ˑq��k�tٝ�)���-3�P܍�%���Uj,�1]�j~0��r����f��ڡ:/Y��"~:~G"
��{w�TRtn�%yA��6/Ɲ@����+�NƂ�[���bQ��J�"b�ω�0a���\n���"q,G�Nj�E�8�P�R�O�4�񢝦tn{���F�h��B�������I�'+��-����Y1y�6�QM��k��?m���%+��`|iWUi�|�����I��ϖ�|M�Y��Y�v���XdE,Y���m�ő���k��I���:n�{ve�ʪ�Y8!$��u�����Y���+m�b���$��X��y7�C�T�7��Pp)���f�E�w$��$��㲐l<�{���gc�1���5D��YVI]Z_?G�ݻ4�="�/b�ב�g7t�,CXb�?�/�l��Aߣ(�I��I��\�_����ڵkןy��S�(�ST4)�c�W����h�F�Z�ő�ʤ��jK��DmD �	���6R�T/��Њ�Te��-_S�,8<c=��i��K�)�֋ �݈h��j|�Wjq�F�9��,xPP�dRb+�U�xġ
��nC����C � xPǅ����I�U�VG,p��L�ǒbq m�D���v#���i��m"d9�PS~���ڻw��ަ3�V/��lm�<~���s�}�T���*�7������a������$]i�r����4�]/��oiӸM];��˓|����2�Fu�w�"���Ӫ��_�u�r�.+�^`�����OvP[u�Gn�^X��WE_V�k|o�SO)p�_mV���L���+#S�v�}��O5˙y��)���m_�LO?��wi��t8���Ϩ?P��2��cu�(Ƅf�E��#)�j�,�r7I��7�f����Ey]��Iy(�v�p�2�@��˂"�S�� E#�D�M�&�� �� �dy�0�R�˺���KR��A-���^��h,���m��y���)�t%��HP�R�Ŗ��*,���s�B��<�4�%R��t/����(�E�f
#K�>uB_
�Qo��D�˸���*ia�q���buG"li���;<�CT���c�4�ڔd���)�K���hsm$c=�_�N�����6O߽w�?���/=��������O�;�?|-^W��1��EY�b-cbn�y�������|=��,�<�:iY��t���.��A��ϲ(y+Y����aA=�Z�ϯ�S�0dD*�Uw%j�|��,�IA�/\ �ь��H(���*�|9�����g6i��ѮM[gh��Β%MgtoL�NA��y���@�`@��1|���5겈������?I*��u��&�P��܂�4>���J|�l	�@(�?ԅ�42�f.YǗQ&.F��_�I�eYJ��LDOo0��Wi.uR��BA.L~�h5���
{+�A�N�z,BJ�1�ląF�^L�<�1�������
7aB��+����
�xH�Q+F�R��_�*
D8(�^���QǄ"n��%�ɩH��P���f�
jxlߕ�b6-�|%p<ˬ���}
��66��ɧ����ݿw���w�"Ͷ���{����}��.���7w��'.�����E��2�|�~��Q{b�η�Ydmܺ���|�1Y�kղ����ۊ2�)���*���f�Y�+t��0T��������|��YL�U��jX��lK�ѐj��6nX��!���HY �z��T���is}C�o����$�Y|�k�/�cmϒ���]��M�)��M�C�u�$/�S��9GRTQ�f�u�����U����G���՛Lqt�唲�p;�&���=_��m�9H��bD��&�Z��BQq��i5��p���UWi���!z!���M1�́�;�ҝ�4�Ni��'&�[����Ɔ�bq��BWiwU�$�h��ד��մ<k�lޢ^+��1&K^�m���y��M��J���M�Z��F��}��h����[7�x9�l˺x���_���O������3����G�:e�Z��J@ri��ڵ�az�����{�{W��z�_��q�\���	~������� ���ݚ��f�<�d0��>���:�Y��@�6H������
��-:<:���]�?<��l!��F�����
:~ӉgŇo�f[��&Ey]��Iy(�m���|�l� P�#g,B?d���@As%]a�bA�����-�V3��A�J�1�����;\#���H
������\�+����,@J-.yn��NW��,~*��XF,t���z���O(z���"�)Is^ �t4K�0�D�-�8=�GF�`���P�Dƥ&���l1��j�`���y�B]UR�b2��A�[bItx�Bi���t��K��t��y�/hkc�.=�V�F��s��Ŝ�c�`<����_?�{x�ċ/��?�|�ҝ7�K�3�X���6��=;_�����8�L.����b�\����Y�?[W�E�	����g�SV�4 %g�)�(���� dG|�\����}1"={O0����]�$՜e��]��Atu�7Ӯ�.��CE��P�j�#fS֕e�fو?�[�E�����ŉ��@�+�<�h�ޏ��ؗ�E�ܝ���Dg,����E��t��	5F~�z�@j� @Ę2Ii6�I���P"�	]���C�Cqx��(�2�Le+QV�X[F�D���ြND	���M�r�;�)����*[q����Â�l���s@��x�)��d4�BBR�a*�k)EK�d*~Hk��y;>�=�r>�Y�nD�3[���I7��BQ�|r���������f��S���q���/<��S����7&���[·C,/�urw�����Ņ�������]�8{6I�KV]_��`E��{��hjL|�FFK
x,��}I���ۣ�lL��]~�Z�I��xrDݰ#���C��`8���������x���*�+�����k��&���K��ݗYi��v[����I�7�Q�,eDLiBT&�
N�4�V�a�,�d>�f,�0|����(Ķģ)pL	��e�om�{�h�/b��_Q��(/Q���F<a#i���hY������}�Ytu�X�k#���y!���{!K�X�����<�gqF��R�ER��?k>WfF&UȢΕ�@S�$�a�6����wD7o\�jxϻ�����������lS���x���;|l��X��V��eL�3�,�������'�`o���<���|8�-�×^~�'wv��c)��ݣ�s7:{�%oxV�����&/��~�z���r}���ɣ��C���S��?m��7��Fs���S��Lg��+W;�][��|L��C~͉�l��#�\���1�,�i��G�T���뿧=Z�%��иֶ���z���O���e��_�����7���s7��p8U��M�âr��fe7E��]��V�!�e��QLk[�|�\��\ƥ��7M-��
��,R��[N���[G����Wj�i>��l6O&�8��ʚ\�g1㊠�ՑuE�fҟ�"�D�̗9M�}r�&,�R��eQ�Q$���D��x�>�,�N1ˣp�=W啤�d�0<�B����$�#>f��ӡs�'d�q�,�s.���������)?gF�۷h4R��%��,Ҏy�����M�<\����v����Ȯ��L��'�g�r���O��_��|��՛�@y�h�W�[;;;~coot���[���<������ng�c�V�q'�pD�t�=�Ai|�����?�Y_���-��p� ��,S׮���"�������^{>ݶ��Wv���a�_e����ݛ�������~��?��s�󉝝~��y��)?M�����n�(#����7DW ;:h��8=$�([�0��I}�\R�2P��|1<��F>�Or�y�XNi?NEX$�X�Y�sA�8=�y��b����(c?��`W��l���H�m��]���XȅQ �&�?� Y��(��뱈��\F���A�Zߢ�׍{�$����Ik}��"���W%���Y ɔS��ztt4��=��w�����T�"݃�B/�ud�-�9�A�a��$�L��qF�3OK
kK�{|`��6m{uz#ZL�(Kbh�������kW��������?��~AorΛ4aa����ï]�����я���/�I�Ζ�A7X�Gԍ<�(址��k\�c��Kg�P���x9k��A�?����i��S���l��7�Çm�=�FֱU��xc'�/���W?x������g_�����0U~4PѤ<,�*v��r�kN�ҨQ�K�L*�-�wyHYV�\8�T�LfR���%x���߅ߡß�1|uN�w�D$IG>·i�������0]�BBX!m�`��x"�:]c8i
�=�GB�n.	���,�����}�G"E䖕���٫�k�c�=��墔a�v�K���ƋL�4�v�ɦ�^@��'��祸�C#�UCw��������c9��Ęd��@�/��(����ޢ����x|H^Еگ8��i1�ϓYtQ4��!��[4���x���6u7�g�v�O����k�n~��/}۲����"AK����ڗ�u��;��?<>��R\�l�v���z�Ne�O�<�H&\㓄v��`mD~���躴������3H��ۇ����^�{��'��ss7�Wd��̘�׵�i5�^�PUe����7���|�[���?����헾���Υ��S�"*�����',H�>/c�Z"f�<RrI������ӭ�|�0��н{;4�)^$TU����:�@��b��b��t���
$��q=?2T�qetKM��̈&L���#�F��C!o�s]h���Q�������'���kEb_�c%��?���G�3����)^�T��10v�oS�,�|�<9��=��k��W�hclL�"����P1ڌ\W��ÎC]O�ߠ��[�H�aU��>D�,��h��h]���>t�F���r��|��_~ǽ{���+�~����o�Z��J@�����˷?gw���&���Ko�&�`��7�p/�#t�\��xn���6��PSE����dB2]~�k ����8y��$�{�ފ������OE�P���p�:�3+�ݨ��ss1~z�k��[߾���?r��~�ڵ�~I=���CE��P�'�i\��旅A�u}�p%Z̦��[.�N+ВMAQ���G�ٜ��ә�&�$D|<k,�I��u�"�}LF�X( ��,�1-��$ɀ^˖�n�5�m��0U����G["��e&�M��(�����w)�:�6�����(`�`�������S����VD^�ɰ^���������@F|`܊�s~\�Q�PJ�m�-����(��T�ce��2��V%�7�Xб7�'4�-YTZT�"��0)k[������{~(�U����r>�����{����o�إ��c7o����˗3R��A�ͽ���m���͝ۻ�����߷��bv$�b�0�����:Խ�IJN/�k���}�drx��-����9��=����E���$��y�Rޘ���⭐���H�I��n��'�|i�xtgv�#ߺ�֯����Ý��}�#��ST4)��n���N����V̖C���x,5BgϞ�#�+���8�����n�/"�b��HSV4Ҳ�&�G�}�)�TRo��(� **]23�\*-#ǘ_z0|n$ʅ�����Ӽ���)��b_ ��A�#��h}M�p�Ʊw⻲}t�]�r���J����և�F���{�E*���71p(�]�K,vBϓm���&�p<�X�M+�D�_@����!�`�������X@Ř�WT��)o��n�P���B���ˆ���yz&ϒ���^}��3�q�;{��-Om��O-4ea8{֊�}���G�kw����l��/Ҭ|o�6��a`�M�~��,���>]���]�����+��WH���ն��vӟ�3�q?�`¿�3N��Rض��5����| ��Q������;oQTn����Ζ����ƍ�up�����>��<~�;˫gǿ���7-*����O�a���i��CU]t�ʍ���!����X,��ξCg� �"C-�АrZ�HMS�;��` ј%g�歌��ba!��RZ6�g!���M����Lf!��Uq�nmy
��/�Y��2�*�����F]��ޢ�W.Q����l�bш�9
Α�)x?�[[RWu8�ҫ7n���=�_�D�.?�����O��Fgl�%��,�� �Z���Sw�I�/�u��	�N29'[���禤2-��}c�#��vP_5[�!g����
��tAY�HZ�	��MrÐ��DF����Lӷ�W��w7���W/�_�WY8夜��0��_{��ݻ�w��e��{uS��:�=�!���H� Ҭ����Z�doA
IE�k@F�v�G����q�ЄoS|�j=�!�V�o ^"J˿dQwHx%�ILv][�`��76�t�3������|���_|��G�7�}��ō�w0�M��&������Q��"���m����"����/Ӎwd�"J�k��7/��ؼ�G�z�tō�ϗb܈$H�cL�	 ��֒���Y�HҪ[β-�Hy~ �i��8����H1#� VP^Vm�ߦ'�^���p��<�<�Ķ�����f���0V����uYD�9#f��oݠ:K��O�3DŬ�$������xK!���qf9f�%b��8��b,C~Q��38��bK�ӡ��1��j�XR/rXxi������O�傖�ES��n@k�.�]�Q�?_L&T{�6�D��=G����W���[w�~coo�gϞ}��?���+�t�:�m/��n^����zD���T=:ع'׼�^��������~���y����i��8oiQYT٨ej�����1��;��߭2�>9H��>�k�]���G���ry���G_��K�~�����]~�O��������:�̓�&�g�I���,��B�|��ZGGGR��O���Џ��>B�,cS���T����;4�e "1���ɂ�H-�KH=����C�T�Z�V�4)��&�mV?��&�r1LU���8�E&)=��j��z�;��3��4����r�tC��iLy��z�C�����^�u�Ξ�@��:��R�{��K!�x����$E��� ئv�m��uB��B�����s�q�r�2�N,J^2z�+7�_r'b��2�CД��ˀYuH�,��ɒf|�{,�����]����%��}��ʒ�߼�s�LVTg��<�ͧ/m�a������
kя[��s^��y݈�Fq��re���L�i�_�H*�~�|������e��3�[�(�d�h-#��ϿS.���wF>$Y�G6��1����l��(�_p��So{��V}�V�x��/��3/�x�g���ؿ���?�����.��QѤ<T΍�{u9�_˺|v2=~��xl�X,�9s�:aB2��D<َ��	uYZJ�͟�B����RW�ѩ�d1e�;��$�A%7˖�a���-�J)����e��u��˿!�Ɍ66�hsk��MX|��aa!�x%�]%m�T~��{����ł�	3�
�����HXj�<p5�+�=>O>%����iN�,�����r��[���Hu�"��6���Z�|}ߖq/��_T�'|��0�"4�Y,�4_Zb�׹���@��u\"�t4�9s�R�;��l�����������;��7>0=���������k�IR��������"���m���L�� ��Rq�/-~>ֶq������a��=q�p�SK�{�V��Ob��>����nV#��JŇ,��y�	׃_[�K"�MeY�(������`��W~�Kw�~�S���Ǿs���Om���M�C��{m�����?��Q�w�� ځ?d#^�+�d�L2((�F��e��T�q�F�	�HR4��Hל���@�ء��+YD��5"�d�X����_��忍&�A���)o�ӊ��-�N<�W���`
|�������8[��෹�AϽ��9Z��O��R���%Y�U��C|Y�W�s�H�O��S�N��:Z���sC*c��X�\��n�̀��%����$Y-�X�T��9��G�k��g-ፕ�r}J������yB�n�x������S�O���q��������?���~��,Do[o�ł�ߙ���mn�t���X O�1��T�k9��}9���������)���{��P�ý��ݽ�?1o���?<5��ʩd�Q#Z��C�d�-�$�I�䴪�leP��a�|���s\�V�Fg��Rz�N����o���o����ߺ��O�<���?����{�`���:l���;o���ݘ'��P�H�E�$%ي-Y��ĩR�SI%�T�W�#?�5T%�3���hRIp%�Sw��@��7���y�^��Ҏ�")����.���;�{�w�����^k��<���4-�}lhZpx�����&���
�7ٶ�Ky�%��ʑ������$?�X�t!y�U.�tY��� ~ `��X�^6��+t�U�B/�J�?�|#)/T(��R�������iB�'�|��]��9�(���� 8���R��]t��vMJlX{��;c0���i*K���&?����9]�;����h�2p��ɟ����$�8D� �3�N��hYb�a�
'h�Q�����e��1@�&D�c�����:����d`C3��?���a������@-
�N��Vw���߿w8��3g�v�]k>��Qmeq�4]��[w�nђ�)4�0s�uOʭĘ'iZ�����ywv���w ����ᛮ�
�9�Ȍׄ(�e����� �\��Rqeg�)�#�v�i��+)�)��Y%<����<]�5�+����~e<<q�o�y�c�}�[/����]�<L'�W��vo��M��#kk��U�o��>���?�O'�Mk�s��mYH��.)v.;t��ȮO#u3����Ґ�z�ܣ[� �BGL�f��*���⿣�_��4
�=w�rM�c�肎����m~�p<��h������?�|t����n8§B9v/Q��^3$�o[��QBU@��1�#�\>��B�,��hB�Yl�ۊ3d����R�Q�S�b�Xɤ1�!>Ou�V�
  q3?��`6�E�%8�%���:�,�I��ŏ�d�F����)�����O+J{S~?d����6���E�^w�4M?=�~ҟ�?��S������'��aU5�����<�l�靲05��{�)-���׏��4�*m,ô�]������Iy�-��a|�(9um6��a\�s���`���#��iST�Jt�@�,��s�I�M�L��Ha�V-6S��=*�A���̶^��'SVM���jZc����/=~��=r��������߿8���v��;{�/�O��M��#����3�ww�����O�0�`��תּ�e�mC3̺���x�^	G@嬼T�m(둮�K(�U�&�p��X����)�����o���lT�I���մ�2~���� �"*�Q�2��ŝ��s꠭�q� fKg�e�B�6�~Y�
�	�m�S��I+B77�r��~@s~x�k�L�?�tFyR^�m;�3%���*WR_@�Ǡ��e�ԓψ���N�Z�G�Х	����`���AH��A�֚45u!���`4��?�7�����@y�n����s4�Z�D[q���_z����g^���;Om^�gQ�Zړy�����#�~�d���k�ꔵ����!;�,��Qk;GAР%h�;���ʻpn�Ã�|�4�	oL"��$!K�t���$�쑦2إ�(�!{����Z�:i5�+����ʍ[6.�I���{�FЦ��8��5z�Z�*[��o�}���g�����N|m��֗U����-EM_�c	���G>n���b��.M
���п?���q�~s�kz��J$!X�2�� T�;HC���s��v� o���vR���n�\�Q*�'�)ƹP"�g �L �)�(���'�����vMz��@�� cI��=�O�Wk�a�����!��|,%J]c3ML}�7\Z+�RQE.B���Zߤy��8ȏ#q ��xC������� @rq�� ��]�J�Q�l6��÷��A�f˿,�9A�=#��KW���Ө��8<���$��i���
��.�	Ɵ���*��5k��|>���t|��g���f��������A���,�'���`|[�	���'�[r�����A����R4�6A�6�L���]Z�x̮On���͍�ҵ��x���X���Ipǽ)ׂr$���=���n������N�!��J�<��6E�aIy�5��@v$�1ߛs�@�^��z�8�;��w<r�c�������+�ַ�<}�R��u7��i9^c����"�-��W��x�����zZݟ�M���1̱ �UD��xd)���*(?:��S9/^(��6Q��,�t�2N�s(5�p$���?�J�M/��6���o�z�腗�ʵ]2m.��[����2~��Y�DG#�@��Q��Vs��No��ZIU�CZ1:���(]jv��A�ƾO�`��-��P�Q���)B+�#̂�� ���i~^�T�pW"���{z���砆g�J� Y���D�{H�R )���I#�<��;�)�HQ�+E��WY�-rQJ^�km��K�=��[�Z������=��zፖu�%��0����dE�W��T����g�ye����R��T� r�a���v�}���Gw��ك�����[crL��(�I7ߗ���'�x"N������蚢4�ŕ��"���0Y�̖�p��B����f<��_tk&eaLoxl�e�$���Ԩ�Hk:��������K��鋳��߾r�~��qj�}����xy�_c	���55v_�y�^����˃�0��H��mi�ݪU�	F�i��a�Z��#/*��\8ObS��CIIB��Y�H�o5G��^��B�ːL}!��Z��C��~Q�^�B/�d~�ͧ�Swx1�,�d�[΃���
p3_~My�'Z=�[��.H��D$0N
jt�A��J�?��5x��h8:�Ş�H�I������WKI2�e(�ٞd��zo�O�z��M)P�y(��܈s:Q0��xV�@#J�����J��x^���ίt� ��98�"�`ۼ�9vZ��:�z�����s/�����y�'��fh;��MP�UՋ��?1,�p��,�w1�W����u���nCcx�[K��&��(��/]�ݻ?�>Vv�b��4�8	��\Tk��R#��J]��T���7�Zk��^����i�Jɋ`��j6Ņ M(Ж����S��'�ry�d����$#K�k^�Q����o}��?��k��C���g�w�kܺ9Y����4-�kz,��{x��������&qg�M���2��d��S�f�����TJ�@H�����R.K�22B
v-B�^,���P�h>�{Nߴ%
�uע�;�T�I����vM2��Z�m�O'RV+x4ZMlI�P���cc�V:MY�d�R���#aF�yFe�J��}�����^w$ͩfU�`]�N���Լ �d�@�	�!a{�c�"��ƕ H���lh���&ǹ!�qKN���@�b�����q�5e$�����X��u�̓)0~ ��[=��٭N'����MƷ�y��o�^;|��K_��ĉ�׫D�Ew��5��(�b�T'M��
��J��֬Q́]�6�
K��4�J_�%h�A�>��L�O���#7���&�IF�MapH
 �rO�Rz�!�2ѢA�A���@f Y$E'�����G�|ŋB�
M% ���q�H�[�%��t�M�13��D�kK��	�TC 8���*���q|����SO\�?r���7�������KK����X���x݌Ev��WW/]��W�a;)��8Lo��i�ߗ��-�{�VY���E�+!���^�b�T�"gK�Iif�x��l���j�g�a*rP��"j����	��6��0T��I����As8�z{k�N�EG �tm������$�KW��K�wx�Z����EM�Z�hm�KZ�A�f�9�y���Ç�ĥ} i�R�L����nq����-�$"�Wm�2� ���N���  J�lQ(�X%�|���M�04�4 $*<yE� ¯��  v�s��C*�>u�=��[V�վ5	�����G�;��W�����vm�бc��멣�� ��[��?�J�2MC�lg����`tH$�yX��d���L#4ʛ��h�f �j�����`~�j����?>/���o�Y��x2V����5E���7'o�P��D'�B���d���� ,)ە�3��L��ec�,0����H����HyH�[����rKJ}��$��%��:��\��w_{~���]?x��૿���z������e��3��i9^�cd�����"��rn���Ma�5������-I˝��^UV5]3mݵ4@X@�e��� ^����b ;7�+=WzMP+�E�?�Ȅ$̬JH�j��R�V�.@+f`��o�ק��K$ldyl�p�slMF	㒌h&��ҵ�t�E��K��r�n;�M�Wy]��6���į �X�����2��xx��{�yr����u #tV8�|a�bppX�m��D�T݇�T+D�fA�_��
:U5ٱ����5�m�#��g�\�3�~�ik���ը����$���}���0��t:��:xB��x^����QBf	�8[tjZ"���Z�F:� ��dY���4�[��������\N?~0�O���A@4+�� nQ&|ð�X���?�)+ C �υ@(C�����3	v�$I�-J�"�d,Jz*�
R�λ&��#!fټ`�	È"�@AޣwR��}�	��M��1%�*u����6�,ژ_:z��+{?��k_<��?zj�:���F��<��i9�0CS����=5�L>7
� �O�q~k���f9�9��m�ݪ*��2 R^҅�����&eq$Y�z͕]k^�td<]wų�h9�F��,)m�C��g��sL����ɥT`����d&�W�;��}\������&������]t��&��]�K@��֔E�>���:2 �����u~ϜV9����d׬[ ��(��QA���O�(-�>q��;y��$���Y�|��� N8��BF�Eq�_oB4�0J(
걐ѓ���8�=�z�u=	�������:;�����_^�|��'N��5:��n+���)K�%mȁ��1�/ (�jY����|�˗3��W�iJC-��5���è���O��tD�a���Π�ᙔ�D�㪅m�&s���.Fi���Su�q#���'���T�	C��*U�F'*:W�3d���:<<��� NC�������-�W��1 ��S	"��k�X(�gV\ew����gZ�?�?����[��_~���c)�ZKдoȱ��LHu��~��lV�"}+��� �O'i��4)�,�j�0�>/t�nZ�k��n7^t�ӹ,��^C�� b� q[�N-�&��Ż��adb��0xOU>C.��t�b]�x���Eղzrr=(s3��n����F+}�NF�n�R�Q��`HU`Q˳�8T��i�MVU�B��A
vэN�"^�xMZ���{ԮYJM�wt��wDF�m�l-�uɨ�S�e8�2D��+K��ᡇ��c��ɟ�4���h(�S�~_��a8b2�5�.U�ԍ����N�g�ǂ(~���/�~�m?����kh̪j%���2��T�V�����J��
��
��:�(HYh�T�
�ʦ�4TɓASaY.�����V�y����gd섺��i�s=�s�o7Ăh8���g;�E�e�𮔦�� ��؀H
�"/��u�BT}'ZQ�^H�(��5���f����m����'����5��[�%��r��0��ESD�p�Y5�7��e:5g�������'�<0����7��2��Ԙ���ˮ��X���xÏE�'Y<��z�A��5���Zy��(�3
��y�ߤ�MF�(�xcx����@�����d6���C�1����:9P�ƣݦz�I�Z�פ<7$m��D�2X.I��L���N�l�J�Ɠ�c_D/^<��V��h��$�%L�$���2��v]
yUF�p	���$"�A֚W���g����t4����j�E�mIY!H
eˢA�I[�Ϩ��&�7]��aC(K7u!���
_��PV,��!�Ҁb� ��_�Ѣ�ʺ2|_����W�=��D��7�?��F��ܿg��?;���x���}m�i]w����(I����ү��%>M "�S[]���z�ҡ)އ7���r�	%*���*p]s�5]�|��t8��(L?1J�f��
s�魭-��M:�L�<�'��AcH\��P�@4N �j�!�L��9������8�-`�dI�`�f+�R�N��2,�A0�=�V\���Zd5�B)��7�<����<�Z>�)o��iL̴u��9����{G�G?i^��uW��5��?����~��_�:q�uZ�x�y��%hZ�˱؝E�8Q�@��d���5�T�go7M�ci���Ҍ��Յ�����J���4R�Ψ��Es�R�������1D]�u��%�$��H�v(ED8/�Kۛm�Xi�p�|2��y�נ�imv� �R�b;�#���j�6��e������Z�ڽ.u:=�gs�����^��xDk��.�i��8�R����e��ECJ�8�~x��K���tF��͠��>��ǻ�X�PM�����C 
0��s��k����@�gp�5�}T:n���O��c�뻏;���$��&�:=�z�x3�C</jAL?����{w��R<�J�8j�#�	
d!�s��s�g�*�� �E�IF�A>Փ��j��Z�{OTU����O���� ,�y�00Ѩ�s�5 ��&�K����T�1o*���_�U(���"��-:�T��ʨ�]�YV�f5J�B��*�v�Ϳj�F�~1�?2s�ԬvWJ�zi�}�%]:_K����ͤ�Dq
q"C]V�H�X���!��fߚV7l�ԭ��VҌ�Hf���l��]?����s߸?�;��ީ�e�UKд˱�՝7�@y��|d0�zxx�3?�d�]��ԩͻY�t���yW�n1�
]^��0���t��y!?���M;�۴��Jud���3xG�ky�
���QPJɬ��G}ED6����\Jev�.;`���<�1����������o�'�y�=���$oT�V�I-~�t0���#��M�@�R�HdJ!&�(�� Ú/���~��/��"_c0�LZv�i:����(J��]d� 0��W9�<>^����ʟc0�j,ts4Ad��9f�w��-�L?0�Ӄ��Bc�?5lz���[U|mee%|�3'~��A�����U���7M��.xŊܭ���:���خ��o�b��>�:�AG�W�r|O��N���S�8o�|�g|�鼡X�ؔ�3Ox#�Q�dTo��@"@>���?�9�{���2�����5��� �$���*)�X-�������a�i�̟χφ�^�t��{M#_w�}+3�\���`���
��m�:,5Sx� ����d��k���Q'�Fߓ��y�Z���&�W���Ń�3�͇_\�<�дz恶6��xE�4-�r�'ƍL��<����x��������ukB �10Z�-��k`.ivp�:N���堙���]e u��!?ϓE|em�V�7��lP��@�_Ӱ$��Y%�9�,+!dd���D��er 6x�*����� px���n���P�ۤ�hFGGG�@��6�Nݡ.��f�&?�!I�ib*�sj�e	O���A4gH��~�[G�Ǣ~m����&��;３6�{!a��9���"�4�����.�{�C���R�������G3m�����c�<��Q�5S߭;��#����տvM�yP�+��7��;8 �����eX6r|�
�*��'4ǵT� �}J�A9���ex�d��B���N¼�W�e�w]w�;�=��!�����:��%��f�dm��.��I��)M�7	�Y)���8��6_����Ì7(|���5T�\��9��$�c���u�1ڈ<�� �|�k����f�Tn2}�������'�����݇�?����n2;����Xk՚F
>T�s������T ��țd���\��(���3e��	�5u��>Ҩ���y�<����<~_8�嶧=���z�����һWj{���+3��i9��?3�/����s���J��]�wu��-Ev��8s�D�Fy���Y]ِR~ps4���Ч���:��x��w;�h7ȩ9��7h�ې�βD:�4i��ȳNq�s��i�6/��8EhΝy���Zt�St�x�R�F���QH�~���z�r�ن4Ȅn���`Ï�`��*�[�pA��O���=����n��$����+>�m��:<ׄ��n%��4e7��J� �/��ik�rs~��pD���VWW���h�~M��خ����a�һ�0��ĵ=�	���]�y��pz�4��n�j?�@ 2c~�</����H���ؠ,�i�6��炫���R%3���_��Se�2�>Mc��n~�2Z��u �~y?}�h�~p�U�Y�@�0D��S��ep�9ፀ���jd��z���)g�)#GA**��jk\��L�[�&��T�� !k�^8	�K/��m�����ַ~����x���^|��3gy���ώ�����Z�l��K�2(r���I/S1.�b����7 �C�Ԕ����*^}�c`���ưȽü���'���Y^�=���K~�Z���X���X��a����W/�F6��I�~����մBSD��	0m���[ͥ���_Mu�i�#�YV�d��l�t0���!����wj��ѧ^�-F��V�Mi��S��hɀ[U�;�3��!���h@�񈮼�<�'}��ܠUg�">%G �#b��e�1C�۵k�-�:�d�R��.�Ƽ�"��v���55�P!���;ٚ"��`���n2� a@����Җ*o��г�}T�?lo0�yZRs�˹X��Ro����|Ќ��f�I?�q@�P�͇�i��~v0>x������������$0��;Ҭ��9�}��M��J��� h������� K������wL�U��x�UZU����?�F��{��3Sj�M���|g��Z(�"#��
�z��4������9 ��Qě� ��'�{�i�mZRJw���0㍅/�+E��d�yj����,��a["�~5h���ܐe��k'���o?�r�u�S;|�j�{s��c_{�����t��d�-nw�]�n�g�x��d��Ζy� 7�7)�Z]��L�D�L�jր��?�B�c�U�d�\�y8�S}^�[�������h	�^��M˱�� ��W�����A�����FiF�(�q�4J%��E��0v��N@H�09��B�3��FT�}귛�l7Ȅ��gϜ@� ml����&y��"��*8CFG�$�[_��αM�1FCEF�gB��Ԍ�#���[����n*%�Ȅ���E�S˨Qe��P�'���{Z���M�vG���VK���J�1����C�����P]w(�� q����M%���:<�&�	�oG�%LJ
F4O�W��
�^{��`�߉AL�YeYu��씤���9�M��.����|���_��nWܢ������Rya|�%�=D���_|L7�.� �I��(.��Ȯ֬K6BK�1']�<H��@
�Y�B��^�כ����uZ��i����Y��q\xAS^M#�N���\��R��T��� Wt��IBa2�I��*���T�y�%�Ϲ������'/��-�(�	@6%�%�f�Jw?ǰ�X�ǹ]���OHG<�#�'����\z���<�⇟�������}�[;��2-��bx����-�� 
ɰm%\+��n�A���JJ熨Σ�.�Z*�\3����-uq�\�W`,A�r,��1][������Q;��,H~�׮��e1I3���e	Lzs1�؝��J�%6˰��;���@�p�$��j�w�]������@<��_�RxF�`;;�h�ĶdwlYT)N��b�os@h���\��1,4�/*�R)�9h[�� �䘆�IY��� 	9h�g>��[��A�(��C o�i�Q ��5�}��C�@���p�@�)tŋ��ad�J,e.p�x��)��J��YLo�T�+XN(��$λj��YD�yD��X���ٺ��8�̣L3�¬y��v���k[�V��'2��x0��/L��� �t���Ku۞�y*D���|�k���J������&J�%aQXg ��T)�>e=�9�@��[��{�<pM�8+*�zf����7�q�c<>�V��Ma�'''a��0iI�v�l>cߧ)��>Ü���锁���I�V�3C�t��_�g-V��_O��c㒡\��z��T�\QYd��tA�n;�׎�M�t����SƗ�i����o�c���O�3����������_��#�p噟.������N��tBJ5����1��sҕBy�������֔��Xo�OHF״乨��((�iֲ��o��y���Kд����-���Ӌ�$~����]a�YZ^IZ_�EDa��i(Jl S��)V��mnm�,��h<����++�f{C��1�E_�7�	?���t��3��>����~�G�z]�KY��(~��.:� -`(n@T����@n���E�1�)I�У,�l�4ဏ.�0��LL�F[qx�5#gA�,E&����u�(�/:� &2E�Eg��0  �[�q:W]L$i(�� �ٯ׉vN�!����L2`�]p�3@�p|���:���{�l�y�s���`L�V�<K�j�U�\�m9;�ޝ�i��ʟeE��ı:<<�޴,��#��:������% �3�cH�R��L��*�d(�&�>W�28TY*������^�<G���˾r��h6o�WvĈ>-u�-��-*yNM��b�|gUٌ&4�#��.E�M�F�j�\��OF(�[Ҭ P��Z& ���n�!�z8��k%R:%V,���5������<6N~uw�^�xg/^����v6��hU��6M�8k�V�����}��#_�����|�g�z�}�����5�HCcƌLޘ��N8s�&M��Ն�.
0ir��3(�x��(󴌧�Ko��������˴��X���X�p����������^���S7��q�1t�"K���<�e ͏n*]|�`�q��uZ���h���c ����N5�CE���T��$9ɜ��:8�N/���{+t|g��WVɵ)?���
*�D�F%����v`�R[��r�HE*��0�YB�C�/��^YH��1lT|�6��].D�]ras���35%�k�߹A�9�)1�����A5�*90aG��"Cg�A�Z���.����#�f$��/��z��Xʌ��fɘ\+�n]�Z�Z=�7���^T$|.M>�-���;�i8��;��T�d�4�凘#`��g."����!׳�c�n�wt	J�q�H�n()A.�}"򙦕g;���"����0���}G��x��<�t���8g0>`�4��7�?0��b�<W��fEU<J���F��H�"�E�C��=��q�E<�]j��Ik�E�i�sv�Y�I\�Ś"��"�cp?�96����y?�}t���z��O��܉��3�/|�����O����ܙ�O.�?��CO���s{�Q����d�r�*}�EA���0�)>H%�� Kͣ��|�m���[4-��xE�4-�r��"��3x�ǩ�`X�8��O�Q|*��6uWZ��*'S�镀 �X�t^��E�:l�w�����nI�VC��A�F��&:��=���n�`Z�{���*�*���v�#�p&HKy�?ԸQDC`A�ᭅF9~���(J"�9��@^O$�|\xm�і�� �)�ndfJ�OB�քǥ��K��A@���Jq��/[Y*%f���Y)^\HBM�un�=P�Ä��1��	E�w]p �vs�3D6�Q�fK�`�ρݴ��%f�ye���N+�u��;���� i�*+)}T�i��RA���v�9��$R�y�^�:J���BgW�He¯�s���eы�N�_�qz����o���$�wo~x?k�ң��4y|����<Wc��xP��� 8	���6�L8P�/T�\���K�&9^�|tC$�E������S�76ߋ.�+���O!_�Q��3��2(�|ո�y�jQ��IA+VJ���;����3�����o=��fwm������KJ�/��_�_���_����ˇ��T5�}��!����M�o�l*f��j�����S�|,�棇o?�����{k�h9^��M˱��@ ��bY�������p�˓��]�6�4�H��X|�uR�q��%(�h���;��=��Q0�v�Fz�M5��P�5T%<�,j2pi�=]�wzqt�.^�&�l�펟ؖ`����!�<]dFJ9�1D�F_��?������&4mG|�逃Hv'|�NL� e��Z��B���(V`BSR�o��Yh�p���Е)�nH��������@��d���p�B��@Y3��v)h�4R�F�T��t��DQE����`S���9Ԭ���6(�����4Wd6>W,��@EaX��0�<��ߖthY�&)&�ps�[�5p��M����Dw����;����`h��_o~��B�q�����_�3��GФ��Ъ��d|��T�XXz)�?	|*yn��j1�^�j����)�&�|c0{�O�[w<���X�lb�nU�����"��I��#@SͰ)���ƙdRh���m;���N̇Z؞M�\�_���k�ߵ����z|������]��m��<�ͧ~�z��7/��,围�#�S�ͮo�4ː�	��$Veu�a�	S��0�����|��ew�+;��i9������«������x�s:��煸�� <'��T�BѾ�sP��R QtF.-��4�D|4�(��=Z��g������=�j��rEΜ���K�84D�Ad}}���V�PBe�M�d��F��:�tr�����*
��a� ��ڒا��/嗣#����n�Rf����V��J�z�-)q��qI��̅��]���Dl���6
�Y�~w��X�d�4��b�� 8'9�׃ќʘj�2r]�u���- /�":/**i�'T�_ Q\�R.1 *��^��T�Γ����D���A�JeΠ�3���?��?�3^������kkk˲��8.&�FA��A������up���D2���ɏ��,�!�*�BYRا���=]��1��5�,
`��)�&56��s�!"���\ǫI6I��RJh����Ű"�Z�!L2��JtS�:�6eE��Uq�A��޳��������_��������o�. ���C����c�3�_����rNZ�	��l(
�)D�p��	�Cc�ek	�;���}��>񶭥�+<��i9�����,\�<��$��?����n�,�ɋ����;Y�AC�A9�^��$��l7�^������I�@���A���C�]�)�.<GJC� �.^�D1�B��u�-�hssS�[�;���ޜ%)�\5,+� �����f���`� N���HK�V�2(��&�L����u�i.��/��A5�XT���r�'��+�d��j�b���!ZW�쵺muV�GO 3аq�k��x�hN�a(]�ݶ"�#�Vҽ��i0$�A[3�����n�B~Up��	�_�@H�(M����rd��+��4�8	*>��z���8��$�~��jUy_=s����'F��d3X�x�E�)�2��1p�J7��*��*R�Ff�v(�xT���@��f��4�)�t�9y���6耟�3H��	��'<OE�<7�K|_��TX��f���R��{��M*t�Zg�p�*]��Ұzm��������'/^~�[_�WO^���'o��kSpȷ�����p?����%���gFV�FM� 9�l�w�L��*�{�y���|�f����-�+>��i9��U������u�g��I��8�?E��(�ݘ|Mx�\��=@E͵x�X�2C��@�w�E��2@��a>ץf�% Iy�-�߼�AG�Ĉ������')�tpp@�=���Ѩ9~�mooQ���R��2@�a30s�#ٵ;�:��P8W��qL���6'K�J��рQCڻ���?����a����C������|$�	]?�*!��A�Eyf���OGGC��Z[�:�#��y@��kz�4j����H*�!)eƊ~E>�����4�Gr��V��i:|.:���s��f�Z%���� B�TD~s�B2\(i�&|0h\��eB� Z��@���փ�����|^�%��??�e�ʵ螃��3�8�b@+	|��AɄ�<M�|����̅�&ZF �|z�3b��2�� �M��,M��P�.���-jw[�1P��}�Ǒ��T���*;�
��ՌJ�wpB�B5>�d���74��TG�Uc�� ��.՜��w��,V��p��{���կ�vӉg����{?u����#�T�5�@�H�a��s߫Q�:��x#�����ԧ��X-���s��?���r��c	��c9^屣��=���o�f�_���Nf����9�t�D�m��#Kee��mY * z��WYu�N���A��{˂���DA�fp�l�x��k�޽��M�n����*�<��E��١[n=� �+ �&��o������_wMr�|��r���ذ-�c�]<tb 5P拲�g�t�� ��2�E'���8���8ēu%�'�3Cy����	�ti�B?�͕������4(�1��ug2x�yuj�=Z�]��ш`�����0�
�|d��i8�ly���x�� �$	�k�T�;���;~%�:4�P�bz��r�3��0�F||�������_�̢c���#�����Fc�P�^��h<9��5��aZ�>C������0=��Bp��R6E�&�\t|2H�b��'T��f���,~/�Є���`� X�u��9& ��ᾈd&Y"��a��_�,��e0֯��Fw'�����~:�t��^x�.�]����ұcd����m��"�k�@�{�\���߁a�� �s���s㥽��w�=��|� +����A������ 5q�	��{=��Ȉ��<N�j��������zu�4-�r��"�0e �%Kk��]�o�$���y�&^�M�44d0�$')����<GW�N��������J?%;  ���h���}Cl���T�QVC		"��FG~^ԧ�]��O��P�&6�V�����j�%��l�R��e��l�;�R��A�FW�Qh!���8�]���)i�x�R���&���ҕח�4p�p��Ez���D�a{mC��
�6g��
��ۮ���BH,��p8Y�:q�ASFSީO��` q��:y���Gϣ��#�����T��c0��J%t�9h���a�l�@)��qQ%�� �b�q�#���L�heI�M���ͥ�p���q𭃃��L�8��z����t��xݿot��@��-���H�����^i��<U
p���V	�) XYtkfvM��Ȧb�aXx�Z�Mݵu'�G#���R����lb���2�� �ϛ��^R�ߣ���=���������uz��st��*��!��.���<��b��-4�t�>��{$dؕ�ZeǨ��KӴ�G1M�J�J��2a�mkJ\5�cNѠ`��7)��)i6���73a>=:��۾r�m;Z�We,A�r,�q,� gѣEU��i��{�v��^�Z���ߡD-���8C���j���� #!�4Ϥ���9�$ت�W�A�Q Y[��e���j-���R��{6�]6��hL��K�^Gu�5k�.� Իs�CQ�F���%@�R�E@���^�σbs��:o�{	���E0c��c�.:�P�A=�)� �<����I5�|��+�5�j�!�>�3��?�4���׻�th4��h��l�G����@���L&�R9�N��u[}����bXS�du+�k\���JsG�e�	��R0����_�v"��E���m���7UeqwV���E��ʨ�z|����V3w�f38IgL3O�Կ6�?y&w�BO5�L�!e7 ؐA0�Ȕx�b.�|'NZx����NS�q`��(ۀt �h2pщZ�uW)��|4�K9�0Tc�00�A�n�&b��P��˿�9/S� ���Fo��4�<�Ag/\��.\��{�)f��ء��MJ�������N��m��Qws�
���F��>N�P2������Bg)�#x<_M^`���Գ��|k���7�v��Z*Ϳjc	��c9~�b��Y�/����q}��͟1Ms��*_�C�t���)��E^JWUU�����6��(����F�	?�N���O�ĐJL@񳵕�8��x�<g`�ƌ���(�������F�VS)^c���@�B���R,���`�ֈ���#��9u�G�䡌�A(�f&�ʘ� 7y*�O��]���b�� ��kh���|T���i V�F���P_��
syG^�`3ӡ��G��N��uR�I Yqp�%�'�1�l�mZi{|Y���OӉ��hJ�e8��\�l�� <|h��c��9��1�+sS8.5�4�aةL�i�ܓ�駂4�P��9m�_�d��/�O�7����;����Yz���|x���y��«���%)�?|��楮t�p�Ea_�q�3�
d+3���*�\|�,F������(���M��}��{�	�{�L̪A�
f<O���̇<���k�!�*D�`>;$~D�V��u�mtۉct��5z��:ؽB���T[ۢFw�ݒ�BY%�KV�vɭui2��t3PGs��Q���P���	h4�8]�z�Yi~�]w����w�}�k���X���X��Xd�3�9`�󍑟>8������C�ev�uW�Lf�{��P�eKW%����U9  Y�:Jx"*�Q � 
�'�-�Pf�������w������0����\?��4�V�%]x 1uޱ�N�Rq��
F�<������aF�y$F�:0Ea�AJ�V���C�Kz�+�:��a�|�բ��*��s�ϳ,b.`R^�s���MI�qr`j��ۑUҐb��s�������fҡ����{B�(����P������69h�� �4�5ڤhcO� e[�l����h����..�ɔ��K�tH"�k��v�v�ZU�[|m��4�`?(��bTΟ?��O]�z��kx�����ٯ�ܬ�?|m�Q���s����sm���K���6�����W��@��D�^�\閔M�$��\'�C�B��>!Y(��M��_9�y� |@ͦ�?���_�)m�:�u
����\x��lV@R�1�A����2Ze�u��t��q��'��c�_��KN�d6{d�Ɓ
��"���[%]�CJ�>O;��q���u
�D2c:�q �hLp "ˠ�6�ɝ'����?yﷵ%��UKд��#��!��?�V�����G"?�� �޶��m�qd��X:ِ��4e�!���>�-R�cPeZ�YC@:��=�(��t$�$2�E1���#)Y�4��c��'���#<����d�fAHG�	5=�n�٢��9�W z�N������I�t9!q�rLW	iF8슃ɘm���[�Zc�g4f��;�=t� �r�0
�LMv�P)�dR
�����S%�O �9ZX^ ��}�_��J�Ǻ�`P6�2:��4�w�c��U�"�;�#���>����9u�z�J�1�T2m*;��Sp��z��)�R�
�Yb�
O�R8.����Ʊk�a�n�|��Uv�����G����(����<
�tu��3�9Zs��k��?��q���ׂ���L�̞�|n�d� �2��p��	�/�ݥ$:���ހ����]���R�u���P��\j(	�"#�k)R|mk��h0��t[<����3�n�f��{�x��*$5t��P6���������7�~=��%z��E�8u��M�SCӂG:�����B�x�7v�t7P��TR�����ɯ[�۩��ߺ��?z�M7-;�^�M˱��� ��8 �ѵC���?7��?ڨ�w׽Z�Ɂ\�=q&���T�vS��;� ��B�w�{� Q"��LSف����Z��F�?�&H�����䝷��������ke���=Ck�6������fh���#�����g�f��B0�+x��<d�.E4���֮�Z�ͯ!��@V-��R |%��!���'�:("C�G��̯)�	񽃙�n�N��$d�J�e�ф�E��eԣ�dJ���qn���I����\������;J��A����1L�`�g�j"S�߱�9�s\�	�* )�9�lT)�-SS�/�g�.:��4�w�4��k��(J>��s��F�׮=�y���L������g��
�r��tj-��{p� ��9_ D�d��"���z#�7��ϫr��0]���t��}W	�5�*��T�|A�B�RS��*��6�	�6t�2�� ���+���siϒ 
�?�s���;ik�OO_�D/����=2�J�1͎ed��L����T)<������6W�����}��y���UKд��(�0pyf<�_֌��4�~.M����Ʀ�o�qGADK@I&�i��- �H�����\e�d��;d��yj��T���~�Z8��
�(��_lQL[#�4P���/��Տo��h��\�.�0j1��ڮyB�8����M�d��6h(MGCJJt�9�y՜�E���2I5g̄���D_����d*�� �D�u�{h��'WHp�S�ҥQs�4\
���8���l��oӯY��V��ui6��n�Lty:���H�єϹ���u�s��E+d 8ȉ5����� �ViIYIegUV,PҔ�'Jy���J�݅����N����*wF�H/�����`�|����#q��r��ˠ���gWF���'<)�`�!~n�(��&���B	�"�j��R%s@B�Ҍ -.ZxVҊ��5E����$��
�2�%�:��Z��1����u�NE�QK�z��Z��\�K@�LJ�Ȃ�jk���cd��Q*j淟X����t��5z����<�9|�9nC�*�=ŋG�{��T�Q}����_��y���x�۾��;-ǫ>��i9��58�K������YX|>��2�� �c�i؞Wh ��l0�E��]1i��(U`@�v][:�?��f��!�&�X�8�{s��.��������
A���[�b�#J�3�>�B�[�D<3
��t��Ur<W��k��[���fr�y�V�M��'S
�B���lj6�g�娸a�����;|Xb8�:#�%ӄ`���$�T6�Tmv�⩷Б������2�m�Z���B�a���D.����U6���t�\SD8��Oa]�.RV���׺(���D�"��I&*��8b.�T_����]�T��.��� 5-�[��aif��B��l;O��se��/j����]���Gt��t�3�}͗���;W��?1��YEZ�ױ�ԅ'�1M�9�&b� ��$34�%$& ��m�x��3 P��KRs��G�C5�VR>b~[J���sB� ������Hl�6Z�C���C_C�Ra����I��#Xs-�MN��1пy�K���h�+���]:8��'��k?�9��ŋuɆ)Ї��yΉaex�����'?�K�YZ��X���X���X��9��}��p�#�O1�y��7�i�u��q�����PaR���Bo	�& �i7� KY��Ȟ@$�B���a;��%���@�Q�4I��t@�}�\Y��v�.���h��e2�CZY۠N�lϤ�ں�:-��i4��`<�ס$���b&��h/�h��8Æ��-�5�pٗ��yb�_(K��7E^�DKV�t��&�ĀXB1D�fåzդ�?�c:<�Vn�-*H��ҡU	��)ZA
���	xK�X\��B��{��f�qn��s�ȧ�ħ���nU��z|g^�eٶ&�P7u�,WʼX��{_��ȓ�|8,N�'/\�{�&o���v�Z$�_=H�ޛ�$��qe�g(Rv��<���wӔi<�Q�M��d�=2x`����� )�Y%¦$��nPJ�$*#\D$� ����eP��E*B����c��*�x �IN���ACMS�w� ������'d6�ا�l,�b����a`v�;�ݽ!'
���I�Ԩ�̾�%]��᱇��箞?�����OkK���X���X���Xt��x��ώ�����Oۖ����oڎ����vВAiM�H��)K%sфp�ա�t"�	�s MuP�<A�F9�-x�)^l*Y��Ex>
�R&|����t�0��X����h4K���� �_Y%�q���z�&
��q;t �(��-R*=�~�9qe�d������F��\4�	*r�)�Y� G�+��7 ��1���%�$�T�).�<«e1���9�Pb!���h&҅<���Y��B�)"R|�c
���n��,]�H�Z�:�`��*W��}���~�u���`-Nc9�B
�ӽ	�<�b��`�Ϗ��e>�����LΜ�0;�╽�l����vk�Z�@�9�^|��8�e��z��,
 � ��\��,yr�X�@���u��3�@�&d��)�1@1�\k5OeIA���<���#\7p�ps��A��ފ|P�|�O�k�l`�G�w[�l)��@��A�#&��������	�&R*^i�h���'u�զ�w��^L/�t����?��`�sO����a����{�`I��<��Y{����m�g3�0 ;I 	\E��It(,G���r��o~��R�ᰬ�� %1`� %�@$ ,��t�t��ךY�/>�����LJ$������[K.f����|���x<�go}���E�#c�{�ߧ�M�?DC�c gaH_>��(Z$�}]��Zv����$�(^�r�	ϩ��:Cn��6���iK� f:�S"���'h����:!0�Z��˕T�'b�� u�A@�pؗ��^o�w���f4>9�����mJݹ�-�B���hm��<� .�*k. [@��?A린�T1�O�8� A-��^n�o�B�JJ���4��#�08�D1�DI�mQ������D�*�$ۖ��p��'���f�o�꼂 ��dj�>�F' ��$A		J��#�5��!J��F�t�D@�q1ME~�@6�R�:PY��P�W:\���Q�s�|��e��3��`Q1|��G���8~���o���`�zc8F$r>�ϼ���h���2;Ӝ��K4�;��A�L\�83�e�mh:'an]��	^^Bi!5]Mp!���IH�d�
u\�3%+@�(�A�x �\~|���N4�����-�e-�'�Mı|:�u�����Z5O`;]��9�YR�;|�"��b>�,mh�ݥ+�}���K�ݤQ��QRced8-�t��\ ��7��M��>����h-1�}kд��C8t��L���ϿMf���a?�
���T��J͈ �ǒ;]E���#�ێHW��ze<�PgR��C��,��T"�dJ	�"l��F����M�@�1zpt�A|���[-򃎀��<�i�4Z��Ɩt��\W�h%�ɷy[�q�FsxM0��d2-	�Ȧ�.���BY�t���xPq���8�$YEyaQ�T�@���Q������Fܥ�YJ_�U�=��#��oPe�{6�n��;g ��ʢ�1��Ќ�[��\�t	���g"�0���?��5�����`{e�Rbl�3L��`C�a8��h����uL���-I��ia�52(R�YjV\O�C^U��</������Ƴ{�������_�s�ŭ~����+��	]y�x���M�Ƥ,��hg� ���6�H3, �Hu
��?8���;``3gP>�&U��@3�,Ҝ�Og0�<B���A���\u�)VanK)��'\�l6��bD�G�Z|^�Crmd&�(�@ȵ�j̳�� �TAM�%Ci�bG�a*�&��\���1��]�P��6���z��]QOΩHk���7$�d�x���>�Sz�UZ���X���X���������8��,�>���'j��vl�)�"x)$岑N2��p�F��3(J-\��0�{B��di��!��RQ-D���VA���d�n0�Ee)]�&�}^���M�A@F�g���� � �+����T���i�u�a���F���dΏ��IN.���Ma�8� �1�A�������Ĉ�%!�IGV��(f$5[,�_�pJ��ik`S��\�ҡ���� ��̋��]B	���K�^��oʀ�b4@��B!��|��5r�_�]uaբ5� ���e��)��;�'��n�6���u�R�jx��	_hK7,�yBG!��q<G��0	>e����N��5��G�X���<~}����>?�����7�hooo�7u��l�k��9��:�b3D�"�_HY�hkW"�橴�)=V�ȹ��S{8���GyK�3��Y��=��*�y�>����`{.9-W �+��%]x�9�.�sszvA:���DF�B$
H����k�
����U�Y�2Sds���KXT��˞��C���BI>r�����u:4�~;��.�޽{tqvB����>��z�����=ƴ�ױM�?�AЂAɗ\�z)��_,�_��_-���c��2]���J�&I��F��DI5�2��R�&ب�u-��*�	����U[uu��Ҕ�"�������+ I���[/�R
�T�Ŝ��]jw<�81�vm � %Ġ�[�l��IPH����-ߥ����xJgSɐA�i�%����r!1Uq��cO�V�^&��V~����EW���X�b`��
��6�S�nT��ܑ� "�'!��snks �`��E�����Xh{ؓ�-��;̚.�X`$�+�3H� �����3���Xּ^s�B�����5E��fp���1`4�]�u��^�!�#�v����=�|l�]�x6�nN���^��æW�G?��l�2��廧���'��$���)�lw��'d��(��{%)27�PFS��4�^�+=%�T��	��BP_@CyҽYAɝ�rlit0���N�*��S\�yJ%�N,�Ђ��d�j�����M�#jG���s��*�]Cu=*�T�g�τ_3E�S$?�E�tNu�E��F	�05���/�ѵ�]�O't��)���c7�~���y�?N�:?(c��c=~D�&�O��E�ڝN��+�&������e�=ϰlh�T����W(����P�X���0`,%8Х?0�@�xi��Tf	�i�e5�q � 0ji]�E��4�۷���$j�e��R	�H%@X!�t��T*�_��'��(�O�1ER�����E�7{��i��o������E�`�P��2���3|��.��lP�G2*��?82!�U��3����H(W�[�(%�h��e���������7	�tҁ��<۵�,-��YڒqK���Ab��O�ov���4\�x���+3t:Z�-���m,[uvY�qb����/Y��4T��]���i5u}����"
�!�M��W>��7�`�o��7G�����������/_D�Ǧi��)EA�'e4dgɂ">G�$_@��H�p��Ob��:)2��nB�g}Hn2���!�D"&ώ�����:O(�A\2�]����o'����耬����o���r5���k1���"�ˆO(,W���w���n=u�e��5je��	Б�����\�D��&��;�޸�l�������>�5hZ���0���z��l���<��$�?^��{�R>�m�r��L��`Ϻ��a*�Fh8�y�H��P��R���2?�$bp��BVi�ㅿM�E�	|d�@�w��'<�v��&R9���%�K�GB�@��� ���.� M����� [ڴZ�/�tZe�3Hs���v�-m�F���)-8��q.�&pSv���ȇE��M.�Y(z�l5�$2
������r(���vJ��kA�<�9M
�J���$�xUR\��֦1��;2�k�5bdF)Nҁ�[|�
M�x��[=jj��d��e؂窱�$opeJK���X�j� ��dᎩL���;�Љ�l8Ou>���`z�w������+6.�� ̮�<:��q\lNc�A@���d��4o�[���TF�]��C��5�/Ǽ�K�F�D��hS��R4�RF��"����ūQz[�6�n���/�4]h� e�Si�(7����oĪG��ie���?�dJ'@wCj���b�҈���f�l���8_ϕ�V��|�����x��_�u��q�5�4�Uc-9�}kд��#<4x�u�4��s:��(�~)N���*�ǚ*�E�]I�Dg T�2<�v������NkI� F�/�L�V���W��/�r�y�yB��;��\� ��I(O-�}j9"�,Y��s���6moMӂ��t�M�A$�#�^�'�������A�C�W	�B�9L� �TuJm�P0�Ei&5jGH� m���R�R�*d-���'���M㉀��nV�$;�$x#HC�@:��	�=�X���gp+��hwO����84�(OBzp��5-���H�Y�9���fc�^�,�	��st�"W`�68��`S�V�V��c�NS�I�7��D6å�g���c��_�$��h���0zf��V�������}��C�!�tjJ9x�譇�w���<A��a$2�)�ʛ��ǭ��Rg�R�@���*�(�$�� T2����xL�(�t6���	�Lu�)�_K¨�y�`@�	�M�n&�Mz҃g��l)U7���e��g�
�U�V�e#�ѥ�Z��Ё�3p� �d0K3����qs�?�'ݏ�O/��+��r{;���kд��c0.���]���ɿ����Ӭ�Y�n?U�N���a�T�b)n��R�h4)W[:Ԇ�L,��Rsr*�9�ܒ8cPRpB�N:t���K&Y.�2U�u�D��ZJ_�`U�
jh�Gpw�Z���;&u��n�֦C�8���f�P��x�9D&Ƣ"�Ds	�%0����o�T!n�����=W۷ɬ��]-m��aQ�7ȪT�f�RT<є9��VrE&��e�������M��Q��Xp@c	�T�^�-�6�b3���Hr:�%d�2x�����L����}�l��X,b
Gcr8��z�@�G ��R��<Mi����
zU�QX)�(��/���%FЮc��=7͓��b��Q�~0_��Z����{���ʕ�ӿL���p�s�>�ŋ��9N�KAC��t� e�̉sH�L��@+�a�.E��05R�T ��"8�L?JJ:�[0��[�.?&DY,����e�|��<�Q���Jɒ6o2�U�m��Z:%���h<�V0����Zi�����wl�:��)�l���LY)�Y���d��U��8�\S�d3܎��'߈�g����o?�/6w������Kvsc��c=~��V�xz}<�~��"�̟���mEM�|'�����Ȉ~!cÀ�g�Cb��p�Z�eǝ�΢��T]r'''�:=%�	Є2ײ$�������0��96VR�hDż �]'hB(�L�0@ɰSQW�������b���90n�i1����H�z�l�'Q!�@և�o��vz���S*�4� J��˴|���V5b��J�x�vuD|(5K�������3�x��(G����2D)Ҁ�9�窬��t��a�@�`}��)���2m��F&����֠��T\(P6ˠ�iS:17P7��5V#��_�9���+x>�%<'�%�h�c��mf�]��i��$������(:���h������_t��yg��;�w�>�x�()��p�{r!��R��B�J��*���Z���F͛��͑K]6�D��5-R�i�^@]�!��S�� ���'�,zcPo�\!���e�D0�Zs����X�Hg�Ѩ���U����|ɯE���b���7APU|
a�S�f̯jT%=[DP�>�l>� ��h�1f añ̓4M���w�q:�g�d���;��u��X���X���T�{���ۣ�>���������Piԛ�c;��2% #����TxF��3�(�\�i��)�2 ��ζ��`	6��h?�w��Q/�I�7T�A�.�M;[;�Zb^2t���� �&�e�����\�Hf!h[����:��ȭ&�2.��]|mK�1����Zh׏���YC^�G��'���	���A��./;��"Z�mU4��'�jP�j!ڣ���u5�
���7�)� ��b�+�Bi�P:�T5<_��|ۡ��m*����<�mA6��N�)�M�,��0"�����G��G ]Ϧ[H.P��2ϚK��䘸�@�:�|	9	Ki`�/[��׺.&XЪ���E<�.���lv����ύ�{������������u������k����$k.E�I��`��o�fbr9���B�-в���
�2=*O���F/�� ��W�x�--nPF�ku��0i�O�|J5<��J>΃~��_& k��4"�4�0K���XJƵ��C9��5�� ���p�pb@�A�~E��@���p٠��xQ�WB�(��k�/�q��\Adtќ��5�n�����~�[O���_���O?�z���5hZ���1<�������t1-���gD|���[m�4�ű�0�����,)nR]��?<!;�W>v�.m�P9!)[���d)�h�D6�R�-�iBP�=�GX.2KJ�Y�n#��}
Ð�ڤ.�Q#��y{Jej]��)IY���/1%� [�� �i����>���|j�\�:}�ˏ(��:�E�A���r�TDx�8���ޑ�\#� ?�D뉤�-��բ��#����� -��Ȁ���n�G�=�rP��Ō�G#�Z0X:c�h��Z�8&�YB��
8�q��q�C1�H��y�H����ө��~�3�%${GHIx���_[��89hɶI� �]���F��w�qx��|�����?���}��e">�?�����?�d~������OIV��7d�\tr0I�W�����H����b��)�l-�LM����h�����mG����Y�.��-M� ����U�Y��!�A�|�%C�$%��c�4h�iB�m�i�U����>�*&
8�K�
q_$<�h�:W5H���]���!]��������nY�>O������gkk�˗/��d񿞱M��AZ��T_8<��N���q�}�/�����u�������R�'P�*�SM�hy����,-���A�	��K�8�2S�6���v���x�plP� ��s= 4��R���Nۗ6sd�~�o����"�Hh��H"� �;�*�J�r���t2a�����z=��ܠ�A��^�AE���j�P���8(BE��}�Y�%@�B�G��g��Φ�iJ��ʷ)��-���cx��6���N8���|�#���..m��4�&�B:<ӄ���հ�a e���>a>�ʘ��L@=����6�o�"%���D�ܛ��5�0��(�V�||��Pd�pl{�@�1a�v1X�r��Z&�a����(2|����_�c_��w��������If^o@Q��8�\@��P�Ķ�̭�G4�4��F�yt��L��Q漵��Q$lp��lA�g��k�� �q _g�A/M�G��Q@�~IvN5�)��ʘ*:ʷB��C4���MJژkS��$ &�?,ǖl�j����nT:U(�ʩG������>��J��cI������h4��x<��ggg_���>_�����M���C�#�sz�Qn��Q�8K����TW]B�Q�%x{)���2�J��(�"�WW�RNhZv�!\����u��v���\U�"�)\����*l���$�e���8����3��a����	��p�,�PQV0��`�T�4�ہ�b���`���G4�ЌIZ��m4�G4cz��ou۴�oӠ����ÊE�)[D���}�Y8LX��Zʌ�j�1Ed"ޟ�����g��%M��IFֆˁ|@�oJd^��^�DJs��`�E;��HLg:��A�xJ ��a��%�	��R��Y�6#Ǥ��f��hQ��g.`	/�<7-��@)�T�<������y^ �)�As����x1�|���.ϫ/�x�/�~�<5��a�6�a���(��\J� ��˵��`�F)�c��.u) Q�ƺf	,H������Ju����^*D��CG�����ł:pd4UIy��b�Q��ejTyP|���F�H�O��d�F��d<j�Dƪ��l�xmC	�6�R�@��ƪ�Nm�IK#glL%|-�	��5?M��C�/76 �=��۷������wv6~����Ϸםv��c��c=��{M$=�����i6�7y�������U�apV�2�@'��N��Ɲ/Jn|�Q�J�U�� ��X;�Z�u!l�3KJ�Ȕ.. �RL�3)w�j2������=�� h��>��L�@g<��%
Z�MN���N2͕
z%�0�E�I�*3)����b�Ԏ��(�)ͦc�� C���i0� �ף�l�D6y�J*cb����/Y�&��8�i6O���X�A I���3���d��Od ��An�1�S8C���|˥�ݭ=�9���>_�<Mi� ������Jg"�V��A!���,�u0h`P��r|�}(��J"��(cVj����nT��	�:����m�q�(�J�6��̦�ܾ}�>�����G?���߾�����G���jS'�q�1��%���h)C�KY�e����B�6,���@Cuƒ�dHV	���b!Ә��d� ��|�����7 Ȟ1X׈lw�[P����+J���|֍Z�VF��\'�e����'Y#�PUi�����/�v��R��"�
�aK�#C���K�o�Ѻh����,�]O#�,�p]����#i��w��>tvv��^�ֿx������c��c=��?9�ό/�_;���`켨��k�llU�h�_�2��X(���@��n����K;;�Z��Qdld��G�M	I�Jq��@S��jz�3A˥�x��>]�h�Ӷ� ʍ"��c�AY��kd�@�ɰi+��s���d�-��%�?��Z9(�p����|��d6��3�����mQ�ߑ�a��= xǡ�h0`���d�`n� �mϡ>2?�I[�=^N�`�I ض���"��<wx_{�}���bJ�"�0.(��Sr�.������E�vEY{4;�R��xDQJv���_�T�,;8N��"�eE���]�����C�l�is���!Dd��My?F��1{�\ɖlm��iL���W���U^�~��O�;�h�V��������<^�.S�`T�+�X� ˃� ������j����C�F'yS�JW	���U+%Fʯ�<��X��&T�v�Gg�\��!x3j�%2GK,�l�j�ӂ�z���d5�Mt%�6��<K����8���|U�DJvˬ���jl3:.M%�������Zʀ�>��˗j�u&�^���v��L��[��}������ܹ�|>�y���3Z���X���X���OxgD�qD�gޟ�'ʢ���8RV)�AըV�%��Hy��\:�p��ؤ��-�j����@�-�Y��L�(a@�Q|�j������m�*�f��¤h�� W �wdFP����N%J��b�TU])��M�v����4e��o Z4�2b�%]f�61�g%�sGd1�@F���tL'����X�a+`�(͞ǯ^��A_��3(�Vx�R��F��${Q+���Z�7;=�v�ÅhR����f�K�f�����е�C����AԜ�� .���q�P��ڿ���b~��s�������S���	A ϭ�Χ��1y�!u�qKL$������_6N_�x�+/��+'�� �}���ۖrd&�����2���ڐl"2�Z6[ ɒ?$����0������J�ےҚ"��ݏ�Ԓ�:��o3(K��'��|����k�8:�)�&�T�1�l�ТTfI��:�d�:��5Ow!����g
-=�ձ�ֈ0�e=�V��"����EG���Q�e) ɀ͏��*1��䷈29�Yd����Ͽ/���~vss��ݻ��+W����N��c��c=��{�Z-�vGa��$.?V��3e^=ZT��8l��Y�?V���h�O�X �t�9���v� ZK|q�n�#$�q��=�y(dlC�i
�s�¯5�������A����@`��-b$*��d1��� ,��Ȓd)߀3�#�E�F��� "����ox4�U�n�A�M�G�h�����9��k�zM�6���A�A^z�>-�/^�<Τ��(��%��6���{;��lڼ��iL���W��B�����b0mLS��^�:AK�Y��tN�鉐��%�Pu�E��nѣW�(a�9[��](a� �a#Fz�R���i`���)��EJ^���T��{%X�v�6i>��I8����п�5����O����%��U���x�:�L	F��Z�vV�(8�u�APʥ���@�Y�D3���P��f��/
K�آT�Q�,N�t1�P5�Q���]t�A��>��k����\*Y��&�Ç:h$�ʐ2^CKG����<2T�������bOy7֔h�p�{(�Z�2Y�4T�T���>?�Tj�dg3�0�ߊ�;�v�H?q~~���d�G�������/驧��z��c��c=�c5�"��� I��E��,-~1-ʷ�Y�o8��paԺ�9�f�ܠI��&ߓ��h$Y ��?�t�P��p���*h0!�Uj۴���|����ї�:t�� W8'�,�O�MЊb��,Ռ"��p�)^v��~]����W���]�ǀ�Fօ�?�S����4�ɲZ����������������� �5���� ��t��#�i��g@6<%r׏_M�*S�Z��R�,Y;��1o�!m���C��b�QI�!�ȯ{��[B�>�y�f�NFs:]PeB6a �B��]2�l�;]�JJ�x�f��Eq(v5Ý���&��?J�a���Ǣ����]���sxܜ_����������Z��O��7�49�ʙ](t��a��߸J$�2��@ �RpzD5[����@0ţ�� $��6/�F8��TNs�Č��	��� 2�\���=>6 ��d�?�%����� A��XJ@�qh�^¿�Uk���V�.�%i�J�]�𦤬����/���u� 4i)� <?�,�+`9�ضZ�y��:��Q�@�d%�2 �{�7�w�0���7��x<�%����W�����?��ۻ����M��!%8��Q�$)������"�ҞR�E>��F	�XZ���e8P���r7@߽����Ζ��#���IДvi�kr6�� K fK����z2$��k���"/� Ä��Ԙ�G M���6mmnӝ{���+���ɉ,����q��PQ���4`�TE�.��踸K�����}�"�iI�a[�k��*S�p�/�"�P��61P;�mM+��WN�j�#���T6t�@�_\��n���yх�nC̍�XȔ$�E+��'H�ؾJwQ�VC�.k�0H�yy��,�))�\��8�m�$s�@��׏��V'�h�'�?�_�lGt�@�����ω̿�4���"�ʧ�y���'>�������ѿ��O�;?��Y3�B&�B��Z��D$�$1�c\�!���貗|�P{��F�e���E-F;ci1:��t ���������LtC�;r�F��A%)Y'%!�rT�D8G�J�/j�[Q2�-��wF�0��Rۼ,�=�a\z8*�C󢖬&�2E�I�.빚#�,[��|ڮ)�7ۊs`e�RI���h�8O)D���Z�c�Ԛ�m��w����7�x�|���\�z��G�B��c��c=~�G�X�[�,{���dy�ɬ�����q}v]_GR�0�
�Ԗi/9���{�bPs�� ���S����ّ��C�g���f9 / ����Zݱ���l������^]+� @�P�;Cy�"<��L8>�N��x�:�]����Э;oD�/]}T��r�7��2���4r`��ѕ���k����dJq4�[�"1A�C�n�����T�e4��z�)%� ��9q.ī����������M�d �i�x�=�r�K��E3:��ͧm�T�ʣϵ=��>~��I02e��%�&Uf�����C;��^�wLc��ZY|8*� W� (�/��R�T^i ;������LQ1������f�)bO<�������������Ջ����?6�.�����V1x,�X�jڼ�$mW�dBc�1E=[i �R�C֤!e�[k)dZ����}p���gg�m����oS/��gss �L�4�]P��F�nJY��)pQ+=��^uY
t�2�<F�t�z4��>K�"��R�{��<�U,+]��r�Js�Y.F2]��DK�eR��F� ���ﲆO �m������}C&TJ;��c
�_�)뗼�W�l+�'�s{��_9>>��}�ʕ��c5֠i=���lh��i�;������y^�����u]Kﴺ���]��� �,�Uf(-r��w@���N��t*޽�=�� ��
�Q*� W�⿗d�f��Mゎ�R�ۗ,��A��$���;����LXO�Q�@�b<'�A��+�Rg�կ}����i2�����47���KY���K�	ݼyH�A�.����Ɛ*���"B���%�n��h.当�3j�;v6y]u;]�B�R�t�y��6 �7�Y��Ԅ�� �Z����B���-������v��I"Jf#�|
'3��9�|O<�(�8�2���?����^+�qױ�C���,��0��C���(I�Bm}�ߢr�����)%��w-M*�z]��N���r��eV�	��tͲ4��9�����u������-˼� ��71��s��-�.��mm�R]e4ŢG�N��A)r㳅 �>��Y����)Ut�,� =ؤ�z�p���S4�����'1���ލ�4M%n)�ָG�YӎDn@q�D��PM�����)`T�*��:�����J礥�p�`�T���VA�֜/��U�)R{�*~�ڟF�ʺ�P�V�̓��st�j?E���f���l6�����~�5Z��X���X���T'�0)����'˦��<ϟ� �[����@M����k��(��Sy/is��$8�� V���� ?�Zr�DVf�{MG�"O$@�Z*j%M�����V�r C*Ӱ&�=��I�S��QRD�]c���E/��:�|�6ݽw��T���\Э��ʵk����G~Х��-�3�s��iH׮^�aw��jJ|�-
�W"u1�08Ki|1�����u7z4��S����*x�"	> v}�|��Ŕ.�܎C��Q� k>̈́7x��ۢ�~��[�(ة)'OǴ�C)u"0��qG�l1�@)�;��FqiJU:���h�2��S�6&%�F���"1?�8>�Hda�<�-��	���J�CL�.ZD����͈Jz���/�����x��oy��W>-�K�je�`�8l�ÐLݽ�Y��C��w��`.����JQ@�%p��u�3^V&��dN�c^@������R����(�{�g���m�E�E"�H��E�@!7R�o�|�ꖓ�{��tYn�^��=)�iФ�ג�-�#T��<�c�7��K#�K5=l$��A��`��'>�_�t��4� �i�� �z�����j�����m�����`�o��Bk��c��c=~�����YZ>]��O�e�3M]��2����V�����@	C�4�%��;�s	#t�moo+{���2 ��})�aT�C ��UFc���?Bs��I�9�!seh�@�2Vw�(����Q� &�4��l,m�A�O=��v�n�;�4�i��M�4./�A�ɺ����ms��nH�#�Ft��}2����9A�u<��ڦ��!���#�N�i��t����<�=<):S�9Ǫ����az丁��' ������8��ӳoy��vv���"��&���X$��~����[|%��W2O�~�v�����Z��;o�k�ߢ+���7��V�a�PXe�Pb��H��	X"�f�IJ'�g��ܤK��ҡ� �e{4�F�W���G���k�|����`L�C�,G�W@�ֶ�30F��!
��ʤE���}�O8U��)� �:�� ��sS񱘈�2�ܖ�&K���EE�����)��9�ZyJqN���ry�SRzJ��
T���c�s��PJl.�KJ<�X�$�,=�[��h�����6�qLd�%�����P-Dyk%�i�ˑA*q�$�Ehj�:��4*ɍ��$�
Uj��Iʞ8�x�{��;���5hZ���|�sӔ��I��*����٦���h�E�T|K�hS}#��'Zh���Lf�nw�ҥ�j�a8g������޾�mP��0�m*%܈� �t�i�7Z���Z�`"�##��(�k�o�l�@�g�| M��6��.��J���������{@�i"�dh���b���{{gG��x@�F&)���_0��J� T�om�iw�2���%��5��4]:�)�����}��gGdy>=��3��SOR;���|�R��}H��:��tNaV�9p^���e0�h4Lx����w6ɫڢ�=�i�e�)�6��@��4�2W����[��ֆ�ᨬj�\q��4��/Dgj�צ.��JE ���4hݷ�X��2F�J��,�`��<��hN�`� ����v�|�����<��>�u&�H�4e!`�@�!�d@�xb��ve8v�y��D�@��o�.�JR-��Er8��|���bXߌ.�CDiSʈ��\&rހ���ڍ"f�[mQo���2M��L�Y{(�I+[CK2-��K� �0h�_�xQ
�[+%V5+2y��'�0���O�<�p%��g�`&2ê0��o�" 
��*��:��,�Sz�M�m�̶��B�O��>��AJE�׃֠i=��Gjh�Rk��7�Y�<+>YT�;�"�)�]沼`�];�%;Q��dHj	2]�z] .�GGG�uAyhwwWu�Y����\|�N��fE.�\���Z^KT�і_خj}��]�+�H������J%\��Ca;��*M�e�sߵ��[������ |��W�)�;e�-�/��M�iɭ��UF��ǂFt6�h<9c0ԦA�-v�d��]��.��֞d-F�s�^��@�[���E�i��?ා��/�D_�uz����]�>K7�N3������&�}��9�x��M��6v�������F�D���ag r��Ѡ�M������	�����S�� O�TU@8ViQ˜�k������w=CW.�r Y<�5#2*�O��%��i�"�	�X�돿��ؐm��C#d(��YIM��rq�Y��Ǫ���� ������varG��a�U$��w�����M*+ShEIK1�	�^>:[�A�l,�"&�w���*^n �w�XdP,j����d�@�0M�7�}��\y*.��0����ѭ�S�n�jP�&+�|��\=M��~Q`H_��N��2�8w!GU��xJ6g�V�g��"�լ���玲�����+ ����q&Zy:��9�~S;��kд��#2���Z���>Z����]�iʪ��J��;MC�j� lP�XZ��{�O;��4���޽{©���5�J�j�
�ԢS	��J_�C$C%1�*aG�oK�@�|I#�Z�@�(�*S��fs����/������������[�^���3�/�}��[Ee��05`+�Lo��c�^����SC�ݦ�����Kc)7���@q�Ӣ0�I�v�ƍG���78��)�G&[b����;���v�św��n��߾C��\=y��q倮��
8���n@��%��˛���|:���5��K�W)0�?�@$LT	
Z?(�L�v:����h2%�?I��/��1Z,�1�C������������m�J���UY	�8D|���ƹdk��� &[�����B���>9;g0�(����Mϖ�#1ܜ��?x7�[�?�)�'���w�m�=BI��c>u�RzqBn�'s������|�ng���ߡ��8�<g��Tۑq�6@��lJU�"M��e(^OA�HV	��DY����&R �T�f�F4���|'S���]RUg^�Y��u$m<�U�G��0ߦ��Л����4�[55��O
�J�A�˙Z�
LA�R�� A%4��\��N��e��J��C8�DYJ�x����;�4��z��l�(9���U�?ǁ�)�l!�(m�|1��A%�8������tFA�-U�>�c76(�z��4,�tv��5��R AǪ"6 ����,"�����uby(M��JHe�\K�eۉV.��dWH�et��Ѽ�׏�������������y{��ml����8�Eѻ��c��q5g O�\�N��� h2Wv$U�
��}x���L�����I"��U��g�y��^�D��\.�<���s��zt����Kn������c���})e~�k��F�MO0�zǳo����L�9^݂�
�����!����-�YE�Oj�KC�� ��	r���),,*���z�!��&��1�{"ƽR.��(�%E���5��'��[��H�Q�E����tO�k���H���\���Kbɂ��Q�1�����b��V�&-�����X����6�C������+d�~�|\����	/�JR����fz��`���P�;���1ų	�"1P*�t�$�t���.�%j�]Y��@M�t�MpO-�%f�� �eYNI���)S-uUL3�s� �!'����.3Q���w�t��k
8���E~+���ZDJJ|zY��C[>��U�.�C�.+�
4�T��#̛5��]}���7����?�����M�?�@)&������q�eQ�/�7˱M�6$�	�Ȣ$��������5a\0��i���<2I����K�"=ׯ^�I�Ӓ@�Í^�T[{G*���x���Z-(=+P���MQ�W�j-Xʃ�bԝ|�.�p>�����N����^�3W���𶆆��[���>�b��apv6�/�k�I��y����gn�hS-H:וm(�y��LA�FKt�
��jd<
U�ʒ��Y!��}�t����=�N!��Ŕ?3���ѣ���p���\Ы���K/�B����X`p�����;򝚼*(h
5C_�Xϩi5��\X<:CV�fDC�ݒV�ۧS:<�0�h���Snk�ܠ$�^�!M)G4�b"��%f%j�5/��fdUl^�������<�)f��j�i����i�1Vv4�h!�)����D�*Q)�����?&�������_�L�����c	�8&�ш�](!'�,q��@��o	��AS��9���	��k,x��^��F��K�5��*�S�m[�4�e/ Sվ4����2�54q�)eq :��hK���]q��R�m�C]'M|o����;z(V�h �z��g�ȘQ�=�����Wz�4	�b8�����w�5hZ���!(��E�$#���y���2�4�}�7=�V����Vk�>jG	�IJ.�\�`{p&�yD/���9P��|�����=y����� 8�۔��)"/��.�@�,P`0Rw��,�T�ZҀ�O�����f�I���7�������<�v�ҥ�/37O��)_m����s�n�a�3iQ>W��yݗ�� �]��OE�ρ����L]+�_���@���;(U&4������OD��O���|�q::>���#�9yA�.ic�GW����|���?�����v����.��إ�]3p����5	���!W O�b��{TC�!WV#��a�T����Ӄ�1�;qf`f*�Q�Xb�m��|�s����� ��C�c23��"���-�R8�7^� e�Jt�x�	��������"��"a�T(˜��Q���T���פ�@���&�;;�>M�N��%���X�q(�����9'���KU�0�И�ʪ��@�ȃ��� IcC-�O��=�.9C�LE��"9��YZ��lM�6�#�$�h�nU�,�J��r�$.�5�	XZ�P������UU:��������K��2�	3���U/}���h���ZL� D4M͟������T/=������׋�v�EZ��kд��C0,������_L��|�{�i:��6C7K�FHԨ�[TU�P�K8h�w!;��C��
����{|�~.�ɏ߸!\&d�p���7���r!p(a��mskK��L�p����mX�a-��D2�Ix���ȑI�r���<��X�r�w��o}���{d��R�9��F��899yi��N�O������s�z*��P�pW��� �I�RjMFw����;���헾�5z���裏��m����g��tz��s��y�[���-��'���:&e��8�E��{#zp��l�M��xB�̀[2�JJ��t���)�qB3+�g����lJ��!���vO�B��L� P.Ϋ���̍��<�Ɍ�n��D��s���q(�����(\�bs�.��0d+J��Z��sNt~~N:�e�b	R����@>�Sv8�~�a�s7b�)�,T�z�yХXe� -GD�R*��,�}�D��Bi�!�yh7c*�$�TE9K �)2 ���l������[%Ė��2
̐�Tٟ�����7�����]y�4�h	zޔ2i)M`�J� ɲ��"�+5�FI ��M�����J�A��N	xB�]֥E/�:M������^�wD��]c��c=~@_��(���ҷ�O��;׏���	�e���=��OQ�V6���LYT(o��]�|�v66�<�wH��ߧi������Xٝ���7:�@�Ev
��w\jw:��iJ�,�L'��d��m���T	+�7HE��y��ir����u���}�`��ׯ��s���{{{~���y�w��E1�gYY�-J��0z��^QT~U��0������.��(�"�����Q�L��y�&Ә6��t�����;w��k3���'{@�����碷�@g	���Ǫ3�0*�_I�Ѷ\��2��m�A�%d�2�RCi�o��q�">��~@����9�����q����&]�&b����ȳ�D��^ۧ)3!�;>��lR�L�t�5��iy���%�D�>��mupWtz~�.����ʊ�X�|�m���|MF��|<��g��.bj1�3x� ���� S���3����X�m�*�IK D�CN�F�R7��&6*X�k:�d*`�2P��Y퐩�������+N��̇\&�)U
8�T���[>4fZ�Z�2V��Ւ(nh.���X5M(B{%��ekř�A�i���z�9���e���k>Ư2`����Ƃ���4��z��� ;RfQ�</?������d���ҙR�& 6�Q�)xJ��0z(��#h,����ݾu��޽+ZJ�N��y��eB0�8��Ñ��kf��h��� F�M�g�t+Lh�ƽ �+ۆR��vP&,H�I�& ��qKz����uۿݿ��ŧwv���yխ�H����8��l��-7�g�������x�Y�]ե��S�����4�$��ymɞa�5:;�(ߦ��]z���"�y~vʟ��B s��I��<�yBM��	d��%��g��?:�y8�;��4m:���z乖O P� \��AݞOO>���t���'3�Y 3��x��=�6z6��Y@�r�ز���p�L�t���$u0v̊�]٧-�^�U�|4��w�2�󩷵ǯ1д4�b;��R1~	��agH�ǔ�@����<H l�����y]C2@�>����L�*(�#ŋ	�"�*6,]TǗ�"5���Y�	ZR����Zi�`�ʢg�}��)�c���,ս��Z�nh%p��j�߫�ऩ��V�.aX5Ɗ{�VU?�$-��d��&���Y)Ry�&QJKn|���C'd���^�-�%I����_�t:�ZZ~�M�? K���$�H�V�V���86�9��QA��p��Ѥ֔v�w�P��m$�8B�zc{K�	IR�k�ޣ��I�h��������C�a�@i)! 0��u�&�%.��
�e�jCȦ�pL[9�M�|���L���[O�
���wf��g[������}鱃�㿍��~����s������~g�&�K��eU}�"s�����ײ���d�0o O��`c4���@�i�;�����:�t��lSN(	U�&L���xdT�t4[М��-5�MAG�3��S�����6��q��B��g`���r7ڻ�G�߸F�E�`w.%�����Aۓ�T<=a \P'����G�_��4�H-`��K�#o�"�8�2h2]� @���v�30c ���Kվ���~��%������_��K����W��	&���$���^�o�Df �s
\8�r�<�tb2�i��V���P��.��I��Qm���3R檵�0��,�"�k��1�%��-����gjr�)����)+�y��|�{
/��1�Y����L����3�k��(t�z:��<�\(�K�ْ�v	�0ޜ�#Zv�*ҺL��nM�����,�_0֠i=��oq4�y�c,�`�zO�U����M��u�~�� �!���%�Ɋk`F�����ם�=	��b���1����6xGמxD���]���h�Z8I $�(��}!��"MK��r��lh��4:�JOF�N��0���E<�����4{�/�������p��k׶�yY����/�O�p�����b�{�8|fL��\�ʻv��K��!�h#�Se�k�ՕC��->qw��la�?v��PHң������R�M�4j��K�ܼw�^:�O��ct�t2�}ڤ!��C��/^�ݍ��x�v������ZR��M|ܪ�.�W�(D��I�dU	�?�ݮ��֢�kS����1HC˾����6d�c����E������Oi�Q�$��� ���~����x�Э����F s##��g2�D��n�hE�xPGw(@�F�2�KIK���Q@¥ g�%��J�T�q�b�	8[�,��}��d�j�b��W��*�d>�@��W��! Q���y�$w��C�M�=bՕ��X+�&)Ñ.c6�.e�n:Sk-i&�Bt�ꚃ���Kam]�]����l���W����@$�x+�qx��΅_��Ϻ=�Onݺ��}���=֠i=��oa�m�����eE��u]=m�n��AP�����)e���`$�n%��nJ���41��bN|�b.�ؐ�|���,]W[�t�!K��~���o ,�%܄��q�E�_I���+��҆A�)K�&�a8���E۰?�����-��#�<���0T��	||�8�RoM�fi�EY}$/�g�޲˕�
aA���;pc��<��;�"�9=>>����v���{�����wНh�)����SF|\�пj(�K
����lS�͏�&�|Ҝ2 ���{T�?��J����
�� �����v�����^b�}r*��*`Д0()��=)<7xm{�I��7t�ԠA�K�(U׼�M�o�&�]�p�rp� "Z�d�B]B&�K�T�4�LQS�M%zS��+�a"\��#���m�$ :�p��`��,����(�n)���ܲ�O-;�V�p�k�U��JS�=�����a�U2�\�Z�c	��`�P
�KIR.t��7/S�ҷ���'�]%�m�W���A+�ehF�����0`/�d)��m9/�ւ�%X���oY�N:C��+U���.c�N��}0����1�y<����֟����:9�?�c��c=��~p���,��}>��Oږ��8v�i8�ėZ�?� eOB"Ĉ�Qw�ˇ����GE�Xh�`�Ν;��@�C���!]HI�[^��6E�΄/�g�# d<O����0%XaP
�JR�ڈ�(.9M��)��&˒���7�.�S�n���ݍWߡ�?C�aO�8l���Q�o�,oVc��uU_�*ӫ9z���c��,.�ޛ�6-�##t��5~ޢ��c��#r:�65��E�vh�צE�0��(��(a`z�2Z4�G�6�ҰO��/&��)�1	��^O�'�(d8�A��
L�S>.�6�\ؕ@$˦��)dPj�Pv��ܢ��6Og�&�����]~���@2F�^w@;�5�n��a"v�B}��{C����Φ�5A����J��U��/�M�dɞx��IUF��T
�  �R~#%<�˒�t�YƊn�┥_pP�[fP�t��-0)9�Ze}T��P��z�0�U�V��<��\f�c	�H�%�'e鲟��Q��G!����`Q�蠊.�»�E�a� |��9��f�CY����J��BVM���K �/,|p\+��R}=K�xvt��h:�������}x�P�?�c��c=�`i�eW�q�q����;��u�/���b��G�I��
��c%��r#G�Y�V���V�x4����,Ố X����}�U>� �1(��:
��pq���L�8�=AZ��R%��4�UY���R�X��*���ο	����׽�����0ߩ^1$W^幼}~����,�^$�GҼ�9>�O�U#�2˖s'Xyx<_��x��w{G��F����
3&�ա��z���9Ⱥt�lB��B��t�Β)m�-��ե�����,;����Uϛ�~L��� � ��\qAi�؍U�ǆB
��P�~J?���J���K'h`	C; ̸���i�^?_�n]��2ϹU�u	B 8Ө�Q�^ի�u��9y�������< ���>� I,�R�1-�Yqc�Dr�����}��j�>�ha�`)�4���.ωƔ�ѐ��F�E��"�C�tӉS���yt���Zh�\�^o*��΄��M6�0�)u��e���T�:���#��l���{�c�zSݰ��.�$�q( pݢ�͒���^pڠ�'-XR��Mz��*[�������;�p�_L�|�"��X-�C������P�_O_xj��T�"���b~٠�$y��L�,��:$'Xr �p�z��@����*J*�(���5�|�w�D�����ht�ƍ�������k�>v�z��h����>�8��?�D?��?�f�O���2
/7p�jH���"P���p0�F��1��Py^YX>���7�Нۛ�7Fzii���V��n��ض%`���a4�-S	W��3Ў���X��x����W]Օ�L��h��F�ǗƼ�1��u�<}�=��^l6��g�zЪo��m�w�������㽻?��h8~�w�S��W2'���#"0����ں ���]�}kC@���"�[st{w�ڽ����ש���tz�^�v���G��b�_յ�o.�( �H҃��9�ሿ�|DA�L�jE�����t$���t�z��OՒG�|�+�&1z'�����|��&�8���Ҭ��hQ2Ӡ;d���y?�t+��l�P�G�馔A�g�6y�l�&o���3��c~>�R"�@�h6z���(3�k�^���k��AmS�j�8�!���V�[��Z�5�|]��[ �"�sd�RNU�^��E�.+*��I>�qrT�I��r�d��BXR�)K�M�S�G�D�#'`�	rm�$���GC�e���� �п�^�_oq���� FD�EG���Fa�b���J�E^��?�~G�����|�����3_Y__�u~HSv3�4��=l<�6Q���3�x6
�?�z�s���,����(����D6�$3D�H4����f����Ҋ94��ظ-������IV��9��9C��J ��3X�
��[t��Z�@BZd Ug~O�[�\%�/���8�%U'�y�	i�AR����P���j��bsn���5z���Y�^��~d��|�R)?���{�$}2��'�4?�l�T��^�+��yـѴ���J���3gh��O[�{4��m�ܢ�4ߨӍ�z���hgwWJ�窲�D����j5*A�Tcp��
��T=:���=dD1�nӁ+b�ؤ�nFs%�:�N�;C�N��hD%Υ,)�N�GWoܥ�7�js��0��N�H�DA�)N9o�

\�.����`F%����G�n�P"��y��{HO��T��*3h�S̷�S�
F�[���[|	b�F��r�&Um�����rI M �c���2 �2�S�  ��IDAT�61�5�H(�6���Q47�E�A����@��i�-��|r�BMS ������Ka��Zͧi?��3���"N��PEIoBB��x$��Z��lɑ��}�)GT�A �:�/��p��T_��U)�}$���?��u��N��ѝ��o�g{����c�@�l���`��I?����s*�%�;�"����Ɇ��fc���Ӣ�D��x��eqqY�J�1:&�����v��E�<iu�'%�RN*�p̅�yi[��o>eW�� ����j)���JUIǁ�$=���ABgO4�Ǯ�.��V���f�������[=���v��a��Y;\�t��Ϗ��^��.󆸎�Yf*�L�?1P%ˋԨ5D�`g�CI�Z�F�s�i�n��K�|�^[*Ӑ2��M
�s�����(����7"���^e`>�erk��yԫ5
ynlm�ҝ�;4��o��S�t��9:ub��5�3��2:HU��0b��[��� a�n�9� 02�������$C
�|i�25�� |���HáʫnXI���ѐ�"�l Q� ��Ӧ��mp+��L9H�I׹F^ "���Ij��c(�ɤjM��m�"1�-���qJm5M�3��3��6��Zv/�|�r5�E*�)��i���`��RVD�\m�kJRP�$��;F����1�T�q��P��se�Y矁��/8�oPYt;��ߗHe�^��/Z	1�B���_�ć�q�?ܽ}󱃽����/~��G��a�����٘��b���4�q|���3���8����؀�\��2[Qx� $��*a���DAR���x��&,,I?8�
Y�3Pڤ�w6%冈�@�k 1c��h=�V@�T˝9sF��liO84]���I�7D�@<���J���1���|����q4�ǣ��6��_h��Z���?�<pfeɖ8��΀�˛��U���]
.���|��N��<e^�gF��`�z]%��T8εFt��6��})���t�v�FnB��K�2�ڃ9�����n�r>fka��\��v���W=`@�	���l�:|:�v�I��.���٥�ׯ��ez��y:�4�*�L�t��:mm��5����!K��$���clHLt$v�5����P樤��Am��Z�	�;�5�T�U���)r�X�ؒ�R`&�)I��F'��d�P�+i<�_�$���^����d&��Jے<�\#���$�=�B�T>���gSq
�rIIZo�p�|#y���+j��K5�gR�r#� �)I�=y�F��^�F!"NU���)_CV�(A\�7�nȁ,�5E�m��j��/���� ;e��V#�\.��|f��?�=���^o���n��4ϩ���>�<M�1��@��ض�§����I�#ͳ���&8 ���褩�q�e���.!���0H��)�\|nN�.�:�q"���b���)c_YZ���ia" ,���le�,1�D �@�V�n̆U50|8lؔ�@7*��'ܪ82b���mk����+A�������ZǗ_}+U����������F�����?7���F���q��+M��$͂f�7;T;�GTc���@�-�s�.ݾ�I�.���.g��SwM$MY��G1ϵ�~H�x���l�7�j�'Q�F	@t8���F�Q�z���'�``� �d^�Ji�L��<�;4��Q��֍�i��u�[��y�����I��+�ߦ[��?d��|�$y�i�x�%�a�#���-2!���c���0l�;@���Fe�Fo\���r@I������ #��Eh��<*�䄯d��4��4
�H4�'�֥�= ��L�+K
���L�pl [����H�':i���r��dU�S[�GJ�N�P����Ǥ����H�U�.Z�@���ߑw��=9��xn r��F��
�����$:��K���Pbp�4*r�.�LH����,������6��b)L�s�'ůW	�s��
V���v{��n������?|��W�����4��l�=�a�m��N�Dӻ�<{*K���4]�\��чA�ީp���0�
�0�wmW�K?��ǎ��*���/`���qN�>�`��= #Tb�� K�d,�&��ɥ�5�@fe�K��(Jk\��p�
^�s0�H�y��%~/M�/V*���>s|�t����q~8	���8�8(W|���W�;�?��OD���a��#K���97q �Ftwk�j�����&X�ׯ^���'���i�A�-�h���s����^�C��X���n�*�!�,�xC�ȥS�.�J�D���F�,|HE �2D�:Ҫ��7�,� ����I��wQ1�����mz���頟Pꖩ>7OK�+�m�>�3��=O�T����� \H��#�
�#(���=�A@�v5N��x��m:��/ q�F2�u���h��DHؒ����4I�4UG�' 	 �����+3=�r��d��-���39��af�JP/�?��R�1���J"H�MoZݧLw���d���F���7��k_�P���H��R���`�|�%��#q� �U@�^� M�L'��;�߄j^Ñ�b���;i������e�O�t:������/<���h���82LD���ג~���~����>g�Y6K-7���Tr}x���|T�i~*)��%�r��f���@�+�m/���!����.�"��#=������+ؤYD��--�X�T�Y�vC9� �pk�&�{%�nA@��=I� ���g� � �o5�������t�v�ǜ�f�����ѧ�x^�����l���#�_�яg�/׫e/�Rg8�R�T��O>�0�I�q�z�]i-r��1��Ѝ�Eu�o3���ߔ��e�U��\[Z�G���q/q�C��m�}�GhyS_���>��I��JE4}B��������ep��+�hs�GC����%�uJ��� �]����BR�A����	-*��E >�{	}�x�cN
��
���=�T�e��\�!����(��I4W�,s�8S:P��p��5t��4�ᵙ�kq�C��R�Qb��8��Z�N}^Ҕ\f��<b��rI��#�r��h:��� 
�*|�����g�����K�nU"I��3Af �	|, "U W�x���;i+��c�Z{U.��Є>�@.�<C��}m����O��D����h�t����׾����Mz�ҥKcz��4��l�����S����(~[�%�,��l�]�s����R���dR����DJ�$R���Ʒ�p�F#����� (�%��9sJRu���L@��L�ʺ�H T�7����R�l���g�Q��#@��' &�a�t�9G�&�����F��0J�M���0ר|b}e�/z���,���F�`����ߺn��x��(���{�RP+߻;�ԨT�����X�ݸI��6���.�1X�ѿ;��-��3 R�)��U����������/|�ϜFv���|�L�:�I������G1 `���q�V�8�QZm��W^�k�7��c��o�ޠ�cǄ���+)'<�DIة�%�(�nS�L�LBWR� +���h:��7���=�-*���^!��avB�Ht�2%h{F0�C�6?=GU��QpL+�T���4��r\���%�2�*�ޚD�&�:/�P�p��p�l�9R�q���zO��W�R�Q�� �&�(t5:��ExL%i��`*/�gBjN$@���X���8���7���R�ZU'
�TԎ%�g�-�* ���� >�G��o�ݩT�
�����ϋ���^��˗/�xP�1g�i6~h���թ7>���}v��O�g���G|ǟ�M�츁(���[��UA��� *�,�����<#�~	��í���jg{OH�0H��:uB���B1ư��p Q%�%�5@���Tš�eh �*muR�Ԥ'<KM�<*������A����ˁ���|���Ź�W/_>���� �4������p�Q�O��S୒Wu���l�h�{ᡳT�ۣ�{��#jU�Щ&�/�P���t��]��Qq�*����Eä�}��';��ʵ���N��ǻ��S��ߙ��üٵ�ܲ�s��A�7�:��2��cz��jy�Tk4��9q��V���6�F�� .��k2Z8�d�b -��4U�����ͿW�-�<���>Uy����X֟��A��SU�F�1�-�hR�/Q!�4j�*���Q:���H���<�)��$d%����T�)�	���ܢ!�hS	�܂���8�4��ɤ}�l�l�h')p˥�N�ˡ]R���P��
�w�M5��^�F� ���v���U~ ���W����]�A�����F�F�C0��iI�v���0�Y-������e���^��Fq��n���_y��?��û�3�4?������l���8������<n�y������g4��M�#|����e����f0��s��e��*���~,�F���z7��KPߝkhwv�$��{�Mm)���s��qL�΃*r4����(�����$ewlM��+]��ew��%�P4�*�*yF�O��r���ɷ�Mb��y�"��G��?qj��'O�:� �[a�z����[��S����y���J��Z�����A��j�&�<}�����m@���Be�['$�0L��]!?�����|�J�@[+����y��v�1&�{��_J��Cn��������F�NPe��_m�+W^��w6)��!��z�) _t�r��Ry�ȋ4�CS[)��=	�X�n�k���U��F��ġ�ӽ4! �4�bI�K#Z�4�- S���"%F
�<+Di�؎�r����oZД)Iܳ	9��"�*>+p�9�HSn��FR�R��j<��Y>���{g�2%�$⤔!=_����@��u!9!B�&R��H��f���9J�W�mOHصz�!<�W�^��6��#���LlN8F�6�8�4��U�V������D+]���ϓomm�moo��_��_����o�?���g7M��]^(�?pzR����zni8�?����@�M��Q�Y��7���	3V��E�yQ?�?0��wF�Q���
Ȩ�i�xY)�I
d��Ԁ�0�h���!�anR�\��m��2e.��������,-//H$�ΓcZ4@�R��@~����gΞ���5CZ��+��w����_�K%�{»�z�<6�|��ᨿ��ٗ�����O���7g�o�a8O�q��|zp�k���T�^b7�2`�����|��iZ\^�+�� Tl�?�L�sK���ݧ�Wc�N�ܝo�kKT!��##H��z��\�ƫ7���x0|�0�B�%`���я�B۽!}�ŗ送yZj�À�ܥ�Ԝkэ�Mu   I��#(6H�4M89�F��iW$�n�	�;3t�0��рR����*� Τ��iQ�>s&FdSpEg�e�ܦ�(�'�=��kn&" �B���gC�\��cA�Myn��Q��1�$�]�� �:�f��F~���3�r�4�)�2�����[��L?��(��%�t����3����#c�ܽ���Ҟ�� 	r6햰�*�2�ch<-|%ߑ"O"ě�&m�-M߹d��K�u�c�b�8���_f�w�_s�����p�;s���+���C=��V�?3�4��������h4z�����������+��(R��2�����>�"?���U6�!�7�~��p�.������c�x�N6
?�:�S^���`)���V!�:$6dm�'���Ί��J��wV�T�Σkġд�Dy?���T�.}�T�{,�3^�>���7���j-�ӱc�h
�9Q�����}4�-U�}+rL�"�Ȓ
RJK�Q?���_iի�k�}�\>�9#w�y��J}c/��������8��,I�w��,��a7�y��l�S�^���ߤ~gHK�%�-7h���p��G��buo��3��O����|������Y���zcc�����T�ϤN�7��x�5�z�.��޸Ѣ�ĩ��;o�H��.�c�#�o_�$*�LFfD!�a�Z2�UR��S�&v�^W"�v���N�
O��,��t�E��0D -�xd{�9L�hXjT��9|h�8��h+)p�
Pf{�I�M�SZ-8���iqNB���y8��2aOLW9=�̨�J�a�)?�T�A�I��V�a���3�. �D�[$<�A8�Ƙ�N.�o�r�:�||�*M��g�ʥ��>f������ʈ��m�{�J%���E�ͳ|�\��q�D��,M����֏�k��c��{�n��֩S�~���v�@�l|���!ѱ�0��h�b�ď�I�����g����i߼��\��W���!)M/˝��A�kl������J������ΏGßq]�ggJA���%OR�rƱ&-#�M�[Xp� |0��H�`�.�	)8�JIE��e�\��ۥ^�/�o�--�(�hF��1�F�G�:�/��+�Tk6d��:t|z}t�'Kc��}�ꍈ��(ٻ?�R�����z����\�?/,־<W��<�C���AK���9��������q���y�v�`��cg�ߣj�I�9I=�F��ģ�\��Z�F���9��������z����vs��߸���.-ݞ~/ �;{�[��V4�ɩԨ����/\#��%^ \�'~���i�?���Qrh��Z%����T���ƉhIƵ(I9?��&���YT��F\���I�kyD�B��o���݀�ȡ�_Ab\[��Fy=���_�������f�����H�DAlS��5b�gqT5�2�e=%�Cm[$��ƺ���T ��x}�`� (���S!�KO:��s��h6���g�9iz?Ri�:SW�w^ɗh�Y�a<Rޙ_��^zI�jq\� 0�4��8!v��r4�$6�M��� ����/dp�7�k�F�`�@R��]�D�y�x����`�� �E�����N�ѳ�A��_y�?|��f�i6����?��a��~{��,�~���Ӽ�^Pvj�������/� ,w:�m�ʯو�y}���y�@��Z����,��Cy*���i8���(�&��~>Vr��y#U�x�5���nn��,����=�h.�̸q�9H%�v��t0�!�8�0�6Q$@FH�HH���S�/i%����C�ǉp�z�`7 $��{��ӕt�-i�\8��j4�=q���5�u
J�)�ˡ�%���Ȩ�Ԙ�]����U_��?C���2LC�M_��*Q+W�|���?~nǙ���räҶx~�O����0��W�!?�n+t�j�A'VQPb $=�k/�Ɇժ��Q�qb4�}�ƭ�������|�k=��G�3K�c��U^��/����|����/\{�n�uɫ�$���ﱴ�,�A�Kc�gDBȓ�%m�MJf���]F�I9Q��R���:� �o��u{{����^�28J�(������r�{
Z��6�N3c��ݟp�H�����c�c�}�-w9����4]F�j8�wLY�g�8#!VB`��4��!���x_	颢�ȅ0���<�ҁ��ԋ%RTչ�ݼ~S�L±ʋ~����jHQ�KT���BG���~���Ku~�ܲ~*�p Xq�V�N줡*�܂Ǒx������������O}�������/?���ofn�4��}��-�:z$I���i��Y�>����t�O@8/�ZG?�kds4rB~��Q+�O��ü��1Prlx7���e@�޼������`��Ȟ����\��z/5�7�mα���w:����DQ�>��.A����h�T&/p�5�6	a��`t"��X��L4I �m��Q-�|1.��j��|��y�(��4�Z�&��űV�)@��Uꣁ+�o
k��iqq���Bmw��C�r%bs}6|%�a���(3�}
�#���q4�˒��%?����§�Ǿ}���������D<�t�_���	�PP�a@�죃���e0�y�$����Q���eT�A�����B޵q�Γwn�|߱�����Jn�Y��ί�k��,/�V?�_�.`));�8��Ej�\%�s
y��T�CD1�VHye��-9ZI�K��+J�e�V'xR%DKT������^wepjR�C�*�ݐJ=M����!ۨ�;�6��PQJW�G�
���nґ�C>}����)�6��+Ҁ�iS��&:LFr�4�_�PwUS
Q�R����f��>W��
���D���W_}U��h��Pt�R�+=�ՈSC�\?_�e���2�bI�rM�s�E�F��� 4�ةF�]W���1���Y2��n��h�?��/~��ի_�x�b��h�f�i6�h>�s��$�~����gy��搓�F�Vc�Z-S���~5��j�����8N���q^0��-Kͳ	���0�x��s����$�����F_�)�� ��S�j�	O,��d�1�G�F���(�6������@hR�I��)U�Uq� �R��l�:��ϩ\q$k��k�(*���Oh�T�@�C��Lw�=�n�����=��V�-�!X�kȹ�Q.܃H�:BB��Rue�O��#�P��k*��p�I0m�f�j���ǎ�~e��t�ᇗ��,=pÀ��y���n��~�˥���ل�R3X!7/�7(�E�}J�W��A������`����͍'�_<y�tu����{��E�2=��U���C5�����r���p�B=�!��+����'��5W��L��x����(���&섇A��]uj��jrj�{�/�"�,^w�1���5�0� �n�ߟ)?;���!@u/p��xob̐�s�$��2�F�R��,R�� 4��I&��@����z-��w@3d�Ԩ��֭;t�fe�uT>�f�sGid�HH��\Iy��?�z%S��.�r&��p6�}��:�|�0&N~�!Ք����>'�������x�G�N��<�t�ҥ.���4͆�)�:y4��M���i�=
���n2�����Z���T�����/��G��=����}?3�(�����3�59�x�{�J�4K�؀<��n�/��>1ת~*���A�No���s�G<?8JF�Q���?!���b�u���p6�W�02�5ՎI(�\���+H��0&D�Tb@��b�PVO-)	 �#�U�	�%�%is��R��EBD�رc�����L��*�42������;�`8ql�[gڥ�ᐆ�^����>ù��5뿵�Z}����g��֜���@kH4w%�>6G�̋�C�[9��$Oĳ��� k�]�8��r$��18�O���>��h�Tu<��!=�5���g�V��Og/��j�F�;���d^�n&Z��NM9��rH*�R>���'"�*+DMp�9��zkA��f�78���h��B�	�'R��d�m2M~�n���� �SK"�O`�ht)���I��`�N�~^~���"���fR��L�*|��W�}e[�h��W��E���t���;�$�np(/��m��ÎX�X�O���64joRD��D�I"���9L�-��m�[�v�T�_��bJ��	�_����������^�m�Y�\�����n��/��K�������ӧ;o��4����ߟO�������<�����m�Ɣ��t�XX)Ru>/R�1�a��,�&^���M�m���~n�fޥr4N�i��j��,�k<m�q�����J�������o	�m)ח
��#*�(iTj�{�b׼�~$ ��G���6S��{�eKT(Q�_�%p�؃W� ��rJ���W����P�� �j���4�4b�(gNs�>$�;�7`���Σ� L��V���u�Q�����y�����l���Qu�����o�y�s�A�?Fi��㕚�����;�yO��*�:Uk�
��|m6�䗫n�6G�ܧ��o��r�U+���ҙsg���S��E��`�}���r�l�V��R�l���c����McZ�[��tR	�S��YW�����c�7�R��٩Q�� ���6����Pș<6*�~���*��'=�9޽���0M��!~Ք-����i8�D����sE^�dZ�8�r.�,��hZm�JF�5�ը5��������>	����;�2�بO&p�^����J$˶Ù��G��I�Q��
��z�)ϣ��W�W<dͅ`/�I���zOD��#{�?1?�n�}�֭[��]i7M?�b�QD�i��$M��3���,wr�c�&Z+�a�HLE���F�zLG�����k�1ZDڊ�L�%-���၂G9'Av� ���k���\���ܨz'�B� �'�ƞ
�rY��������C�i#; ����rvSف�Ύ����I�u���!@���B�\[[��h��Q�^�>Qx�p��sc>�0��KLsM"�[��� %{��Iǟ/��� ���<'��j������{�>��v%
���XYqz�v���۽9
�����Y�>��N�^SM0�Q���DU˵*��Z]\%�:O#���Ô^��C#�D	�rJ�h�hw{[9N2G�Уc��,`�%�S쏺��x�Q�6,$��y���ṁ��'1�l���J�*���0���l��H-��K��p� �G۪���F��L�-��Q����Dn&���t�����Ñ�>vʶ t T�A<R���;
哵-сC�mS�eJ.`���x�WHu��ͥ�i?ح�_�¶�#@
�-v�ES���l��kt��u����T��G�d˽A_�ڈ��0h��B�L[\(}	��;�B��6Ha��X�P%5p]2�A���N�{r0����|������w����3��C8�2�1�Ic�	^(�'��i��xz��03%��k{e�2��LtI\�)�Dd�̴��kx�N�<�˛�yA>��ˑ|:�i��:䛪��z���p)�KF�3"mF2m�ೡ��Z+	�!'��F���Z���KV���W>7Rh���D��9��%�Ʀ��_4��^���@#�*���l�m�,�Ch��<m�(bC�NaC¼�����.?�B�����b�/揭_}��c�L�{6������>������:��?�y���(��K�Z��2�@5���
s�AJ�����{��1�ʩ�s�©����J�i���؜�B`���3M��D<L�G�\Y���ng�J��T�<�GH�����Z�����/�@��M)p��G���4!{����4�۔����M�}'Q%����@���?aOF�!;V��@�T-Q��(��P6�����@�[�GF�a{{�^{�u�M�\;��lk��@�P�lf�	�9ov��h7Iɰ�Y0׶R�AN�l6ҕAO��Ԫ?��u�+���ֳM�UӮ*q^q?��c=s�n�o�~�}�~�w<}������0M?$#W����璈~���eI�O�*OrG�=!7��I��<�Z�,"���}�9�h�B�-���JCI�0��+�B����L���&�BrI��?�")3~��X��"���8�R=�R�]�&��j0�	ʁ�` `�%?�J�dUq� �&�>'Q�� D��U�hi�I���FAɤ��:�>uB�NLڍ�oB�#-P��7����?N�h���/T+�G�Z��?���(���7�⬨}����߃n����뗃ˮ���&8�"�k3�o����E��1��e�5ʴq�'k �_����DCYQU"���T�툏] I��!��
�bCw�\2�@n��y�3�ߚ�c����]{E��.�ƒ�˄(-G7i$)AD&O�7$t��Qs
�m�i�r�Z��8:�K��p��#��T�e�DGJEq]�F�Әz�����l�H�B�����3����4�u�^�:�h$^c�/��}�W8m�vlk�ޤ~�g4�ܢY��TR��ʱ���D�%��)�z�..��.:t�����HQ� ӶZ�^�ı��Qi��A��p��,��&�O��d�������~���|n0���իW�z���[��띁�|@�,�Zy�A�{x���'�|k�M����Φ�	�b2��.&��1��T������Ns,GJ_;Cy.�^��0 ���B�R���}����;%�.�J�2�fY"=�FE�ss[bݩx�r�oGy��`s�H��V©rw�`F�� �p��M6
UZY��r`�C��@�\�V��(T��V��e��#��f(g)�i<������皟�.����o��,��w3̼y�֭��ӻ/���_R���g����W*3����:����^��������������h�i�x :�N1�y���HH�Q�O���C1��f���&V!H����s�IJ;D0�<�?P�XHu�:���3�=��H����_��L~�~��c��~�M�ɰi�7��cyV*{ �3�Hwzpۗ������-*�FJ��*���#��m]G(�7��ܾ}������a$@GԿ�D����!�d*��|��Ơ<+��Z�b[3������v��}�[�	�qp� ��8*�z)C������	�UO�����R�k�7��,�3��v���t~������۷?q�ĉ���^�@�<xr�x�~�'�0�t�f'y��P�6J�zD���dJd�"N�WJT8dKjm'l*�:|�(��J�k񔗄�a͜	�Qº�S�h�u/$I�@,,̓z&��.�j��曒k4+Ԛ�j���STnD�-��E�T�y
�r¿2e��|�X�C* $o)��[j��Ғi�R�L4)p [�r�eÛ Ԍ�~��L�R���4�MyC
���;A�������_{�폟�sf|����S����Om���w��_���.��K^UERSק�~J��ݦQ�k�\���s��kk��O& k�Tg��w��M��I�$�.W���ة3R����ǆ�Y��*%���d�}��D�Zp�T�^"��er�<�
�h�q��S5VD,4�-TE27Oh7���
I�@9Z��J?�� "u�R�}:l��uou�ܷ'bFv��I���DE� �h⑈�TJ$��Kq�#D�5���'��u2U9ܓw�i��^{�6��i4[��F� ̬�+ZW�[�ȩf�i����4�?tPX\���{�Ν;C_����Kj����(���7�K�T9�<����8*C^|��<�c<���8��8=�������k׮}��>�hz O�*O�wFQ���"�ǋ�Է�,s���FS9��ҡǌ:,���(�I�8V��4`K֜���߄;��(:r���a�E*ᤴ@��K�����JH{um��T6W"EZ�QJ�8��g��8�esp�����BW"�U�j4��q�8�<(P�����G��$�+V!7��X���p0�T�u�p�����r5����<���}����{6޼���)/����n'��?��8M/�^�b'���]��t�G�8������/H$��FՆs$���=�@Ã}�=�Pw���z�~�8�J>U��Tơ?���j�1#��q��DX�J[8�pt�^���j6h��)%TiI�%��8	��1��{n4!o�]��7M~}�4!�H�!�OA-�=7egs�RוA�8�4&A��T�t���p�҂ɑ*:_����/
;��.�8T'Q���-��ʫ���A+���9��٘�0���W��[(`��&Dx�1�x񼜋��蟉���$+�?T�@���:S��3Ԇ�p�12���3�u6b��\����Ź�`���z�����K/}�߯�������\ s����v�'�y���,K��ZV�A	zf%O�R2mD�R3�1i'�4��>O�J��OE̟�Ǥ/H�Nf���M&%�9p�q$��s�N�R��Sċ��� ��Bx��Հ�֗�g�m�%�!��:K�ؒTXXH�p'��$%k��\q�4~���"B9�0G�V]�.�;2׈�T��k+��D	��@3��L����&��$I�f��j��zq��G��/_�<S��XZr����qg�[��.8岳�7��v�������S'��G�2L�a�e�E�F��G�~��8D�'5�5J���ͻ�[T���c��qO��)3<��Ylz�)�S��T�]�MZb�UB��	Ua�?-��4�8�*=���]r��������7�t�?"b�
�q�8Ӏ)+^bS�Fk	���	��P~�U��zƼ����B���JH%��q�b"�]i�h�v畗����]v2+4)�B�Lq�Yf�s{���'����V���&r�Ϟ=K�Ν��h(Zt��j���L9o2�י|�i*�c�T�bB��T^TIN�w��%uK������[[����^XX�����2e7MЀ� {��	���Bz�o۵��z����L�$�<�7ٛ����V_�E'� 6�ގg*��"R�g�[qܚ���+�Hl��+�h��t�2~��)c��j<O�w8�g����ñAZ%�y�]B�[��iI6.��{M*�1 O	a�J�< t)�k�H$z�G>��]SQ�m� �����C�8�ܱ[�Kߨ�+_\Y��|����O�����l� G����بG<�olo�ޠG���;����	:��@ݾ:51O��h���R(p���?�ߠ �UZ�u�^w��>u6z�ټC��c4��H��U���T�P���kI�w��c/�3���Ǯ��y-��[�To��O ҙk-I�Lx2�[����qߠj�h�i:zt�q�?�F���0R�i:j��I3\�M�H�v+`��Ƞ���@�'-*M$�6Q��8M�t�2�%-ѝ�mi�b�J2}�/dJ��Lա�L"v��\�Z���y��O�#�<$ i�
P��p�;;;r��Vъ8O�W8�ga��H ���S�S�}��<���F��|n�9��Sb���p88��t��v��իW��{�,>M���O�ƿ^&��������c�M���B�p�X&l���Ֆ��1z(����BڴUna]p�)�E��f�J�q=�/�qu�D<�7�'v���0�h�B���@Bеj]�F�@���i�D�9}!@��3�c��7�h.�Z� ���e<5p�,b_�:���l0.�� � M��dc>�<�^�}�����O�-�^��v._����l����^o����e�o'����i�ۥ�Xu����9yJ���Ӑ��0I�(�<�=�Ǣ>��2�Q'��ۧx�����nnPwo����ed�h�7R���^�F��q�U��w,�=jU�-�ww�~��d����#�V�����k�7�s����f�S���k1���W�M���y��$ϛ"���h�R��n|�y�H��_a;<Dx�Iy��C!sb"���GW��Dk)O����WK5I�0��홨��r�/��	�"�Js����lZm�rZ�U�0��`�D�$��i�}kkW^ W )�D-����5�8�2���*H�=�p��	UD����DZ|G���_��k����p���ǿ��/�����7.\����ZY|�����O��x��q�4����&��q��Aƴ�@&�}�h���7N��)�F"Od#V��zSB" n~��yM�9�z�=,^��`���J��G�9�i8��� �\�nP3�v;�1��Xh)���Q�&�U\x+å}I��G���5���x�E��P �i��4����g�Z��l���?q.�٘������V��$�W�,��6���60��j9y���q��N@�QgR�A��-��O-v0��ޥp0�N�K)�HM�&~Ҹ�G;�6��h��qZXZ��F�F�G}^;�MI�=(Sk2��vh}�I�Qn���W �x��36t�>�s��4��j6rE�'�0F��;�s�TO�3:�%uLj1ub�x��z2�v�D�.K�fA��B`�Gtű��$)ν�}�~��8oZ~h��~ 0S�(��$3�#�j������8��g�IjN�eiQ��y�^o ��}k� &p9�bc5�
�[T]�D8+$"�+q�"fS`�F�˦"Xj���"J<V�vw@�`��Q��K�Y�0���c���z����k���;�x���h�D��^�($FJ�	�fEXӢw۽Z�Li!ffD��\�Uf�v]�`Ѐ3��׫u�3�i��P�ʑ���ch�i�Ա������ 8A�?��R�2�4��kt^����M�VU�4�T
j�?�r�ڹC�0Ѷ(^&�ڠ(�~[uG���i��>H�� P~V4NU*ɴ�V���(V}(M%*�<
cQ�����a����7[��-,,�ҥ�W����1��wwO����[=�5�݋�v7�a^�Hm�R�gO	/i���Qq�l�"H��7�us�	��-Z>S��mC��Ow�(�ߕ�Y�ETS1h�y}��cui�z��[5j--Qku��Z-j��{�.��Ր��ս}�u*���:kUj�C\(�w��1G#�e%S���t���C��1Π��F&�gۑؠ������"6��F�1�m����mD����RB��i��p��q���R	�'5=9'��L^Mb+�9 qPX��5p#D�p}<u4�f�z�����!�p�b�*Cc	�����3�T�Y~�o"w�"�w!����qZ^Zg��N)�|��2����8(�c�[�vo��ن6�8!�_1��,5Q9i������
�dN�o!��h 0� ��`�WC�ЫJR�A%�z�x�9�D�/���m�}�ƍ;�����Ǐ�!�h�������Em���+8����)R��CUS�����DX��l�(6 �hŜ�݆z����w3����ȑ�(�~nAbO�x�����І ��r���t ��cЄ��h��j5��[�5�9U��3�|�g�B�l��#1qTh7Y7��d̾X�f(��x��R)p��ı����+��#�Rp��f��+7n�w��%
j~g������.�MkiyU�!����+��(�(�6)��%j��
o�A�Es+����穳}���4��o���#p ��wnR����
-����ʲb��B��[����lP�-9Л�ת��d�,��h�ܽ�����t��!�8�Na;-��A�բ�I�i>�T_KW[6e
��|Q��>��J��o��mi",͉
�Rj�!"L������d���;w6��͛�*J�������=z�i�Op��C�$����qQ/WY�T
i�b���!�j%�F<\S���0 �[���jG"�+K�"�����a��V�xu�a�s:R�i�IH&��������'��@����_��*��=̏�a��}�~��_��<�p��%g����hz�z��S�A���}��!�d
%�@{��P�QY��������p��>�/� �e�㹓���l:�>�/�)�fIj+�����sE�����ќ)�*�s��
�I�	"GR�3!�� À��@>f���$�S.������ㅅ��y�����gc6�ǫ���3�W	�S������}Iu�H�)����lMuh���um�(�F��-�U�$�R�jyYz�Ux-﷚���&l3�\��6Ү00���Q�\��i�ӡ�ݦ���,/P��g0S���X��7ɃF�L�Ј bN%����h*~NU_M��Q����=�Tz9لem@�u�cN[�ؓ�Ҫ5_�J؎":�F�+�F�ȁ$��RqV ��fqT�/8�g2.�cD"Kb��\�Bw��5�jT�l�~N l���v-0��^'�P�_���`á3g�����4k��A�����&|������*�&}��ն�a�)��d`Sa��}ר����vs=�KO�BL������
2N�	�q���F�PE-߅�[�Ǭ�g}��m?��W����K����Gο��=�x3��`C�z�>dE+��H���i�4]A��W̥E*n8�P�~��9��9�U�ߖ�b�j:��C��+M.v�p�x8>x������Be�����"{3�^!n�T���C6�b�4}h>�%8�~��K%x��<%�h�x�l�>����O�}�m��"?>S7�x��Y��lo�{��81�!Ⱥ�9-�4B#i��e]&W�6��lĢN홊\�"�.����K�Z�Z'֩��H[w�4�i��JJ�1DJ�ܣ9������)a�%1�A��9�I!�
�*٨�NP�=0e�4Dp��J�9��+���!��M�d�f8�����([KT.��M�K�n��)�E�2J��7��j=4��0X��P�f*�+&�o?/l�����%�L�"SI'v,s�Rp�+��D�S[y�8�}�[�$��/б�U�1�=�a��U�������rmʒ�Φ7Q'��a�+�G�ە4!�_�>ͺI��L�|E?=[i�N�Z&�cn���0�l��쉤Au/�ߜJ�D�t�������h���^xዏ=���d���h����$�{S&��O<+��7�#�7Z4q�S�9����r:�g�=�;��z�_�	��F�S��2M{@� �{�3`�ƻ���쭜:.B��O��j�mD��?
G�IC�ͦԤr%�#u j�����$N����}��}fu���ե�痗+�._�<�E�f��>.��x������p�;���b��Q*kmeu]��퐽t��qTЂ��C�B֑�D�t�>�n�p~|�"~n���5Kt�y����vh��Oi��.��ϩQ��Ƞ\��<���@6P���H4�J�#pU�;C�=��NG4Q��E��p�,h:J��������d�t���e�)�YAFO"��?gڡ�3n���X�V�(W})|��+ [���V��riث�k�����6mܹ[Dɥ�g�kd���T��Dg|�V��˵�Н���^|.Ǐ�S�՘j®�*�����?�- �T��<�Ia��GQ)�掶xI�$���ߠetz]vR���)4� ����s���c�%
'�H��ܱ@��I�.��=�|����~����ۇ�����ׯ�ٹs�/ܙ��h`Ww=�v"EN3I̤��F�E�E�r��{��V)�*o�o�ݷ��QGA�4p��sVY) �(��i~_�i��Y*߈�����	��@{�i'm]ԩ4�U��|w"�=��"����Qf��]7�S���znn�Z'Z���Oϴ�f�62�V��w�qF=v�F����ؕ=���E���8�I�;�*�\6�̔sX���pN�a��}Ԡ��k��B��E�U�-.Q��vve]��D؊��}�*TO�)SŅP-6h�M�@Ⱦh��4��s�l�� �0��v��PLE$��Fzݑ�<;l�����jJ���Cj���P�#\�>ۛ��B���j�Z��%��KE��5�&�/V�I���lJ"37nܒ(�*}��1h?�2M��G�4i��"���6���=�`���u��Cߺ�T�9*v��x�D���v�2�����Y�b!����Sn�ʩ�Mw��Go�r-��4�k6$j����ك"U�箙����!2M��z1S�m��騜�3}�k�\1~�Q�ރ�������~��S�輘��h�DH-g� c��:���ׅ�y���\�im��|gۧ��}�L�mX�w����0"�ލQУ`I{�9*l�L��:���h�E��H��C�@���[�q���m��tݲ�TF	E|�A�=�a,�K�sq�D!ʳ$F����T���O�<v��>���,�4o��Ǝ�4��F/N���j���$��퇒f��8��.Z����8�
�"��M�m;Y� K�ĕt�x0���S�7х�uZ[\���>�ܼC{wo3�H��1KD"��:LnY�2����Z	�=�q��UR�l��iǁ2i��q ���ؚ~���
OFZpgr�H�^S����h�}�ܠ���PU�n��Ғ��[����h���L6yW�PB�vD�YoB/�t��nn3�(�ޓ��o��YGמ��8����F[���t,��'O��%Q��&T�	�q���!���m?*M�!3 ����(މ�ȍH���U��:�q��Tn��O#s����i�>r<Rw��W�k��Ş����i�߾`'i�S*D2��M��>�JZZ��2�Ng����	w�_��:ڂ�3��`��'R�po�6 v� �B(���)5
Ű:"Vc	���1�M�%Z�������hnӁ�yR6jD#�#a�۵��D�L�x$�	��0��P�B�F[T����¡�WꛈZ�J��V���f��ыg��g.���J��V[�Ć=�;��B�2:���њ��Po0�����(���xO"y�h���I,��$�8D �y�lSEN�Z�(z��>�%������1^���:�o�F��>��:�#>Io5�	
/҄�r@i5��$���r������'M����Q�Q�d��M�Y��]U���b��PI�4���J�o��xM�IhЦ)/�ڹ�QW�X6����h�R��S�v�-�"�4ј7W %���$�f��N�M[Z����V�	�Y[[ˈm�k;;d�!�&����%!t��;Ew6�
x���-�C@���c�Si9e���3N����!�<U<w���!�P� ��H�X�9����yM��V �,w��Є�٢t�0ٗ��^�g���?yc�����h�bHD�2A���N7���ÜIӬH�)j�M�>y����c�f����P����ˆ=��1l4ɦ�`νx��	�WU5�+�1PѴ�i:Yb��P��j,���K.`���Ry�B�Kkt��5��آJ�.�ݠב4\8�a8L�q�w��:�/[_��O����g�p��`�QD�6�ﹳ�mluz�4ʴ�vL*��:}i��t�D*��A�.����(�h�M������&olȔ �d���K�l��'��P*�$* G�wc����'hy�B.oƛ7n�h8�*��H"&R�oj��`E�� ��4p�apCE�pJ.��7��cJ���M�X�Qg�znҌ��$5���Uu���p�@��3��=Cz��ר�2M۾��ՓrE������9W�Dv��F�'�/�x������&��߶�}�D�wB��d\Ӈ��%)���M���-���U��J'h��z�粼!m�N���(gN�����pz���8fz���V<pd�Wiu�m�^�9��]��蔆����9�[C�BDZ���
ތ,�;��V41�=�>�oܝDI�m��qYg�?k���S���E�}s��1M��%��&���XOC�֓p줄_�4�{��t4�tT� c:be�%�n�<�n�hfHe��<�'d�{Z_C�R��*�X��I���A9/�V*0��p-Ξ=O�nݢ��=	�2 ˓t<��p��gߜk�}�ĉ���t��k�.-}Oz��l��/�[!�c�7�|�3��j�+��&�PT�t��f}w�u�]:}��[�6&�J@)o�A_4�*����!���|̪T��i(�ၧ�Ө~��D	�A�or�,.�S�T���["��8�;5 `[j�^��mt��5g����4���6*S׃Ȉ'�3!JO��i�v�Z���y�6NISn�� �ˑ��Mq=)tɋ��t�^�?���!M����U�`xHZ<6��{��}� Oi��J�D�N���'�@�D���U_��JcM��"7Σ
>������&;����"��e�H�����j#]H�J��3��q�B��#�/�%�IMT�D��%O�����Ѥ�I��S��ψt�������;y�-%I����0M��/�/��@E_�m5�k<77�����d:L�p�9.M��^�StG��d�tɆ��HЄ;��C���H�V'G�����A��ɤ�����K��Rr�+w��q鋴����wci����K˟_\^��r��y�ҥ�H�l6f�4���9H~��Vwa{� )s�G���"��S�ߓ�����_�n瀮��*����U�$R�WOE���x-��ze-�M�H�}4{x��M�%��ؑ6����*���`�'r�;�v���t�����! ��.
\)�r��DS6'��ܛ���! XXqK�~l�?��[��i9ی%��j88�B*�K)�$��F�lt߾?�	0`�Dx�hD~Y�Z�cQ�Hz��+*�哤&bF��&��g�d�u&x�{�}e�jW��@h4,AzB$Ei�T�fVk"6F����6�o#����~�je'fF
qDO�I��-��}Wu���}�{o�w�MR�$6�6U��|�����P7����H�&F��S�������UW<�P$�uzM梫�"�x����"W�mr�G��,}+U�
-
Y��(���8�u_��ct��[u���\L�h�M�)�S,��L2%\8[��n��T�AaBu�[$�.��T��.��7��t�I[�����	7�nto�iS�waU7�M�xϳ�����2��f��M�nD������R/*�MǙϘ��#�i��d�8�c��X�� �����XTE�ظ�����j�]yr�ğ~�ȑ��4���yc�h��k�����N�SA^B��{�x��X��Qh�4j�M$(��#�6���m�>L��85y궫U��C2_[P�o�W�#� ��ޓ�$��/` ��n���WdfǅZ�xc�^�CS[A�"�Kq�jh��8Ib�^�4I�3WD�nQʍw�ޔ��-���Г������Y�M���c����ʱ
�g�IN�ͭ�D���|�V��Vollѹs�Ե{gRM*�nu{d���Q�V�դ�H�'@���!��)G��L8�0��d1I��
8��vP8F�`�K�ٌ��]���5Z\XR9��H|����F�)�)_\A=���>�V(R)Q<�d%)�i\��(U�~��>!�߯��TU�Z{L}O|Y�?�7��t�����h���^�E�S7 �� y�#��QM�Zm�F�&���Q�� )S���%ʃ^þqcK�x~/��OW�8��{�3��;>�jL�r� }�0�%d-m�CuH�TD$SM���4�-����3�4���D4<�w?1�Q/�W�5x�ȎɜA��N�?�����%*�s�B����4�I�ܭ�<��@���a�T���G�P�ZH�1 (�T� I�0�'��}���T-�)�Rz�~���v��P�����uJ�����"bkRx����3ևmn4���C��_ۘ�+�u$F�fߴ2n�$0�Ň�^sJD�b���'&lxY�&�[%�l �7٬w�����cBS���e�4]G��N���y�����P/�&j�dIE���86Y'�_�¤X,KU��ݎh2)�H�����2�����(<9N�D\�Wwm����K�J�"�P��i4k�����`L+������굦�\1��	e����U��g*ǭ�C}�������^����M�h���M��4��!jLX�of��m�8��L�T/����� ��32�7�Q���n��[���z�~Һ�2F���UK�o��_��3nw|�`8.D�rE���[aј)���X*���. �`���s�Aw_ZZ��Z�h���+mR,����Ij2��H��hC-Dh�Q.)� I��H�<h&uxA
�h�T���%�G؎d(�)�b���k��B��+���Ii+�b
��>����c�.7�S4�(N�h0�y7�N�Rp��YzZgΐ��X}zMd8M*�'q�T�]��Z�o@\}��ֳ`��r��SwU���4�,�J4�58~�JM��qN�O\R΍�k�t)��=@��}��y�+졐��I�u�z�6c��*��5e�%�,@ ��
�� b�;J���\�)2�[P�;ѐ��h4����@w�Cm+g�S��4���o���ۦhum]��n�
R�Єk%�,����-T�=�G���p����Io�fZ@*��HH<�.ߔT(:�4 ֑H+������hݤ�7 M������7@���� P3�Ѷ(*����	29�~��_n�qsE�V^W����9�݈�$�cT�|׵���0u�X���������2��&:������	g�2���-� ��Q2����ձ.��~���`ƭ4f��͏,��ݨ���mv8�!͖
y5��W[�T%��������i
�B�/�)��?R�@�K5j1�qy��%�h8��-v���,>a��3�p�H��`��ףl'�˴��J�h�K>Fڤ�4��)b[�O�".,��!z��9��5�ql����ϧMkB?�c]7:e"��)�l� C�Hq3��&[�Y�
��(�k{���-yδ���   3����Ҳ"�{�n�ͤ�_�7���Zɹx�i��L���A���Ӝ*|�Q.��<$| ��͈W�H �Ч��-��,qNm��5	irr\�W`�E�k�󴾙�5wf�']ܡ�}�P�� �kB��
׫�Q� ��SUvѐ r���k ��R��*�IT�5�,�R�w�oߞ��;��[h�R�v�\��n����8��/�`6����54V�]O{OШ(�%a������~��(`ڧʝwnș�J��,}�~EqW�7-�	�ػu�5r�pU:V�U���������vC��a�Ѩ�d��"��^�t��@�{0n�.ӱ}��z��\�K�y��M31J&�T�թ�N�M2���.��T+�(�H:A#�ϱ�,U�_��(�L�s�\ߠXfH���!JF#�V��µ�R��S�z�H&Os+=^���4�1 �{$���$R��K��G��t�b�v�LU��[�t	�:�g+��BZ^T	��7|"�?�TL�=U	g��M�#���H�]�&2��TTL�7]�LAZ ��2eB�c���/����K�>��8�J�	t�s(�����yj1P��DbP�bT�U#tG�`rN�!�d�b�`�H� N�Ғ�� \X�G*J���C��@E*���v��#B��'��(����+��ٲ�i묅#z\NH���*���7ic+G[[y}���j���$�=�;=ǿa��C�=_K�!�Ui%[� u��Cv״�$���J������[|�����x�r�Rm�ؓ�����s[d��B��Z�m�A��<�#Z�KT/�G�-��������IU3�H����S�ZɎ� ��lٽa�s����H�V �n4J�W��[T��U�_AP<3۳�!�ɎO����GA��R-_��عH�1���X����7[,M�	��P�nP��/k��.�ݠT���bT�M!�g1
�k�{ǄZ��
�B(�a�)��[���*�6"[�"ex��6r�֔da��>�b��Z^0�D��P)���*���d ����U�޲(l�U��V\!��E��	��8�qDʞ ��Z��	�4��/!�[�O���������@��8ԯ��R�|���>mt�T�I�S����:/Ъ�p��a2��CY���;x���C4��@> �*�l�?�����H\E�I����Pl��T��|�Z�N�k�6�;ZM��ay�w;l��(�LP�R�����u"�@o��<*�J$��"��ڡ�_`��fԛhoG7�ŋU8W**m[k6����X�He�)�;t��KU�(XZZ��ׯK�s!�.⨔@�I*
l{m[^�����	��C� "P�z�2�����;#�)߻��Z����?in@�-6���n�HW��U��T��>�u��OR�ҡZ�ݍ��EB�N�����s���L4p{�q��޻��?���T� �^o��ӁQh�[:��58R�.�G(��+X"⤚@z�aR���G�x�`O�<11��={��i0�3�Z+4>�\�?Qí�K��"'c	��;T��=�<������J%��<�.4�I�0d[u=$M��
m.�u�����¼ g��w�RRs\&+��P�E6H*m�H��HX�����Ш�������XT�"�`֑�sF�������m��
�� ��(U,�a�l7V��]bu��Ȓm�(����-EYp��e�C
H��s�F(	�@�V�����,�HY��Z�'txx�fg���sy��H��G ��]�uv�xn��F�ʆC��B�\�s�����	�iD�%b����:#r,8/����*�~�*��:̱���u+���G�n��ڈ�(�{�%OG��]��aRdl�2C)�(�<�����A��M
D�z�A�mpU�]��V����)����z�;�11'p��5�F��s���/�4	�h��F��h��6�@	F�l�V��;`/ �7V��T\�۲���EC�È�Q���
��N�Iʌ��R��~��6�mהi����\(��G��mmp�D�FÒF�t��]%ۦ�zk.V�K]&�"�5̉g@ԭ�3��10y@|��(|�->B-ڷR�}~-_�4:j�}v�\J�G(�HS�^�2���TI:"��v�J����ũl��OV��q+��;`�V������.Rs�LRT����@�I�&}E�H�6��hcm���1M��d���3�*�Ɠ�&-�4�|A�j4K�!K;r�.Y=I��{��3���R��7!�]Uq���f��H���p=�`�@	\&  I�y=[��  "�%��ӭ�3|&��<s��YJ$�J�R��#R%`#�R!��Z��iAq
�h��>x�j�� B 8^E\�`Cp)�n����ۜ����;^ǹ�3�nQӖ�'c�U7@Ň�n��\,�r��m�$Ⅸ���
������"�j�}�jC\OD쐝h�S�5��vRݖ)���D�d���_�o�w5���� 4�"ß���KKo�n<�FF2�j[9������	����xr������fO�oNq��&F\x�mnLj]iP:I���ݰ�i����-M;�T�0¸�f$�$5WoT�d�S��A$�ժ�>�ƒ>�O�o�7�������A�i0n���ы[�'r�{�j�]e�Өwx1��*�:ϝ|�IUp>,���u�B��ҋn(�����*�%]�t�H`aG���^ݭ	Wgdd�� �\((R0r�S�,NH����Wfy�KU�+�.���(�KF`1��W���3��֍hX�����|�q2$�~�ӫ�_z;��9)��(J���~����<��H{)��Te���lEPj�$d���ש?P�MA��4F�	�"�@��st����K��������vz�Sp��!U�>=�tB�K��Т����<�2����
@]�o�ke8����*2����G]2�A��;=����� yБ�x�2�I�)G�zEҢ �H]�<�S���u�����i��	�U�����}~6��<?==�S�����|���N�����GW����ٳ���:p����Q�omѵK�hzl��vK�t-G�;A���� �a2���j�}{�d?����tm#Лh7�QZ��m����"��B �o�=�����j&��3��oQ�5:R�ԩ<�M�$\[o6�|>L�1���jҎ���G�͡��ѻ��E�	�K��9��BQj������hR9W�/j��C�t�� ���D�yN�sT*���|�|B�*/v ���J�b�"�T;a���p8a��Y_�R���ﯢ�� ������� Ѥ{�d��
��l�'�V�9m�.͗��X�?%���.�p�tt�Z��dw �]�K����l�6�:}�5���V��"-��>QH�\J8R�ѵ�BZ���ЄW�:���3C�	Q!67�������Cĩ�5ՙ��C��*j%\*��Dq��BX�[��QO����� T@1dt��o�\��i�n"O��xi>�t��Ig�5�F����8nw�5�d�����om���<]�_�J��"iB�w�{@/R��0�㕵��  ��k�t��L&~�+��_���CW��;o-^����O_|z������f�x}�����O�d*)�B�L6���󴴲B���i<�j�1�8#��ʪ(OE#���b�z'9!%��+�{����㕟���s=L&|kLB��Z$F�g$��q��P�������0�odc�����[t�����B�q_�I���j�N!,q�?�V���*�n ��Kk�n`���<�<5��8
@��R���}��NDt� �&�o�X*N+�9�4P��Pq%�����m6��R-ʄ���Ds\Ӏ6���X�-���$�����5I�h�n���
h	6K2Z���y[G���d��|	�������V��=��޴�L0vmRQ�z˖�=G��:�J��TXq5%�e	�x�xs;��Jst�_[�E�x��3��τ|�9p��Z݈�i%�*H��ȶ(G����D|�%gn�Й�`stj�B1׍2��:>��/��k���Le5���>)�ڲ@R����c4�P O�����ޱ��-���Tޡ�}�F��)�,�38R8�z��]/��\�����?�{t �~������!:{�f�x��̹ǭ���r�f�]~��ݨ�)O���ym��&'Fi����$�I:��/�����`�O+��ϑR�,�bB�D�*���vwA18�X���!���B��xd��P&���C���-Dt>n��B�X��ۖL$��dTah
H��� �tc�FOaܕ��k�Nǝ�N�`�-8�Vit!W��zg�OU(sw|��e�kl[
,Tȣ^e�?�I�}P8dK��oe�?,�>�T��w�vE?��hS�ޢ�����S�١j�A-��)�U�r'.��f�syl�Z����v�P�	�/�����_mj�T�L8���PS*l�lɮ�O���k�C%�t�L�����5H��ĀD���*�48��#i��wf��j�@���,꼸��?�n��D�Dh�A�h�=�`����F��:uJI ��&�;
�
���	�sR��dpp�A�[�7@�G�۰�r�>��P���2���~��2�	2F��P'��5�z$���\C��EE� �Q[']������8:Zf��"m3�%<�k��>�@KK+�e���Q���f#F#�C�b�Z��i;�nپV:�~��q��@ӯ���t������B'W��X,5�y��Ѕ�^w�[9
T;E)�����L���+�f�㰑����Y��w/aZk|�A�' �C�K�E�_�}�7*���p����(1�gT�&�ږ� �h%�Y�=x�"l�	��[�p;~Os��O����nV��(���t����5�4�-;6
t�J�|��t��E�ZSJ�'F���/�X�}h�Y��#���d{T�|����P���꫐l�x��B,��6>>I�
,�Ut���A�C.�����*@��g�vD�1��$݆h�Ĉ|Uq��ҵ��tKW�	�et�#�|�AJR�4�)�#h0utk��j�t�Nu�U6�*9"-�k�7r$g�L5p�8$Q�#��z�*��� ���0_[�TY2鏢�b[����J2��Q ���eB��Pו�B8����*���#�c?6ڐ������8�4�"��h7�cJ�E�����_�g��>�����Ŷq�X'&''��86�p8� B8n92����� �����:p � �Te[D���(��bs�Ѣr�'=D�E	{�hmmC�M���5��ojۄ�ךh>)�z���^I&��a�T���� 4������^|������v+�����4�K%�۔
���Q����kz/wL�f�DǾ�v�{Tz�@X��ۢiF���,W�[Ti�e+���u�Ŵ2��c�m<WU8@Y�QojO�?��醫m�v�Iǩ	��8����X+ˋr�0#�a5��P����s����$%2
��_�5�<����X��~_�T��ܐ���������-?����G6J��k3H�Ey��1�F�ꭶDeÎO)^�ꍶ�y!89:J�L�BV��+�teu���Qr����luh����T(Fl/2#��s紤���6��Q�.@���.0�&��t�Ǣ��Z*�T�O8O
�X� ��Quu�	B��~�� �j0�[� �-��B�Tj0�a��bK��D.��>��"N��N�ϳ{NY�.@!*֚m����p��HP"1�tBiIi�H��Գg"O��	H�v�0D�N�8A++k���(J�Ī�>�\_E�Ħ�NW{H��:y�)C2����#C�H��#����O^�mƣ���?c{�f��;l��]�Q�(��(o�Q�Q��7)�� P���k�s���D��2������K �n�T�~�\œ�mTC�x��Eh(��{z���nڶmR�;w��#�TjG
���d������>���CRq������������co�YZ\�#1jV�t�{�@|�i��?B��sh��Ѥ���/]���Ti�U��!��_ZY��V���C"]�r��yZ�ڤ����N!��I�wJ�g���#DJI�r�%��{C՜���Lx9&�dn�~����Cu��-�oH��MU0����=��4����t&�_��w� uJ��K��T,��l�&'$n%O.?���-7�<�rt�Px����2��jå0"��!�� ��ۄ����;�օ\]�T5ihb�2�6Vi�^��;H�5y{�D�HT�\�FG�y[�nU$��&��P�4�/JHav�@�^)�J/�t���64sY	��^r��R��HE�=�T���\'W �j�k��=�%����0���Q��v��{����zwgN�T�=��R~4�6SUi��������j\���!9x�~`���f�ҥK�+��p$�W *�Y2U�D?q�T�N�I�&� ���IW���r��tzvxx�k���k�p^�|��iD���g���نO�qE�<l?���chB�?���8P��
�V7Rf�.t�u?�L�B�|���ӫ���B�������� ��EE#h!������˙L�簾�j��������ܸ����ϣ�ǎ7���ݫ����^�bc���=ɤ
&�V����f��˯��g?F��0-]�����	���F��=����О]����4ϓ�����W����S4}�~��7Ov(���'�8{I���H��Y$xFe;i�ߔ��"���E�tŝɪ����w��S���@)��'�aRn*,���g����?+�H�S�'�*�I��w�t[�����T�P��V�3�hx�*o�c0n�q�L�����V��=U
S��zӣ��a��ttH�G�HȦIs=M�j�����;OPC�qvp<O�5
��գD��-����6*��Eg���$D5<R���'	8`łD�ca�"Dy��u�ȡ��5�ܤI���3pw�����׏NZ��N� �b�J�&|,��N9Z�IRr���������5TsŜ�\I�����%�	��
�w�!`I����X�V�v{{����_���tLg�Z�@5W�����
C��B�rչy�exU&b�cB@e(���LF@����(�-���畑��S��c���%��K�����֖�c�����>�	d��N��"Z��� �!�������
`��U[���H<J��Z�*
� c<	�PnG���|@{b �$`4`��~�5u�� ��yK����x����|��Ɓ���œ����w�����|�8������O��}trsw,�����;��?Z\��d�>����ѵM�"mň��_x�Q�ً�鍿ڠ��8Y�嶶(;>A{���;i�ѻ�R	:�7��c'���葻h��5�
EcQ�:M����-��Pi���wH��8ި�Ǣt.:���A:�L=���p�M�'M�'������n��j[���=���Ç�ǯ��u������O�fs����>�"��k<�/�`�-4 9��z�޵Z��O�/�58H� 2�f����� PЊ���T]hu��[�Ս���Ȑ�P�_[/7h)��Cu�qM^]��S��i%�g'�R�$�D�]��ja��Y��%�4�vFǡkNʍ:n"g"�\q�|_a�@v�T�&[K��#
�*߷���g���-�2D���7`z�i�*�	)?�Z���F��� e�0CT'ʈ���tq;�n7�3���*�#f���իW�a���y�]K� �cH���y�Os\*Z�hhLY���y�����*b`rexx��۷o_��h�>��~��ӱ\nm��V�AE���j������tF�	@G��� (#�ixQ���yS����Y�0!}>�R�tZ�FW�kk��n�yS���3��Tᡁ;��o�d2��?��t������ynyy۷���gN�<�����<����+�mb[������,O:Aw�X�W7����*�S�U+3��Q$�� ��	��3S;������oӅ��41���w�ɷoV�oAo�'���9z��O~��cq�\X��~�}J%�tρۨ^�R=�%�:���|���H��D&� +F�r�=�\�q�G�R������I�À'��C������;����n�nc�T������4�9<�:���|�ľƟ��s�f���4G���ʮ]��h0�Ǌ���f�[kt���]�!*��5^Pxn�-*�������Lcm��#:ލZ�3�Y
�#�^	�B+��K!F�P��2��Rjt�����u-�T�Y-V*��+�HQz>�2eSIi��Fd�略dQ��R��t�N�Y�6�K��R`g^�*;��	��L��!�� ���vT;��%����J9�&�_����t�.U���<W˩�*��z�F8�'�a�١$�f��2A�*O�w<x� ��l@4M=��h[��L�����})f�������Q�*��z6������kZ����!�������Od�#_��6,�˿��?��bP��8�`D��^�����T��E����G1��q�:���8!u����2C�x��N8Q�B���M� ���[|��w��E�gh�> M�c���۟�����_�S �@e|�'辣�Ы��AC�L��I�ͱ��7����T=}Z5��Ì��<��~�*~�6��<|;=v�m���]a��p:C�S'h�\���8�9	���{���m;h��hv�b|�W���]�hs~��l� ���{ǎQ�j�>��g	أm���
���h}}sM�1w���g��F���(����.�I�&����Ͽ�.���Q���Lx���,MNN� ��6u^?c0n��sW���Y,4>��t�?�`�AM(";aj��@
�P��'G<I�#Ҡ*��ò ���b��cֈS���8;Hh��U���>���잦0;P�J�� 5#��rq��4�d��� 89׮S]�A<.��Y��8�OD���`����{�%��kR�.-��n���!;ZtWyV����+�����3x�u�*hYQ�'�~��\�0��b�};$��F���q(i�ž��xʾ�#*����tV���M�8�|�x`�y2���(�lQ��}�
0��Į��7�Z�(��UqP��%�%���k*3$���f����`�j���'O�|kss�K�F�c��{��;� �6�t�l�(D�����0�r:^CT
 	�I�p�y�&���( ^n�g�E��}����ջ�h5
��G�^�Y � 4��G.�K�ş�?�ӫ����S����;����<9�t��h��6�r�
-��ж�1:�s����y*׷(�o�jWf��`��r��7�ȡ���:t��U
�����e_"@��=F�m�O�?����k4|�"�v�mgø#>DNۢ��}�f�;C�>LN�Bw����_�A��K�W��l�H��vc����1�56�%�s�D%M���f�ly
�(O�#���k"LtCZN*?<O�+Ł0K	(8H%P/�z3�Q��\��`��~0�V�������g7��L��C��AB��@�\���.U �A[@�D%�65��ҍ��1A�g��%+�Q+^�/PU?Ot�OfhxbB�y��ج1��@Z����(�6!��!@irx��FKRtx ��T �!i�����;'s�n��DF-�(H��;K�8�6�V�0�c[�+� �W�>DO	�j��j0��.E#�6��ʌn��y���B�T�IDʩGM�%��QN	�I�	�iw�$l &Tz�f��!�J�t]�w4����K�e&�٧z.�r>&DUD̖�� W�);"\�D�j��2}�_���܏:�������.//?����h�����w���e
)B�nsk]@"O8V�FA��8\< � �� K�G�h�C��*P$����;��%����y8a(�N�~4��������i@ӯp�o��K/=z���g�N0�1�.���ӏ=&�o.̜�|.G+��4{�=���������L�]z�ғ�T/��S���Ca�������P<9�e 4:6�6�V�)�}��ҥ�c�C�M~����s|!V���s��t�_����N���0���;�m�J�[N&��-��m�Ѥ���@�S�T�I��Yr��m�)Q�uM�^�]���Y]��{=]�,8�e��)��)���Ws~�b���J�uw�cS���	A�'N��~��h�NL�
��&~C�S���jS�g\$UP�["I�H�F���5۔N�8�(����u���VC�SB<i� �/�
[A�M���d����Sh�fӨ�����~�\_Y����PZ�9p�L*&�"y@4k�H��gd`R-S�H�+�����l���R�n�8	���#�f��(����� 8V鯎'<q����OxH�]1p�FcB�O&�4�2�/-R ��@��q�A���)���l�~�]^���C?u���1@�ޢ��zB�G5BWAz-@�C�3�L�;�w�n�"����(�w��+Wf�����r�B��[^������6d�ёq��P�Z�M*܏������ڴ�����#%�8�SCv��VW�	�@^��	jb���=����顿9r����s~��+�11J>���������a�Ȳ������ر������!�u��7h$��Z��&Ŭ�=t��g.��^�t|�VK�-6���O!�J�7_����&vOS|8C6l�����r�J��q�Ӂ�u�D!��FF��t��өQ���thz7U6slx[t��$5�"a��yJ��R�'_&;�'f��*�k5���9!�G�V�)����XK*dD�N̉�)Ik>� >�V���C�ׅg0�ݎ� �P��.D*�r㱘T%� �4�acӢ��ړ?���T��9b���ҿ�Qd�6�&���9�|�@�n�C����(��s��
��h�E�QJ����uc�N�j�*����!�K$��b�g��y��kUjWk�I�E|1�1���,�&�l#"AK�)���n�<2/���Ǥ%��~�# ��ԝ�V�:�D}�W LCe� �Bd�S��� ���hxm(~��+�C�S)=%��)&	?W�*�A��Wi�vhn���I М�@��&�ۡ��P��hJ���]a�7�zK��x2%�2��d��&�����A��U=!��|,U�9�T���Z&5D�-���C����T+�d�A���㺅ɑ�g2��_���S^����t���������7���m��)~>�Te,�ǒۑ�R�  )����H�g0��pskK�x^����Q�� !>g��x�h3�K$Rs�����1��?6��W0�f���w�
}q|r��Z�J�)e��$��;oE��8�q�������]����Wh���M,;�	������	�J���*m~���+�k��#/��:ѡ4��*�<�Ii6�W�ΐ_(ҝ;w���-3h
3̨�7������|��v���9MK�-���4��� ȭ|�.��@iY�<�����KͦSd�d�RwW$N"��D���&]-΃H�+��H7O�4�NP>�����4 H�%� 
kk�����ɱ7xS�+�>�q+�˾��X{`��>P�CNŃ�%{֮*�wMs[��5q��G��!�.P��VD����ݭ*�`��A���աvS�U�^��Wb�E�
-���s�ݠ2/zဪZ3E�o��U��t�7�-s��mO�
޶�Ru��sT
�ᮎn[F��p�<E&'��aԱT� 0�B���Wr��BJD1��p�Z�����\}�-E�(���WE�l#x�"U�&�bIP�F�2��1�Ѳ �D�T�ϗ��̹K���.Տ�z�qb���ܐ>�@,	��D��@7R�E����S��x�H}!R`fR�:-�%���ȫ۷o�Ud�whpr�����2p����C�r��`0<�j5B�"  ����1�x-�{qqQ�G��+���j��4_� ��95���	���M%��
��[����l�����KH��4�7�'j~���t�]G�$߻�nZ�2�^B�N^� ݯ����С�hv��hr���{z?�w��8~���M��&Ȍv,Z��HŅe�L9���R1O��E�|��R����q'm..�^y�jw�A�Ω�Q�<���wӶ<H�Vh�P����$�T<�v��Cwn�W¥>O����aZ^]��c�侙��6��s���/BĮo��F�*�.2&p�T$[B�mxm�]��.w�-]�C<����!6���_�s��%�^狫[�333_��;Z4��0xڏ/n��(׆�-�ʼ�Wء����C}Q]��tM@�0$ऍ�b&XP[.��xApDE���#�$L_	����X���b��Ëv-��Td�Q+�)n�M�_R`�0��~K�5O%�6#��V:NMj�mG� G�y�� ��U�uK�M+(R~�i�����^j��'Ŗ���I�.��^KdԱ8�"^K���vG"�ғS/��B��I
e�(ʶJ��+.SG C�T�o�K��4�.��KfҔT�]&#�����h�׫���ڵK 	�Vȱ�N^�D#�N��cǎ��Tߵ_d��;�������ɇ���>� �î�Ce�B��W@��C����yI5�SJ<3U��b�!ׇ�]ALD�Lc`u�����þ}��~V�w���_��K����v-�KN4�v2h�8=���������[�~���=�S1���F�r�ξw���$��
R�X�ͭ2}�')�����>kU���SG����屮�� �7Q��4O���<�9�.����g?C�j���9K���R9O�/�#��NC<�]�!w��G�}��d��E3�kt�G/S���#O~�^}�u���ȦT(J��$5
%
"�S�AW ��*��;z�ފ�B����)��7_8J���⯴���`ŅjC����u�?e ���>K��ҹ�3�m��zy���gO�������M�\����_�������ʭG�
�ZUٷ@o��B8�oG\�V�趥TE��y�+�+M}y��:Ү����C�A!�۶Ւ-�CR<Dj��,ΒKA��Z�|s}���2�6ݖ%�N���T��%	���$~X
H�]��MG� |`� Rs��e*�\h���+EqE�V�:G��	6@D���KO R�T	 ���2º���YJ� \�&��d�����F�_���"7�ƸҸ���3`u����}��e
��k5�n�S�i4�~�^�lڭ�DY ��B�	�FH�"��%ctt�vFHP;u��f���4:�}�U�~ţ/m��_�z�G�|��\n�ߕ˕:^k$���Y8 ��FKKK���*�D"%�	����@s�[U�A����Ġ��>z���_@�/8��
ҕ+;���/��ֻ�����}��@Ȋe�P,H��0#�O|���V���_�r��-@l+����2}��ߥZ˓�?��lf�~���4}�Rl�^8?C��Q�~�]t�/�U����8]y�M����ɏ>M�7_�W^|������ΣGha���49T';�r�F��&�)�h<��;����3�ۼJ;'��x��|�Y�&��	F� ��r�"l����A1�#&6{D�F?�j�*E���TZJ;Ť樂N#_�Лm�������[+V(`Dۥ�����|����@�kkb�OV0�@���ѩr�:�)7���X*�?�ٲG����6c^�ynJe�
6Q�V�Њ����mI4B��l�ZRJ�Ȍ�m(\��	��k�tUnWG~:P����PʎHL��v*D�B��2��R����5����miAE2J�*�b��ѭy��
��4=���K��}ΙTP4��A�f�"��iQ�	p�ԝ�%���m)rA0:#��s��:4:������f�*�,}�_�T�!�����:bs:2�:D�ਢb�P|������h������7�F�.?�5�͈-EZ���o�m���#[M��{1��FF�_N&��~����;���[�k��.̔��GJ���Z�íVs;O 	�Q3ط6�uBꮿ�
�+"PR�jE[]WQ].1 �S�~��h���r8���>q���w��cO/,.f����^1,v4H�|_87#_��?�)!�];�2���v��t�^b0��hdlECQ��T
Eڹ� �F���ŭu���i��շO�z�Hé]{�$��1��S���-��W�Ny�㴰�IM�����S�ȡ�(R�ӵ�3���Bo��
=9>I�=���ht��/������V);9F���f�P]._������v��C@������`�@8�JS��S�U�M��W!v�
�����u�x���[oѥ��hmqI�PFUF���b�`�h�������iߏ_��>�R�=�ղ�eס
/�`@�sN��Dxj~�7d�Z}�RoG��G��J�����R��L� ��^��ߑ��ۛؒ.j*�+s�gO?Qnk��P����b_PB 4i[@��� �Rl�N�!�e)�o"�2����X�>]=��$uv��!�{ ~Җ�4�\.G��C"�I^K�,��ٲ����8�x��D�V5j����
�z��J��ƃ�$"L ��KH��9zf.����
��qKzI=ف��@�;��HHq�t�8��m�}m����ᑬ�(�%l[��_L����s��1^�.�������_X�X��b��v��h�^r�F��H$�ȑ#"���@�xO�2)Y��U�����_NLL���
4c �~���ǂ翿9��׿������Z�:,��+�`��_C��;'�&�^}�ua�q��F���{m����)�_zbh�.^��3oS�T��}�3t���T�(�hk�:�&�Q�ޤ��B�|�7Z�N��������|�S<i_��~��裟�$��~
�!,��tey�V�W(ēe��5z��FG>�ii�	Ӊ�,�U
��MM�`Еo��aCSa�t��i�vZO6(�z�]K��Z��&�b-�_h6 �=s|U-#�qW*8�B^B�;'��U����i��iZ���D8JIT���h����N'�Z���i�����4�q��^]���+��J�=��8��ty�T�9��'=)uT�6* �տ�-����q":b7�s@��V�#�MҨ�Ӗ�;��&S{2��j	�.��P����NԿ�����(ن{$`��b�:U�Sx��� �I��v�Q��^�+ ]I�RlF�H��+-%�ۄ�j���E�@jqlLZ�R�����s��z���3p�yH��ᲅ�JI=��:t��r�E�@˱�Iq��;|�� �;�֥�E~yu�ff�H�S[x8��:u��ܤe�3mW �y��-\@�i�6v��[�.E�|���ɤ��`�䯒��~��������Ͽ��Q�����g'� c��f��TjN$�IZ���8!%B�zh���f5���9���}��_Z�q ���@߸|~6U����/_����o=�x�ħF���)+D1�ۥ"�#�s��,��[���w�C{�w���*��hkc�<)�0��q���~��i�{����ŋ�Z���~�s��R9'��ŕej3@zi������C��S֭0�85;��`#���＋����!.\�LY�Aw�v��&��7���u�_rb��J:T.V�O�w^{M�W##���=)����o�<�i�
�R�u�PR,i�^�x_d�j���l\B��d,)<��O�닋B,�61A�ZC�Q�n�Rh�MI5�1�Z�=/�����u��������[�O�W�Gr��W� !x��9�xF�Igip"|���%</�/K�MB̆����>av�:~��v�j�6U�m޾+�a Kpz@����V����-
x�x)�4���iy]��:����z������J�	C��|�1M߿�L�Uކ�a;�qm\m���'ùT��Dyf��� %!U#*�\Ǔ�Cihn+�f����J%�Z*��,Sb���2 i��itU���w�|GPm �D%�����ҢD�|-u �h��0���VT_�I��`'Z�ۄ��gS<�G�FF�466"�7�) 0a��X�u|tt�+��������H&��W�֮���Y|ps-�@��:��e04�� ��H�)u{�T3���������855����~��7 M�c��s����cǟY�t���?����Xx����p��9
�*���)_ܢ��u��1Mw~�T)�)5��{��/��W^��_z�b�ϭ-S�]�-����k��m׶)��g�������Ju�6�H�e�	�ع�vO���z��SD�x�N��M&t��ߡ�����K�TA�i @O=����C�	��W����C�G�mr�F�Fs/��m����YZ+l�"�	R�]��kWic=O=�Z����!
���u�T���G>�(	TX�<zA���Yɱךti�4?~��IEJ�=��~S�=��Ĉ��Y!�J톻U,�;��Ñ���|�O�{�}��\z�1��R
��3��Om��T�Q��	_�\&�����j��r�����,/�-Q�P0 )+�^D��C�1n0�R�ڠzCj�<��,�oS���x&A��e�fa#\G>�HP//:]�����"u�H�dwE)�t����n�^TIHJ�b�KŜ�.3"�D|  �Ok-y�J��M�;OE��9W�z�5��F���t���1`b.Ɏ%����8'b!���u�󹹶��Gij|T"S��J�3�P�Y�E~e}��|�mIɅB*���ͮ 0��Z�WI!�� @���֨(C�X4���wK�z�{�n�&�H�ڠ�/J�+�w���###g�%�L�gh��u>��l�o����8Q(�����C��Z����+[�?/�Jnbb�9L+������2YZYY�.]�9��~�g��n%����υJ��:���S��_���,5[*-�)؄@Y��\�{?|?���܅d/�������}�������O���]�|�
[��0�X(D#�'�l��t���HU*e�Xk<��lȢ�T�:�⩳T���|�ԙ�Ny���Vi�'^u�2�(�Ӿ��'?6D�/�Q�\�k��х3�(�����F���+���BV�%�����o}��h���4��D�Klm*J4:2EN8LB�5��(%��B��I�i�%��8�NS�R�^V�y9�	�sk�Uz��W���Y5�&�ɔ�|�}`��J	ǼR�y����F������|��|�����a���_Հ�P�;W+��ߨ��Z�������t<,D��p|T����#* gۊ��Y�V�$iu�$oG�>�>��`5DY��Ϡ����D,vv�l��E>`�s(�� QK)�"��8���_�$<s�����*���T�=bDJ�Zq�,����j<$�]��3�,�SD���B�71([���}��3�<�cÅ��O�B�C���u�}m
��d�#�R:2>����_�D{�5�<sf�Jl-' �/*,N@s�z�Ǟ�]�V��P�Rx�ۃڣ������a�8!���~�iG����#߃ �+���8�333�0�����p�Z}��ҝ|M2|<^/VS��+���?�ݱc�/��t�����Tyeexce��co���[/�������ߎNM��Ah�믽H�<A=Lg�"�I	+�g��W)���2�@���.����t��2=��34����L��7M=�05�ഋ%�
�]�NW�����Y�
�<�:�2�d q�#�Q���s��N�9O��E���3{���F��z�lb����V���-�K���Y����7���V�'t��l�V̍<x��N�X^��J�HW���(�a�d%"t��#T���^.��;���
�����f�$�6,� �M[4�ІF7��!|�8�{iMZ]\���O�����~	v����3[���?�Uu�W�Us�E���c_������Y����~���c0n����Z����R�����=�j��6ݶ������Y�/���l��-��C�cxK�,!�T�%�嫴��B�ʍ�5�٦Z�!�n7:d�Q��K��i�e;N(Hq�I�J�� Q�_��V�-]%�n��P]�Q�����);���<vSs"]�I�DE��Q�����T�\-�)�ej`"E*6i�I���ۋ���
�V��p�Q��93Na9�h8��U�|�B�kN�i���{4!m�T"���Q�}����s���F28�i"}�Г�A�����'�,	�Q='Ⱦ�unth�o������ȿ��z|s|��;w�{�Je�뺻�����0��G�W=�&= �hm-v�;?�=����;�<��h&�(�;��C�:w�&&�B�{��i�Q����I����R9_�R�@5��^��w�c������h$�F�Z��/^��];�P�R�ĞAD���Kt��wi��y����<؛C%G~i�B�����Nљ�����<�s*��c6���[����yz�/���U���t�W(6<F���2�&O���v�ݔ:��
<1�{�*2�*-m��ǈ�I��(oTh�=$g�^&��K���\a����ŦtЮ�-��M>�������0f�����ڕYK����iB�$OG������mU�^�٬��gC�ȷ8��Ǐ�p��0��߈�t*O�k��7��P�Z��I7%j�.��e�x���;��~j�dm+����Srx�}��h��T��ꀚ?���΍���h�5^��A�R�:��@�;�?�*��D�Vw��i�utSU�Ŕ�"|�_-�Ҭ'��E��DJ뉴¶�+}���u���%N!����Ĺ"���SſJ/�Ow��(���'M;�䄅F��-֠?e���u[J���%iq
k�l+����"����qp@TeA G�0`���ynӍ�Mh�#�H_]�a�"&''��T)�$	��M����z6��\�ܡ_ˡ�O9<���v���:�ƃ&K���[�}~���'��?}����#��d����=��>O��ʌ���"��._�J>{^�Z��]�h���2�V��^����Q���#�����t����������8C���gi۾�TY���k�t��%�,�R��,%+m��P}c�
�˪+y�N.O�
�.���GSd�$��o|�R����ie~����;�#B4ϳ.���nP~y��U�@$��0D��sM>�0E����"��7�I��Uj�K��(�m;v3����+���;(62L3r^}�%r�=p���y��z
�!��H�F��PūI�;G֠�Uz3g�Ѕ3g���ձ8%�"3 �j|r���v�/�k^�^�5ͳ�d������'~����P�_k�}0�W1V���*ݛo��ŶM5�K-%mK�Dz�Kы�ߍ()1I�lW��mK�8 p^�^�rWs�H��h���1�+H�A. ��l��C �V�B��!B��)i��Q�X�}�ƨSoj*�R�$*;��I�%1���Mɿ-�o M���3�9�O�ǙO�*@.�i^lA��t�:�c��NxX$ �tDSE�aH�!��)��]�&@���ݡ��u�H )��i�勗�Pj�Ѹ|7��̯�VG�����z�kEpB�ώ�X�
���Q\NMM	)ZRz|ܞ&�7�Mlhhk�6q����}�Z��v����Ƃ&#JY���.���3+�����;*n+�mǸ�Ǯ]�H�wl�>� ]<y�6��7^���y	C{����^X��3�c�`rhH�U��$]�I����Oi�����d�R���A{o�GHVx{���|^4��w�4�@v�(�mǜd@��SOS�٢/�����>F�~�sTg���k�Љӧ���{�Wi��Շ�x���3?�!ͽ{���������O=�a���菿�_�����|�m�z�J��,,Ҿ�m�x}�N�{��|�q|�D�?D�J��ַ���1��ݔa����
���I�C����fЬ�� �M����3��mI���P&��󛘚�[;��jg�XX+7�ϻ��7?����G�e��`���&#�V��6%ˮM^�_*�@Nh�]տL�O��%�f���mR_���,�J� �$·4� pp��6
�;�&��!k�x�cΡ�� �ޠ���$j������+�_kB��Oh�]�(u�3*��u���tjJ	R�5
�jѢ�U%��+�m[���G�2 �$KiY����Z� ���\.W��	Aݖ4�y<�d<&�,�Ѐ��i5���2w�V�X$.doQw����Ɏ*"E�"����m�j�j�%Z�U��e�,m��=<�m�FS������H�\����[Y]�㍭�׷��O��͝���^A������ɿp!��Ʊg��9��/���Ό'
'�D���{���{'���E*��5�T��I䦺�'�6�����(ݾ�vz�A���,-^�Hݯ��7kvx����MNѿ}�)ٵ��ltV7�x҅�΃i��d?�����Qr\י����Y��o�*� A $@p)�Z!Q�%K���˧{|N���Ϝ�i��i�m�ۋ,��(���/"	� ��(��Bm��r�������*�ힶǲLI��TU!3##^�x�{�~���Gz|c������X����OKX&w�ٍ��t�-�������=� �C�"�I!�;`��:z���#oX�����q��	t@:����0��pBX�]�����^�ͱq��`lx�R;wo���u��p���:��׮������ ��>�vF>�]�󘞙����1zcD"Kv��f�UD�����l��/_)Ւ�x2�I]����oܽ�Ǜ��Yd������a���_����2]��u(_ѬE�6)4]�tU��Q�z���uhؒXL9�L1�q*-��E`���Q,=`�fZ�f�K���ɶ�X�Z��b� I� ��7�CG�6fn:����t����D:L`��o�L��tb�*����)f��X�i[ÔNh +%bPdi�&�k�S#��Q��7��!g��HPm�sDR�������Z�(�����)�[��M���>�bY�v`�=��8�T)+�4�j�o�btt���K�m�J��IngN��\Q�^i��!�e�d�*��9��/�~m|��tu�٭Ve����<��p&��{�8K&S'�ѥ7<�G���jq��w��M4���}�;���7o|�֙S���)ۀ݁�����	���=@O;��I��$�f�Id|�&��%��l���S�ٹe�hmڴ	�����!�֊�u���A4������"�8
��.�抦 �'�&|MA���C����c�0|�,&�n"���3琥;���A�Y��7�ɹy|�˿���.�ǯ�,��<i=��kb���qb����:v��PL����ſ��%2�Ə~��>���A�ij�]���><��C���¥��Q.��G0I;�N_��C���`O�p��4�G��M2A$�1|�|��܌���n�J]9�[��=.�~���T.S��D�J�nܵ��{yd��'��c���զ�s��|�h.�t]Վ����]RL�TX�L=5�?�8Z�h��%�&�����)*� *�)
�-ۏ(}$%`c�"�( @Tbq�ZE>�Ap�O�(Ȅgp6Ð�Gn�f�Đ�5�r�P�'$@��bx#�`g5��Y�fz�z��jԖ�Dܤ�M3L�3^����f���5�Ĕh���D�[t�Y��P��,ጉ*8��^��F�������?W����W��E�%���*��k��Y&����Ͽr�b��Q1�)��b��:=�&Nkr�!�[[�
8IJ**����DT�K�wq����Y�rd��MQ�ӻ��d�3�N�%�G���_NOO����)`����4��.�l{���#�/]��k���y��}�G=�]?�R���*����u�W���X�׋�o�ͳ�����^)��`��u�?�+���e	g����w�>�uy0�i����yq;�@zzy�M�Ϋ�9L7��BUv@�,�3c2ɴ��p� ?��Oc��8~�(�_8�g�2l~>�姱q�f��p�c��jnƓ�>L��".\��D:%�Wo��3�<�/�)�"�	�,��F1�����<�E�������x�������q߯}��} �[�X��s5�����A�hcO:��"'0��	���abd��7ŕ����ʶ��
фP�[��n��>���*t�.fS�d*u�P�=�~�W��'o>|����a����&ͨj�j2�5{ z�-��"k�9m�2L3"6~5,B$���*����6"!YS�*;m���Z6�EUG����r�e%J]U�Jq[�(�
�G�PN�[�� �q���:��)�M���6n��R:/:I�"6�!o]��3i��/���uzp4M[�71 ��
8�f��*�q�Ԧ��GC�ID0-�Y�V��f}8���aC��j�D�/���9�4����6����4�]V�.�u�����RU�@m,�!�I��'����r˱o��bbj�����'�Q;z��ߺ	�T�͐H�T7�a=c1ł59O������yc��L	Q���L���_�.	���\.��V-��c�_ͦ���d�ڵK/��8�[Z6|�%	~���
4����k�\�P(�����,���h?��g�9y���F.]zx�������:��ڻ;�:t���F���rg�}z[+�=�)�/�;��-�c׮�x����\���(��O���f޳��vx7o����F.��T:Iࡄx>�X&���.Qoomg�$����͡R*���։8��KW���������*�ݻ���w��e�P����;�p0���W�# v��=�����K/#O�s8-�8>�[�(�؂�m�p��(B�k4����>���
�s�ix�m��D���^�Q��pKWo YDO[3��4֭[�N��hK��G��G��U��ϝEgWd�ȶԟp`��V[O
��)�6�@O,�cS�b��кM�宻�|�k_+�������V�j[i��{{<r�r1�ƪ{4�B�hN��I+��ҿq�)/�U��4�q��PA��f��PB��ZC=�& �yE�;��Y���b�$�2M��j���"�l¦�Lz洟f�й)�7'���
˘d�#Ujʬf��S�l�bQ�4(�g�*��x�im) ��$�4�<�5!K���UZ��]��umE��)B�1��2%����T'E��᣹���Wu�-A�J��W���l4����b���+�����##��<�3'�IT�Pm��Y�5���:����My����ȼx<�lv�����撩�D�J�7�;�<N��ex�Xi�k��]�䵡Hd��L�p2��ñ��g6͙�p�?'���crr���>��c�o���y����7^|q��'���<1`��QGt&�������+�-k�^��'���#��(����ލ]�1�&P����P��������̩O�x��G��,.�|'O�FK�sKl?���&����c�n ���m,�cԳ6��������W�ͦ��8��awz��x��]Z�l{O',/��Զ���K�]Z@o{;��܎����;ￋ���we'�~�f�l]�t�� ��������ν���hi	�����׍d|�Ǯc*���͉�@t��z�e�����w	8]I.���8N\����<غ�7ĩ��G��m�}�1}�*N��왂%�maؼl�s��uЎ�ׯ!G@�B��70�L�d�f�O��s��;���o=q�]����ϯ��W�j��@п�ZJ�VS��u��V4+��ۺH}0��ʾsU���REDhq�J�����L���Z���4.@����C��/`KS�w*��=�a1��8�bK�*���Mn+��X^T���y$)�Dpe��@M�H�eY���O�������͒*�g�V$�R���F�`C�0�r::M��&T�Q1�4��dr��N�|��ʕ��n�lu�mb�ˠ��mL��j��I,k'-�� s����-��aW6Cg�b�WEI�,2�n+bf?�W�>�Uw
2���;��@�#\QњT�0��Z��*�-W��uW��|��!�x��.}L���2��R���F�����|��ׯ�޸q�OՎ��}lA�H`�57W����o�7>9���Ց�G�}'�ϗ4B��D$���us���oss����oNv��o����aw�5:r��l!�{�^��}�H�wii	���!�V��ݍ�z�7q��Ab1���߆�{��Lh=r�Z����`jqk6�c��e�׮���'N�ƍ�1lٶ]]hnk����͛�N�nuX�+��Lwv��IJ�Ɠ���ց�KE��~k��SG��N;�g�y��w�O}
�g�%���dC}=�§�����0�aH$���^�����ٿk��1��<y�SS8��s�U.aln�{����r��t6c��C>�F=W�*4Zҕ�oس��N�эy����-�L���>X�Nj���h$_���pz1nz����G?����D������ն��ǭ-�HkG�;s���D���`��ּ.���u8���i��!_��ȕ����aQj�5Qv�����V�Vv�t@�U٫�X"���3þf4G0�a�Tc~�����:M,\2_1�����QU$�wM#�rZ�f�tT��&���K��f��B���k�f�@C����2�P?�\Uuy������HM]��bS�|��x��E�I���4�ȴ	G�&�+b��>0L��gqЌ���W'31�տ�>�ў���P���0���s���qm+�Fc�
mTْ���#M̧b�e&�O��c~aV8m�K��^Ü7>J�ǋ�,���~�^���5#�I�\*�t$|p��3==����c�̑��%h�Ab�u�����ا_�#�ht��x�OB�я^@<GOW�7:3����~<���j���Kg�l=s�l���w�>����j��_E��M��C$��?܄<�Cܾ5����`qۃ-h�VQ˔�}Ro[�޽ގ.\[�F� ��}{qs��:q�9�h��}�Ql�{ cW�a|fV�Q�t�B�%t�����%�C�}1��	�f���i���E�i�ew���y��݁���x9q��a�W���p��p�,�����qt�C�|�$B'���Ž;v��ED�b���D�Ӆ��O���"_�Ѝ��Y�������w�h�9h3Q̏�`mK��9��
[7�rp?��z�#����3��G�&AS|"�Yb��J�X�]�V�u�C�>�+O_?r�H�O��m`,����j=�Vx;o\j���rKm"rHK���R�dZjX�v����&�,@��A�t^ח�78�� �&���hAg�r����vژ9E��L����jt�#X��N��4;�d��,�L�L6�kb ŉҍ�Jj�a�R}Y՚�\Uը�&A�nZ�@E��K=��:V,~���!�-S�a�~6��Q!�(B@G�bO�ƀNU�).%'];W:�E��4>fpX3+�L9�U�$j��L�C>srj���&A�T�6#S�@h�w�g���޸F]u(o�-�o�,̎1��9�43=�ťyML��Ƒ�L�$�%�/ �/��-����9;WЋªp��h��8	ܭ�V�k"����l������GGG�]�v��/#x�؁��Ȉ��?w���6:>~�X.5u���lׯ�@0����8s�b�<4Do�����?�o�:�ա��E+j%�oM'��a<��� ���.��t�Z1�|<��=�,�N"�xm4P]�Z�[1��xs�7oD3�K7n�܅$�(�-����cp�l p�#I`���w��̹�RE&do�1�(�EȠ�Z�"�oC� \��\3W������#�L)��`� I3Ξ;/�ן���)|����f|�W>�x�o�����C�v��BVn���ߏ��چr:#�Ʈ�FgO'�.�`���Gi�K�/BWsq�g�� L7T�z1O�p�j���t���4���!�;ɀ_��E�=�H0�*���NZ�p�}��o|#����6V�j[m����aX3	4Ӽ�Tʊ��+�%�Mb�v�L�BN�6x�8mu�U��5�RUEw�ae�)~���)�	/��f�MWN�1h*��Kq:�N,Ҽ�W�Qhu�Q�*�5��8"͈���rL
�M+�L2K�Ub�&K?��m�`�p�L�)`Ń�U��@<�,&ZZIT1)�P��:LB��j\Vf\��� ��P��W��`�5�D]��ƞzV����a̺���S�&�� ��Y�);I��].W���P(g���Q�(&�)>��r<�G�S[I;��0?�A�W�1�ilbR<<'��8����EGʤ��f
�I/�NE��h���v!�Ӧ�%%�*���)��hQ����^Z�ڣ�轹\��x<򃩩�ӽ���_&���4q:�ƅ�����#7o|�\��۸n�}~)�-.."�/`zf�DRU����X�V�[�ѱ[�dd[7�O��]�)��n
��G��o����z�D]A/օ���ʈ�����������pR6�_*c�΍�=�e��+�P-���#��]{����l��Fjj�0:��'`��=4��Q��V�i��,Ӡ�݌���Dv�V�6֒t=|�4	z��R)!$z��C_�xmm-ho��ȵl�=;�ƹ7���f9G�Í>?�7�.nݞ���߇��|9BD5��tC�N�y�BW�!�K�-a��i�Ȏܠ~�A3���N�Y&��ca�6����={
��I�t�"���dJ��?HǶ#U*�i��%�雺��������ݓC�?�*���V����� pyv�H2�Z��`q���0/F��uUFϤb�r��d�4�B\1��R���{�n ͌�T�_+�V��B(���Ų��!���ZJ���P
z��v ��M�U��]U�����/#S.��(�r�]��ҍ#M��ĥ�j5E�B�E�����0�c��?���Q����|�a�"������,ZC=\��X��ܟLeW�&&`2)3}������ƒMҙ�����8į����3�3iƚ�j�e}%fVG�פ����xӪU��]4��XX�"�QA<ڊ�Wߕ��	xK^U	
x=N!�3�e3a>����RMҾ���.G�V����_��r{���[�t����t��W�411|���:��o�����������������։�+>P�W�;`5�ź�.e117�/|]����9P��D}{mgZ;h���V��'P�HC��f��6Q�oZ�,�iB��0\vR��o�
;�,=� �K� Z��K�9/lJ �e�ۛ[`�cdh���C4�}H����`��	�W�c.��<����Q�dq���u�^8B~��p��]\+9��V�����@�?���><z�Ah�f�&�F�q����y�@8��ͫX�%�~�:�ٶ���t�}��q������y�D`M��
�w&���l%��h
\����a>���5��6�T��n/�����������|��?����J�^m���x��Bq[$��D"��2��E�ֶ0�b)虼R�:Uj˨	)�v/
Lq��j�$GE!�RUM���/�����FM-R��Dp�Y%�ĩ=o0�Z����\�L�� �Z�t����g\�g(�]��r�f�6��aF�t�X���w��QJ��K�S�R�΅?dh�*���k�E��6�#�!�j�*r:���&ӈ����+M;X�H���07�Q!�L-* #�s��dH�ԧ� ��ׄwT,U��Z1���=��
 ���A��6S	\�M��������R&��Y���jU�Uv�%���:��{�s�$���ŀ�v�(2�M�Y��KѪ`q��m���
�ң�X��/_~�
��E�x�M�~���/�/×�~���mnoi�ǣ\�~��3J@�������P3Fo�bnn!��lm-a�����S�(���gѺnk6�@y6�׾���8,t�hǖ�� O "�
��'�χBwg6nۈAڵ�,��`
�8ָ|hjn���+8G�6[�aǃ��tts��ʖi2I�����dK�TF�_@_G'�t�{��"1��d'oc~~�t�#���0�{5G��Btf� P�6nĽ��Q�t.+侹�E޻N��lV$��$n\�?��z@�oǦ&�A�*U�"I���"_(bdr
��<�;�}x~���iU��*A�>�� fT��Ү���_��*�T�j5��Ē�썺�ub��?����{�|2�;����V�j���7fҡ�X�D�4X�,zŨ`M[���&h��seQ�-�?�J�7buZD9���áˢ�zF6�E�n,r��BD慑�M��%*ũ:��XT�L� y�6
�p��BM�z�b*�C�@@gS m4��e�K��3<lnk��ǝ&�HR*'����
5�>8&"bKC�.�KM�)~������R&�3���4&hZ~V�k1��%�X�P�	�X�����W:O��fe�	h���.�T�	�c�;]��攍����Gr{<tL�T8[�XM%�>3�Z_v��(`Z��i����S�X���� ���qT���R���ة. �� �������<������K�*���yUqW��<����XbPh���w�O&7��
�����iӦ�/����hbͥW_}���W_�J:����jmvx<��[�0>z�x�&+�^���Z�;#~�29"R*�%^��ժ�r�ۆ�5!���z���������[o�p{AB��l~��ᛳF��঍ho�Aw�v�J}�lv'h4���>>�>m��G1_�!
!�Wx&��c>R�&�b��VK�nv���|���FD����� �P�N�fE8�Gdz[7@���S�ٝ۷�M;�a��ܜ�ن�m����s��/g�}�7|�<�_|�w���O}�,&3q��ݴ3���I��۶�N�*�/�=kp{|���\Nd�,0�׭(Z�(:�0­t�����t��GR�d�o��Ł��O<�؃3[�x"�]Zm��ӆ�~e"�`,W�tI�yS4y�a�y/��	�����.�"c� `"�Λ�.$o=�X��[��B��D��J�[�Y�t��t��7�ͺ"J��(�,�4�Yh>0�gmhK���n-D1´��fmD34������ص0h�*51�5� DӉ���3Z(c]CE~T�А(�$�4�8�'����T�fOꦚ��
��;Sv�^32ea�N�&�,1��I��S��˺PJ}�R,);�˚�Nq�&�	�����F��y�!�Yʆe�_M"{�J�G��Ua�uwF�Q��A#����IU߭T≾~}��Uȳ�J%z��y��z�0΀���e�t؅�V.�?�d-�s$<l4��H$���{�FGG/���~栉�r/��`��������ժ���vKssZ��N��!ܚ�ً�D�w)�F%��`af!.B��jV�J���6�GH��(t������Nh?[>��G�M֦0�a4��{h\�&�.,�R���8~�8��2IX��(^�wSV���4��>�0z�m Bn��A�.�G�¼�A���E�r�~� S$���<t����t���Mcvi�&�t�ɩ	�c�M�w�O�\%�I�[�aQ^I\i�7���-�ܺ�:�ݞ�[�5�S�p�7#��N_qO �d"=�G��WX�f���(�s�("���ٗ����� �\�j��L)��N[,�g6l����'�qQ���?Xm�m��t[=[��^J��m�X*�v�T��3�ƹ�hC(�l�0�nC�P��%)����I����R�j��5K*j��Ԓ�����9{e5�RBd��,��Ej�{$
�і�����ݢ*��:�;�J���h��.�1Oa�����6���s�Av��͉J�" G�LC�T�V�)�S���j(�/�ME������;�Lu���[���A��DgD�AW�%N��ue�lz�5�LԹ)�b�kcK*&Ls?��;���S�������qT�A�9�	�+�
h�L{�e}&�q��!� �@T�@EQ�4,�кy�ֆ�KE�^uu�{�Z�p��W���uIֳy�����@���`��ž�]��">{�LF��S�\i� Te/�����oG"���fS�Ξ=���������(���)hJNM�^y�{��=}����3�;�Π��У�˸{�.<x�~�ŏONɎ���򥤓qz$��ފ��
�ˊ�M��Ê���}�S�K�T��W��6�����^�x(�Srs�:1�{l�a��g�41%f��x���\Ӆ��[��,��h`�Ϗ|,I���{��ݟ��]��7�R�Fo�
��n�%]��v����iS$��Yl߶�>�
Y�LOa>��~�N��|�ߵ�K]����;�&@u��)l�D@��c-XK�'?~���;��^��s'Z��-[r���&�pu���x��ױs�:��wN��}�n���A7����	oktw B7O�R)G�b�zE���u�����{�l>r�����Xm�m��t�d2�'�'�-eâ��ht_��^�BܪT�A�xҐ+WբO_��r=g��@��)(6�5jv������b�j:^Q���aF.d��	8�Yb�����E����E��J�3��^PA��F��%��Gya�m�)��\�S#`U��@�3ȩ+�hK	��)�m�n�hfe�nV�A"@���+�9I�	Ph�~VRsⵧ4jfƞd�ˠ�+��pV��
�)� NJ"�A�R�~�>�����d�2�3��� T����]s:��M�u2�Ԩ:/3�WkD�ѥ�2}�4���eZ�Jj�e~]MK������`������[��r񨣱R(Va' ���N�A(�,�X���EW��]EU���q��iwh�@�V��ה˕�����x�8���n�::88�yO���@����;�x�_;���/gәu-����������s7�sf�'q��	�ݷ_���Ȗr�2rC��W.� �����Foo'-�	B~�g��������ٳ�����������Aj	J�լ���(�� \k{��A�?,R g/�̍k�lEyj[�zq��I!�ݵ�7������/�lj�3a��h�D��z֯G'�15%�h]����]�~,��A��DT�I?-�%D3i�!�<�%5��96*���@#��OON �8/�0ݘA�7�����A9����a�>71E%�����>}��{�v��2�����������iӂ8M�s٬+��b���7o��������O�5m�{�����( ����J5WEw!�����X����%]��&Ds�6��`a���Q��\A��G��G����灝�>;-к�D�T�5)��٤�q���&Zò���hJ���e��`��2#l�]aaGO6otG�MW�6��r�\�~m�����m���^-J:�ʕhX�38�`�C�H ���c����J��/]��RXtj,˚Lwڐ���e�#%��8O8M��(����uS��nڥ��P���L�����;L��`.�W��U��~�M���� ��~�(�ӐhD�Xˊ����L�um��N�����M�U7�t�a5���w�P��3W	5��3�I)EhB�O���|�@ #��,|�v=�|I:�#q5إ���K���A��s���z�֝��>S.vr��
�̳���+���?���v�t��Y���������I���)K�=]z��Z�:�]Ѻ50hwr}�*������p����/���!&gf��ڎ��v�<<p���\�Å`s��b�I1,��q��'�	0N �<�زm�f\�=BH�}�ܵZ���/�^E_g���.|�����/��܃�c'�4�����?8�k6���^�y3@*�J( �����>�sta��{���	�eG)����%������:���l���!�߃*��|��[7.a��n�W�_DO{'6�ۀ����qn�!�M��]��͊�6l��N\~���y�+���T�A�,_*�ĉ��,n�=�ӎ4Ewe<��,&�����\?�������%ʆ����V�j��kU�^/�k�rMbsz���6���m4g�	4)`ĕW�.�hѬ6Z�8�/B>A�6`�!ڔ���%a���W��R��7<��|��mM  ��u�<_1t��m0�P]]��M�4��E*��]>�h�Ȥ�Y�!Fsd8�A����奅9ϙD�q���V��D�t�2)��&�a�g+3��H�i
\-�EbE,���Q!IC�K�ʢd����r����)P���M H@� ":E�Ү	Ȉ҆�� 8�~�OKD� G����B�cY@����k�[���r���2.ՍM2=�����S������hZ�D��D�8�ȟ%ZTJ7����<�E�̜�������ȸ����k/���%>ӬX-��߯�J%'��B��;??�`�f}7��<O����#x�gM�]�z�j�o�y`x��b6�nz��u��nBOg��`��J0��(�޷� ff0|�*��b릍x��G�އ'j
#���@k��L fl~c7���"�)��oB��rmfiG��J�ji�Rv�]��%�nw?p����.�������a���������_�����qt�ۈ�Lq��X6��T;>�t�w +������>���,f&�16:�'�x�k�e��hR��0B�i��ņ/�$+�84���]p���yc��|ML!R8�v���{�c���&H}�M;N��;0��i�/�L!��cpYh��P�����EA�"�ւ��4�-��V[}.�'2�y������^_�q��G~�k����m����MsX*q��y̰�����r�H��r����~�׫Jǋ�X�ʕYF���U�dv�� @*W�ŻH��"��B^�"V� �R�H�f�e��(��.�e�z�(���X�M@���5��ӣ[L�JM@�n0���B�.�ª�}t]vŜ���b�d�@��^rzM��6M�YD��*�H6s�_�0���&F��cj�6xNfuL��FL�aD|'�jX�(�mM"Y6S�@3+��O�7S��N�&�$�^x҅�L&�o�QAv}�~b���>�>H�5�_�Ћ�Z �i����&�kX�U��A�.�G"S�O� ������ �C%�D���N���ȓ�M1hn���L��aA._���mx	4����4�X���r�ř�&��K�$ _6͕��.;���kؒ�凪�ǲY�w:��ˑH�&m�3�9i?u���"�h����_~���w���=��鰶����tw���A��ᴜ�v>�C�RY�nEx0��K/��L.�f��vmۊ�d�t
}�=�[0r�&������]�N��̏���I�ba�i4�H�s�^�΍��Y���?�ɋWhnqa���x�Q�Ȣ%) ��`G�<�ۻq�ӟ����P�GY�w� ���qt����M��.\f�*>�駰}�v�5-�ϊ+y����b���v��O>��Aj�I-/7���Y4�5��-������0qus��ܲs+�{;q��Q���˰�N�M��儫T�%��Y�r~vS�м^ĳ)d]yB�����7H���H�V^�s�t�V*_z+��yl�Ν�~uǎ�Ƒ�ն�V�ϴmoo�=;<�_�S��o�+�.XH�Fs����h�����׊l� ��2-XVN٭�f��H��Q��{�d�y��\��`犺�&�t�Z�^q��pz��>��U�
�\�_Q�il��!5�l���B�b.'�:!���h޳���P�;Q�� ���T�+�%:��vX��i���΀�mo�
pNSѡ�>L���a��e���
����T~�u�"��0f����$�YT�E��P\&�T��E�0�t:+&�4c��rŌ@9U�-�/�����.b�6$�#��)B��8*Ť�J��ꬸn�#zV[�����+�k3#V�2��t��O�����@�R)�Kt�O�yO�2u:�r�TZ�3�=��X����\e�x7m�+̳�摡��U�,c@�I@ ]��^��-�fdd�P(gbb�e��;�?����*h�/�z���M�N�����'�*���Ͷ�뇴��N�8Z�����.�9Ku���nF���L�	 |�n����>z333p��ްfH�EN�=��O���]c�7��s �~��{���km�k*�����-�J��o��##ױu�N,޸�o^�}��[Kϧp��	L�̃F �3Kx�՟�������?�������L��_��f�B�M��i�&��ਪ�ѩ'�o�^t��Cnc��3't5q��`�������; 11;���i\��}�a͆5�z��~�Eu�Hu�{z�n�!~�2a���+݀�B���[Z�jn���q�s�:,F1��,�SSI#�c{���=p�+��I�ȑگa�����/Վl�_xu4���Xbr|)��d��ͭ�|2�k����%�!
����.G38�S���H�9��9
Pg�i����ePq����N�V)�ar8W�U��*��|�ќ�H"��I��F �mW���� Ut�d����(S+Un:&[�� ��V��N�~O��%:�r��.%�p�|h3��s H��RΣV�Ӻ]�c�uy��CpǑ�f��T�N3|I�Aٶp[6!i��+�9!��̀�0RY/E���L��̍Z!����N	bҚļ ��2�Gn��D��,����d���&�KT'_Ns�ػO|�LqQ�e����3m�M�N��[��4^ը�q�{f��b�w� �rS�T�Iʏ��@�c�i1Hͼ�1�c�t{��%����� B?�n�d�JE���H`pb��A�]���V�F}��������O�X;�N�_M�Rp&>����Xsiz�F�����ϝ=�㋑=v����=���A�1G�����>�ѥ#	�r�U}{��ηJ��s�ׯaz|
;��"�����0�]F:����资~+4�^�HΘ-Kr4�rsq�X*�E?��֡��#cSط};ʅ2ݘUlش�Ο���qLǢ�d��>�=�V,D"x�'o���/����]*4ḽ�x;X���:]\z{��	�D���&�,���"��LB�effi�p�wM/lN��f|�+i'`�a���LO�F2����Q�������_�%�3�q��ͰCHM�l��;K���4ir�]�p�!�@7���� �9�H�t-,F�����p��������,���*V�j[m���Ps�]�x�y���b��L�3�f���|.���b�m*�м)�7��su6�t2)�$nZ�d��4��;�����6�p���׎��+"¢,��%��+��/�a��J�����b���L�� ��Via�L�i ��4��H�D��%��Ud��;�ؖ,��+� r�<2�"�\vt�y6Y	<�_+
X2j� �	i�I�b��)�r��N��WD(��R��Yr	����Gx@u��R�J�D������0(0�sD'�@�fS�9.d��d���V�Q�WDB�/��4�,���^<�(VBt��H�f�}4zT��EhZ�S�@ �� r� +�R�(�<�仯�/�y)�D2��1���$�$��pԉ?�Z�
Y��Q���μ.�S��阾j�zw<��I��H*�~�����.�����1k�d�4::�x�wv_:w��cccOԪ�5�����[�l�Ĩ;�֊��f�]nB�E�r9���îm�y������g��܉����m�lp��5�hw¡�MC롍�a>�J2�Ն��I4��hi�T.IL唙d]��ä�p|�1���0�0��ÆŅThgK�Q��K������I҆�����;�`ȇO<�8�{�a�:�90��r�Ϝ@�� >q�q�~��ב����$`g���\4��)�n8�)�i�c@p�D�J�2n���)�������'��\}�=|�O��?8�YחR��rh��2���䖫�P���G{s�m�	�:	���#�\=^ȧӥ�Bo�l?p���O|�֞={*Xm�m�}��aM��3�B�?u{��X4�ɥt�~��X�t6g݊T<�۴`9�>[Ze���8m:��xq$����i��în��Y$"���BqQ^�"������م㒠9�-:Z�����J�Z����ܡsZЮ�S��ݨ����_���������P�%H"QU�2�,�P�%׮x�l����М=9���E�Z�fz��tK��m�r2�Dˎ��T�ES�9%P���M��e�H�h7��@�rzo9�dQ!�R[M�9c�����V!pS�Y%����Z�%����Ze��ҙ,4)�#�J\���zN|j*�(�GS)��;%A�\ig���w���Z�@d#�|+��[}%���I+�����`�&ѱ�X��"9s��;*Һ�qL�Pd�晼���~�@/s�A�ƙR�gS�^[�T��_&�����}������1j�$�ĞqN�̥˗~=Y��t8}��� ����N��v�����@H1�sv�d�y7c�)>S�����(�;��������V��/^��/"[(��G��D
���B�n��c�P�g������a2�����]���^|�MLG#8s���q��*1>&�%�|�q�u`�p��uDg��F��^{G��;�d�9��D����Nn�@�F�P&�F=~�!�[�;u�&?��֢nA(�yz'��<�;�$��Kg��G�bd�l���Y��+����G���S�����y�L��`�����6enK�P��Qq{P$���<�J��[(���[^�������WԴ����ն�~ٚy�&��k�3�s7�^ZJ澜�򇼆֚�y-�B�D�L��Vh��xݢ��dp�h���x!������ps<.JY3I��^4s/m8��M�Z>�Bl)�b./�a;m>�;-�J*.���j9��\I��!��4���!�Б�	⅗ � ��Ȅ��hTJ���5Z�+*�
��.Qz�O��O]�J�����N�N���q`R�z#�gF�TDJ �ֈN5�Q���'e6EE�Ֆ��|�
�h���S�)=#Z+lL|'�Q!��)=��&���J�Gc�T,���;@��H)�XZE�(h�B��;=���cs%��b��R���E��ajQ)��̗^�M�l�6T��l�|�\!��̝�u8_,���R�%�pz^p��Tv-�s
�{J�b�Q��.--�����,>&������}�FF6����_��,ud����z{{�f��O�l]]]��hw��넲��Q��ĵ8���qangN��ｇ��9�6�0���勗зv ;�����Q|�{�����O~
�H��Eė��"����u
�s��%q�l���%���_�]AU�|{�vI�2���/d1;��/�vcώ��������o��_��j	��;� �.�)!�L�ȯ|[i`�����:���>�ڱ����.`av�c��{�R�W�I�Y�b������:x�Vtu��q��N{�>�F'�M��O�kv���A۫T��	�J��F;{0[K4m9��b��f��l~�p9�شk�sO��?9���%����ն�V��Oۣi����S��K����Ǟ��-�6���d��e�Hg�)�\�m�|43O&[�#C��^*J�����^6�bEU��0�PsA''�h�4Ӽ�Ϧ�N�%z��E��7��`/;N��m�_T��K�ԗ����+,��K<Wfe���q�@�8�e�9;��u:C��J�Y��F�n�t��%��E7�ϖCHB�V����,G�V"Rf��?�a���i@�Fz��I��`C�VVM�h���Z�"i�Ȃ���nA�yd5+*���p�ք[ėUa�++�9Y$"ƕij�\�V_M���ؖ�G@Q�N.�Y�)p�,E Uz�'XQQo��[�[��1�W҂����_��cf��-V�>�3��`n\Ss�WlR�r�����E��?M�bk#�kV���h4�o�O�������Q��/�ҥKgO�����O,.��r�4w0��0�v-\/�Tu�;�Мҗ �j���DU�y�ϝ��3�p��Y��It�w`ӆuhooE�^O�7o�z���v��8��^�����X/��0�|�[6�C��x2?��]��z:�Wn㶭�i���/ ���O�w��O�FjOO/��g��o~Q%�����c}G���/⍓bx~	E�����t��54u�16>����0}���w��nEkg7Z�;��s�R[ \}W���]�/����&
�� d>�󯿎W��&F�!��O��d�����VMH�6���l낍���Q+����,�k�T&�,��u㕾-[>|��G�L��b�������>�L�\��3�Sg�#wO�s�rj����͕��$�J�<���dNfp���S�Q��)�<���W�P�N����J\��\�����O;�L��`[���Tq��C�ϥ�l��G��H�\-�|�F8h�������'Xt������� )�
������4Y6�e1N�k�*26/�z4zFUɩ����vS�)if��P-�h@��6�XI��!��9f� 7&x7lQ��P��Ջ2�����Y���@]E�8�e�JH]$t�j��E�G�EAk�e�T�;'m�k�6��)�;@�@�� �so��+Ud�ϯ��ldDuQ�����\7ySXN
��U�R,)��M���j�*�bE��u�h�*B�>��.�V�\,4�r�#�`�}�ُCv���)�D�����O糹0�L֖�;wl��u�}wtJ��N�˥�r��C��f��ݸ�S38�4��{�3�b3�c��%��D2_0���nttw�RLL��ޅ����+�z��� �����Y\DKs k�X<��t.���5غs6n�.Bk���p��rsKqq�LZ$�ݶ,�'j�
����p�/�������t
)�QY]	)�XI�&���O"�\�]�9��o��ͩy���!�mߎΡ~�	8�a�B��-봢J���j5��ܭ1\y�}�}�'��v\����A�'ʡ�
���@�L���	N�8t��X,dR�=;�I�-��l޽�խ[7����/���V�j�k�2�Y�xkm4�����fc_rT�G��MM�h6��4����p�8����fw��{�{����)�X�Ϋ�\W���b����$ZC!��t���\&�mL����h�(��>�nl���92b�T4�2XZT��R�eQ�nC�	�R�t
no��T%'K���u��A�P�"F��@�@�T�!G�Hɱf�Pi˶#w
]
��L`c:�:�bn��>-g���W2�r�I3	�ʤo0Y�7�,�����! �(�(���Y�f���sTmv*�$���J�UVD0�L��M1M��iD�Q�e��9��4�ˀf��ZYyL�h�ߐ4�K�XL�U��L3,��%�u��/I�����q��wus:T����h��4O?5����z�%z������AS>mkj
���͛��v�zStqI[;؏~)͡ !JZ�Z�m
��#��p��و��#�+S\�^��ӧN�ʕ+�S�4�����uĄC�߇ �5�]����E������h�1z�&6nٌ�P �����*_F���T�C�>����ctbv1���	����x����M�$�������c1��N(��Ս�p+�tgO�Ca~Ί!J��t��휣u��װ�@��ĵ�q��8�s7��iܤ�^�>�ĵ����=�S	K)��hwfJ�ߋ�(��(
�K�NO��4G>�^}�]F�d~�&�&e�� ���D�e�����Xl�n�}g���?ܻg���#G
Xm�m��B�#J�p���˽����M,�~e6]��[��rՒ-��O!N�)�Ԃ�p|Mʹ��1�I	y��,mrY��&�k���4r9����Rh����#��\*I�ɢ���<n�J�Ѓ%
%��8��gL�� �0�%^(�\�g�H�q�JP�ƶ/N�9e��0b^��À�9c+f��+�5Mj�Uonjf�N ���*�����3�x��a�~��^6�Z+.�,JRᎾ��R�(\}��ݤr�G��4u��72�(G�jֺD���A�nF2y����& �_�ڄ����� '�
^�H��F�K��r���?W�q��fJp�L9M7�4M/@���޵  5�IDAT|��<��u�m�e�Ò��B6v��&�1��{���Z�~y���(�.U�UN�itnzt@n?G��XԷ�j�Cjw�u�6M|GGZ��M �%^����7���k(��f���M�9uϝ��¢�w[�:��o@T��Bi�G�!��Cr���?����d�߸�=��% ��[o�pۑaB"��9jj����i�v��9>�ҏq��e�>�8y�,ff����isHP��t=N'r���Rp�8|4I��itx�[l�7�MDi��97�.+���-%�����k���-��fށ���7\G��38v��Ma��+JIskz[�q��Ugf���N�w�����_�*�]b[w<�7%��r4xc4IŲ�J*_����޵k�۳w���~�+��ն�V�?o3��»�����o�-<<I}v)ol���D�f�9%YD>���fڠ2���mEZ�8�g���E�9ę�:-�N���A�Ls�t$&��l��E�dws�Dcb���{YP��m�/ �^��]"-����VI\@���I�ge�\��u��a�5�����w�nn]7��p!���bd�s�Re���roHW%����l]7A����Q�
��l�r�@����ҭI�">k6�.p���j�(��:!� �hM�n���i�]�y石�}���]j�����18��8N�I���)�����|I2��j*U3UY<�L����`�l����6ZR�z������}�sn� Nr��H���K��v��s��?�����x�\o*Qh�5m��t,�XW�L����NEL�aG��;�5��zn��w�>�ڱ�S���O��{�5F����,P�X�Q7�ؒoW#nnT��6�������q�uD�n*N��nC�/g����Q9B���[�t&�s��ɽ�T��tA׿IU�}�F]-�ZMlCKK�l>�+
�@GG�888����jK����q�x���7�Z��T(¥���k����K\@u1��;0��롳�	�X���i�D\���O���D�yv��`��-p��Sp��Y�w���۶o����)��3�<O��Gp�����7���^�~M\�7,�䰝��u�t�V��:7�l�}�g����S�Lн86
�l"��"Ԍ:?P�d�	��ѣ��&��m��p |�)����C/��®u�`�a�{@̤ؕXܼ����W����AGٚ��?�pG�ض��Ud�Gg��JŚ+���m�������C_�ڬ���'�S	��/�^w��zko\�^88�+=0�-�-hN��~Bl�_Y\�v.ÑJ�D�a?�r^�͇���9zƙ���b@�)1\��W�P�T!C��c�6~^/�* T�	ƀX8v~��*FC�" w�f�U�gފ�Y�.|QO(Ll(V�rN��N���}�΄P`���Ũ"�_-�_��[��+��.��HVs��E���V�2��c�9[�x��m�����
��߫��<]��K�jĨV��^��J���r˥�W���0A%cy
�t�nzW5q���jw!vݹ�H�׽&�#SPHbǴ��1���ܿ������Go���Z�γ"nt��cnPH9�[���l��`��i�G|�~�y���z�N��x���E��5'��\;�+��2��:��ŀ����c6�b�x�t�]/%�Wcϛwz����i:���P$�@7����3�Ln�d��h�oҴL޵�i�3gށ�Ǐ;�O�b>�XB�� ���J$!�HA,��V�p�O�;7�o�?9~���+���zŀ���ض}���Fa?|����,� v�ٕU�X?��2]��!(�Ws�xx�B0��>��n����	7v��^�Fv �,.B�T��TJ�ͯ�Af<E�`���Q���G �R��K�L���]{�?g`�T�{��f����흐��Kg�0ŭB���� H�( ��L0��l��kf!�X������]?޹g���]�f��ҿ#kJ� \
v~;}T��)�lt6���b�������8����jl�]HV���]�i>�#��iXkԑLs�Sc�Qe�5��*�~LvQ��֡���+�2�gҐI� 	���g�l!��C<z���L|��9�i'0t�`�G�G'T4���;�KLT�L���hʄ�3���|&E|_^}f���c�R�҅�����+�ʝ�e���^`�m�G[/~����"ݨ�\�`$� P ����l���%xu6<M��#��e�Iy+O~{S����eMLL�X��_/r�^����>��.�D/����\�Y3�����Z�P�E.j$G��%��j
^�dbۿ���=���
*�pM��7
��HDdAP��R�ln��x"�q�:W�qK�l�paW����{�:��L
=I���$]�6�!u�����c�{>ñV;�4�͟#MnZқ�'�<�#�����FM^�ߋl#�ľ��n�?�6��nޤ�J��T߼�v���"���_�)d��J�"�R)߶-[��!�L1��D[w�m�W�Ou�0d+cӂ�rN�<	�z�g,��0;;:�=�vJ����D�=��2�BQ�l넥l�R �g��e���h4�r|���o�f/�h�;���R����Q$��f�{��~Hu��F&bT&���-�N(�
LD�~���j����_:�:�RD�8��%87r�����+��]���98��a����.�ɶE(*{�=��A����r��P�M6l8�ȴ=s���Ǿ����"4gA�O``m������'ҳ�ό�j_X����l3�Wem
.�!K��f�vd@�[Pf�;'�/�-l/r�5�GPx�A�R���9�T0��]!���&Z�����/�qQ�cG�䆛�Z	4K�QY	B�-�82E`뀪� `����ȑ��of���m|Ϟ��;����U��j��`����^i
k�ܚ ��� {~��-�6��R�g�a�C�"DM��Sdύ��&��~>E�.���\`�����Z\\�Ζ�k��� ��~�<֌(��!x>Q��z;�
(���y���c�Fg���.�p�x=���ډ�Fu�)�'>��Pt2m^���;q�Ղq�aZ-��q�Y�v�-Í�5�8��r���v{%iM0�Bpc��6��W�m��R����fa�Ɵ[���՚0Ӫ�����^2)ا�;X�썍�ː�%��6��Ƹ�Yiv�\�r�9|��t�»���`G#e˖��-�����*�qvu��������:~h� S哠v�31>���7�|.\8gE����{v��۽7�I$�ͺ&�>}��O����o��ه�����![��+#r��Vs���k�u�T�bb"�%�h��v`�	�E�������S�Q��������?��?��Ϗ@(�ev�,&�R�p��9ф�MC���\����<��a����\���N���������Ad��Uv��U{�T��x!�������|�w���y�_��? � �V�j�Fvٙ��-�zzj��ѕ�ϭ�澸��م^ey�WV �h�D�R8�	kv>�����*�-��(�
����E��K���+�vnG�l��s��(iy^��z]|l�F�0�_�c]��%���ė��.
��ƶ�K���K��{���Uc_F���'�"�������/���fò�A�)~U��?�'�q�V��i-9�~Sx�wǴ���&���b�����Owv�<<8����t���2c���/�������#�1�.��^G����-��`a5�×YW���Ļ��ʇ��0�[^��������;�����u%יհ�_�ݵ�����C��f|F��-<#M[�R��{�y�IU�׆o��3��s�x��Ov������?
&�ơ� 6�#7�xO$�)J��p4�Twww�>�#8*l��ٷoXv�߬Z��JM:r�U�ԩ�Av se���)lݺU����$o}Ţq���Á���歑x�����Q���G^�So�s��a��rv��Qڱs��=�}�@��WU�%�R7S�"F�N�<o�q>���w���7���C���Č�����Fy3%~@P�d�e����pU�^6��l��2(�a��.$���$��A;�bє-_��Pء	U�7�ª�xgaڋнqmi����¹s��믂�W`���ɩhkoc�"J�6v�Ǩ5j����,�W��oݶw�Oz�m�>x��{��@�a��������ً����׮,�~k�Qo�|�n
P\Y�*v��R�i�������T���cCw�	�F�leU�1�Q��)�-��{��o�Ck�:��`W���G@����T�{Nӹ_.�a�u������Z��bJ���t��ssso�+�G����՚���X���}�J*/�VC!^o�hh��,�$�.�M�l�e��Ic�d�;[�����ø�G�:8S�Վ�s�ߨ�K_b"f{\����Fq��=���^K��l�W��]�a1���<qg�6}w~��4ǥ����/�8�Es�2�q��#T9Zu����Ew�����մ��Ό��KZk�X�/ʮ�ێ(���ncX���۶A��ۼY7�Lc��U��O3�4r=eU~�1*�`̳��%G�K�B��ٳ�;�O�����9�;:�h����u@,�p[�8����l��q��\x^}�8�w	�G�έ��Zڴ���Jo���73��]��jß������9a�����q���}�����O��ǰT*���=�$�9J��7BgW��">	ۏ�H�
���NL)oض�}�Q�+�o���`��y�����qG��P���U?F���
L�h� ���O��y~l�|��a��`׶��}h�������V���P*��M[��q��gi>A%���rm8�Ĵ3җn�����o�JJ���;�\]�\nr�*/�M[ܤ�d&>p�C|~*�"/A��e\��6&���V5�+�b��oU���6/x��oK����,()n�)�؉�^w����M�Cߵ�c��}5k��������7�y�+�B��Z������Ý7��!Q2y�E������8<�%y�\��`rUZ�d���'��� B�}9���\�9}��|���z��e۲6Y��Cr�]w�9�d��<I�?��l��Nq���U�����cD�p�߱��[��Kq@�0m���c�{5�9�[4븚��%��>�@lqWL�gv\�E�l�,gm
���B!`"	��y&�m\L~O��ko֜�������L�	��#~遽��՗�έ���Y?�Pua~��u���͛����?
	�?Qt������b{+n�F�
2ۈX0�t�e���c#��<�;v��m[����Q&�^$��o��V�]X�[���Gc�i���	�2	g�yv���9p&����X� �h��ƙ�����^^1���-Q��U�n��c����͛�����ݝ0:7�ǫ���1�`*:K+ D��¼v	]wMv ᜺g_9�J�R��!���5��{Y&޲V�6��8J&�ܴg�w�q�Ϸ�qG��)	��V<�+ԱN��������-e??Y(��ֻ>�_�-W��<W�\v	bLe�:!��_�R����!�E?��Y&�t��h�XD��|�/�8�QT?D>^�\�W��[�
�1wXp 砙e#e�o��%���?^��ԙ��	��{����[����"X�XzL7�ƒ���L�f��Y��lnrl�6-g1}�����ݩ��
���e��}cny�B���Z�~�c�;I�I��:o���j�qĵ�\ow���]���u�"	h%��q�%r�#p/$�/�Ĕ�չ@�-W�� jF{�ƨI�K��0	�b���D&�����h��L�o_n!!+^����SD>OE��cT�7��p�)���:�M����gW4�������w�=���UlkkcZ&@?&�H\����9N� U���R ��N��C�_��'OB}���`�MNo_!�J������7�r��k�Y&�����¶��u��m���~��w�СC������[�O�@Gw8� >[���B-� s�'�<"�p�8Zp�[5v�.V��i05;�^��N �bbǛ�����F871	g��a����T����d�'���qȄ"|ho[2ů\p����/j:�kc�R����gn���3��r˅��{IpgMA\S����+�����#�잋K_^���)�eS�]���
h��3�'`��*���Ν��AO:��g+n������/���"_ ��[��)��f;�JX6!��7FSO�w�&?��������r�ʩ�B��B�xs��x�2����B?�hkM�#�w��&�6'�������~�+���e^
9�Z�}�T�?S\Y��Z����Yq"L�x�ܰz!��$�)7�L�n9��8�;�W�f���V��\�-L�`��-x�v&Zoq� �����	���F��*\pnM�W�.�%��s/ޖy$֐�|�s2Lnn�]s���u^����`�G�*tL�=wh���B�W���k�>v3���QD��R�'��}�ʕ����B:��vtvg�ѰK��<�;dW�ͼ17�m;59	'���CG^�+WF�N& �@�wyhh�d����A�"�gW�p��0��'*�ehxc����瞅���C�i�&���`~~�;�c-�!���^+�":S��DCn��cl��DL�]�PP� S�K��@Y�A�/1v0Fk5���!�#�� ��AM���&<��z�}L����]coMלR�a�Ɯ-^�tӶ﮿������E���8�!sl�z��x��pgv�����-��;W1S���(��xB�4����@�0� �j�����PҬ��*/x�} ���kUy7��r�!,Z��2�:;;U3��<������0-�]dѪ������0W��Q����l����qI�%���t�PVT�t<�������>����9�Ğ���6�bq�n&,��E{EA���������δ��:`�-n���=��#�\�'WX� \�	V>�ΫMr�:QpI\d��a�<��f͂튢��7 �Yk�*�`���������b1�}����ׄ��o�E�<5���f����P�G���:�#M^�+cccg�t��w����PUw�z�AGw{�m�VC�T(���#���G��ɷa9��[�w��۶m3����@8�g�������������w+�F���_ݰck�~Y���ކS�[n��vX���g4�f*��x�G�#�$~�ٕ��>��ׯgɂ���@2ؕV�/���K�����o����剉+Peq�ov����`�w4�W[����>!�p����-?ںs�K}t��A�^�	�3/� ��|i�x߻�K]ɗ�`�[��FJ�%�CО�A�P��b��)�D_� z�`�.M7@�� �Ӱ����ͅ�@�hU **�x�7uD����gQ.�����=z�l4>Wo��6c�e�~�fL�]���d{����m;-�ݽׂ������O�j֋�j�K�F�L��d�#�:�NX��4G���EY-o�/x�L�t����^���+b�I�@��BoY��^�h���3���f�� ��yMnṰ�z&�������뜣l�E�%�n�����G����_"5{-�HD�}Ж�nH��}�����r�Ϲ�jc�����Sp��7`r|��w��{��CO�F(|;������3����o=��sF�f�*7���u㑛��U-I�������f�ɀ
2�,5*c/�ʄ�Qg|I� ۑm��F�`y�ҷvtA[:�3SP���0!�
,��z�:�ݹ�	Xa'
�=I&�����	��0?���"����%[�w���Ԟ��v�����֭�]�� �[�'O8��=��#����\|t��o\�t��.͒	s�,�Kaعq��`��i��8�����ϼF�f���<��)!�� �@�'��yw*x�W���������R��L�\��FH�}�`8p�/IS7n��*.h���������ј?R.�V��v�N˲�f��=^HWl�'�ӌ85���!W�X^��Y�O�$���n�IB�s�u�F��ݹx����k�P<y��r֌;���ڼ=���(��B�@��p�{w7���^�R<{�z�x?�hz?���<�6�lk�eJr@�$�X���S���K/�;�΀Ķq:���;w��͛,��+$�����M���D�9M�0�V�R/#�m���ק�ܡ���!�o�����<�<�ه�M�d	�8@0���0��+U�?��(�J
���*>���Y����<h(�d���� �bap�)�h�0�>��sˋv�֨ɪzi`�����{֯�#� ��=�����:��lg��ř�GǗ���c�$�S��<LNNB@� �	�]��V�󺚐�x�%��X�v#�ڏ�B��#X�X&������G�kO���Ľݘ��q��o��V������������\�7�P��0�n&(dUT��#y�����kj�]�#�H�(�5��:�-K�f�4�`��O�Vá��,	;
��nM����4,�*� w���V���F�X���$�q�4�>Y�7P�{�z 8�ױq�5MuvY1ʶ�2���W.^��;v����l�7�|����[���ؓ�L��tz��*|��B�T����i*�sǶ-
�*PU�0}�m��sj�;L7$��ep5�5�:�����&���vb��=Jʹ,w�1���X,�vrHuwBM�!�nH�$���L��k�9��T�m{�k��s{o���m�w]���;:� n(nI	x
<���ɋ��g/Ng�4bUo�"��l�	�t� ��@�`_Da�0[�ׇ��N��ԝi���
[Ѭ��t"t��*U�^j�u���g�NM՗�{���o5��M�:�P	��Ќ6���_��iH�L��ܸ��[´�íP��� ����y����ټ����iF��h�5ŴPD��$n"�6������~��(��W)��^��
&[��+�P�Ɏ��Y���֢ɮ��:�6n���:q�8LOM1E�6l�`���7C�Ћ=}o��i�̯�'��iG�w�^Ku%�;�o��P.F�l�J��#��t�r�w�X���}�>AZeh�:T�� �C�V�S,4	K�x]V��D�}8���"C���e��˹�e��?<���}��2������eA��'A�ؠx��h2zj]��{dz�	�p���,��299sK����I�e�rbI[u}x�Ҙ`�2!�D�',W�۟��H�'ym٥K�������]�>�~�����"���Y�
��|��9 ��B�7='�)"5�E���.a����<��Ǩ �T�r�B	�SΧ���(����h8½���p�)w��P��O��RG����k-���_ZZ�*�L
���x'[0t��ۧ���f������֋�R�(�20��v�3#W�UC��D&K�
�{n�rRh�?�A�R���AE�Z��bEU��X�^�3�F��.5�9�Dw77{s~��$(05�/V��r�Q��K���o��y�O������M�"o� >Ax��hS�8���L셑�هgK��.ה�r�.`W����T
:�)DS FtvC�=�,��uNՆ��׆:���y��~�4�5[�~422�r���t�V��i��{;��h�)4�J�z%7}&5c�����r~7{t�Qx�aY`Ȧg�ď_uSg&��6�j.���-�4����ر��C/	��)L�9�ɍD1��[o`STB� ئ�_�,�'c��wٱr]v�]�5M����ېeF�Qg�Ν����T&�z2�=�i��ר3������l�xwBR~ۧ���_{�z�<�H��ހ(H����A  C�L<�
�5&�0����{v0�X*��OW$��5��Rɖʧ�m�ݴg�O���{����A�'Ϧ`�ݞx�X|qv�p��|�k��͋u3=_�)�SUX.W�=��t8�pD4@�eقZf���@G�:�+@��x�,��|dd�h�R��R*}�0����R�$q���A����s����i4g�6�wȹ���t=$��n�<���P�������%a)��l,"7�=��'r�C����sFBA�EB|�/F�|8��2��h�^H$������1�<�$��9@?����q|b�Z.�/������o��X!-7ZLOO���|qC:����Tn��}�4�0��!��*�6�2�� D�������z,��H�9��y�,��r�:,.�T�k��m����s��m�=z�m�}��"Ač��X���p(�83�T�k��xxd>w�L��5*07�CE�C=�t(I_�Pջb�c�Ɏ��o�M�6���y�ҥK#�j�X���Ѝ�m��@�'ITV�����fmS���闈�XXP�.�"F���p��ç�%Z �������`>r��Q��&���֬�*�>.�LC�F��7��2#�
�^��,�\4���a������?P���{6�L�����Ją��sְ���u}�r��M��}�C�]^��s�\5�WAg"��h���W�Sa")�����h-���!>-zba�)յ"��8���������A|���FCF�x�Z���џI<zq>����٢��8��<�@L�����Md���;rݶ�_�x�����'BWbo��+w�����4m�(XaUU��������[��=�u�q#t��/���v���m�,��v���qn w�=�p�+�G�@F{^�nD;���A�O�b���������4�;�,v���[9��Vt�O���/k��K��m�����wUX���aH|=��50 ��.�ba�1ȳ��n��n/O�4V�Y&��oٽ������2]!A����e�il �|��r������6���peyJZ,Z�~�PR�}U�&�Ͱ0����{��r���ժ��a��v�N��n��U@s�������Y8�����P�<�bI6X��ǲX|����7��d����TQe0�·w����TT���D:�s�v�ES�kQ��*1!��m���P�����~E��vՊ��SO�Y�@ww7�A0����@�l@I!o���r�8��񇢯���o���S;n�m�>�A�2�x:����}o�#|�����酅!�0�~�[����4�����Q��r��P�ڸ{�eY&v��Ap���ءX�
���<yf�6�Xs�~N�Syܛ���������U�S�H�>���LK�L�hZ�A>O�?��,�įL4}�t�"��L�/�`#Z��}qY���6z.r<�Xk�ܨAղ!�vr����l~T
��sϾ�n�s����K�A����ό;Υ��ؓS��6G3�m1������F�s����?�l��z�|G�T�����E���"�u�	n��'v�T�͛G���Fa2z4)�y5n��-�i:O�Z)��Y����z�G�$E�
�S�����g@���M(t��5_���Vm_�������� SL��*���j[P�4s&WX��_ߴ妿ޱ���~�Bi8� �Ϡ �H��F\C������ϟ��#/U*����=�D�>��%�M���	;�lὢ�G�l/�$xi<��d��<v��� r�w]��g���W�cb��6מ�=����D⇙L�7�ф�
B��8?�W��LQ��Eǉk�04l
�ӕ�S,K�Z��X�������G~g��Aq#Ҝk�8����#/�*�/��&�6��\�&7�W	����ݼ��Ȁ�sw	l�5��c]�Θő)�q/�W����e�����'��S%��@^mo�Ǣ��Z�-~�Bp�T�J�d,��S�d�n޽�[�;�M��W� � nd�4�����7s�ܩ|>�^�	�M�(�0���*�&	�5Ms�M���:�݂p}�$�5��>IígB�q�m��0&�� SdǱ�\0�a,�<|���|�D�7�w,	��(f�L\�c�P�����{^ؿ���]7��A���������J���b���Z��9˲�E	�\;Lۡk�{j���9��x�%����9���w���~���"�/$�����S'���m�u��é�����={n��G� ��0xk zc;q���p8��j�a]�a�m���,����\(�OSs�w_3
����H��?����y)���͛�n�f�O�hj�+�@A�B�`����������r��L��P�A�U�F��@�F���#K��rMP!���L��L4�F��o���h�r��S-�� �XM۽111q9�;R�׿j�=�g�fj�j�N���89kv������e�~����^����9$�� �hf_�0������r��j������d�'.���E��E��wW͹[K�i�^�ϴe�p o>�h"� b�fg����ߎF��r��=�Z��iބ�	��y���F�V�����M����������X��h"� �1<<�9�sNU��R�t���~?N��pJ[����6�׫m�"�(�gR����?��	�H4A��"Du&�N_�p�,�O����L<= ��s�:m�	I�$8��`�7���	'?������&� � �U<���x��Sf���-+���MNQ	)wo޽�I�.]�&� � >���8G�(��}s��)fO�� � ����Dz�[�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA� �&� � � �DA�$�� � Z�DAAD�h"� �hMAA-@�� � �H4AA����e!�3ۭ�    IEND�B`�PK
     eO�ZIRP4#  4#  /   images/2dd92824-eee5-446a-82e5-cb3be823b6e8.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  "�IDATx��|�\u��sڜ3}gf{�%��)	����Ԡ~p�ދ, �
��(!�BIB ��Mv�7�����v���=�w�z�+��_���7�)g������<�sfy�I� �dq�I� �dq�I� �dq�I� �dq�I� �dq�I� �dq�I�
˲�ҽB7�'�)4�z��8h���h`�^_^ �r�,�0�W� �a"��Q*�T�P�A ��`��`�j!������dt�'�	����˂�➃�<���iy|���ލ�gWc�`M-�J�� v�(�Y��@2o��!�	H(�V��PNT�� S.L��g|/�2N����</
�������Z��"<�`�	X���Ï=�=�gq���zOn��}�s9\~�%8i��3�Q$������
����q�T�)0�b*�%.Κ�}Xn1����7U���j"i)(@�\P��:4�@�L��*̠�T�E>�A6�ʦ�����[������o�E��p��	�5O��n�x�8uA&su@�LADi����4��>!���t�
*:�Z�O��yp��	$�
!��A�9$�#��b:�Д�F���w8�����dduJ:���X��-��=c�(������פ�n<�د���+.�d���E�1D�Ĳ�o���Z��
/�k��L�?��	�БS�&@WUDr*�s|DޭA/��2vGdԻ,ԺM�T��TT;,x�M�t��@�$ ����Օ������ˆ���`u�s� &su@\<��#c���/�S5��:2&G��@��"�f0��Q�`A\��HZ��kr���>����a�N�e蚰{"Ϲ*���%9:R�l�ˁ�X
�Ơ�D�̅�`�R}�]�Lo(G&/��r��9<���͙��_،�I�&>�w�ʣ�^G���L��v�霪���'&@Z1Q��L�����#N���)�M��`Zh�t�ԧch`��78�HIa��_wka�+ۥ�"�v�3C�HƛM�%3BR[�g	�� m�stKo��'�f4TW_��O����m�w=�����9���1�����H��R3�~��x��X�qx��b2,4"gZ#j_��!�SM�C`t*"鈋Ayu9
,�[x�<	�!FtB��s|�o��3�}z��@�N_����q'2��<�$�'%�XO�n^9ݷodtV2�]�f��-K����|Ak�5����è-�+����y/�We�?�?�3x,�:�}w����r}��f�\~[*��yp4�t��Dږ� 3�S��0�xe,��I�\r�pTE�Ü��Z	�w� g�H��i��Di!	�u����c�Xy�Ixe�zl��5C��Y�ֳ���m$�J.�]�;����%����;��{�e.��oܣz/H����F�A��[�ˈX�y+.��M�hy+.n��_�����m.����J��$G�'�;SV5�����,��2���@d��JK�0q��'U7�G�� K��{یR߇�|��U���t��с�_[���Q���De���%��3C#i���Y#����݌}�Xg��0�����_�5�W!P�dEOm�rݙ��74rʓU���W�B����x}�H���j��zu@�ne���[x��=?�ҖnI��j���"A����NF��'u��qh0��.It#L�]����.z���mI��S[:ֻ����toL��s�W4�'�s
�|������=�˃Ґ����=���7iKiX���7]��J�#�UeQ�4��:9��$<�/��ό��kI�u%���O�c�w<�Q+�؃�ּ�^r�{Z������9:�BBþ���馬Z�4����ȧN����\򎡉�	R@	��P���� F�)$��n���b �Dy��2�:���u�m�|��`�7���}��\��X���GM�)��SrL(���z�s���'�<��K��-��q� J�8�L�G��"%Գ�NddQu�/˰�K�5㒅�}M��3��{�:��u�>�������6��H�{+����������|�1�ۑ�Dc��qxKܨ(u! @��� �Y#	U/$�mpT�dt�\֓V�Er�����ܗ�-(�|k!�̧FmQ��{˛�~�m��Hj��X�����q�Ny�3ܭCޟ�A5L�/(�R��\c�Y��3�xh�����3t�0��F"�ҽ����8����V���O>K<��=��"��r�Y6���Þ��p4{k8�s�g��A"#y� rJ��t�$��Q�Yh�W�3��t���Z�EU�Q˄FvJ}�ƹ�PN.����2�����h(�:��8�͇�N>V���S�=�x���w��$J�v���N�<l�+��Հ.�C{!���$����9��>&�����(VM��Tjca1>2��s���_ǒw%��K�)�/�U1�~Z<� �:�����
7/�[�PB��n%�^#]1�L�
ޓ,0��?�3�ݤ^�s}kK���Ԟ�]��=��� J���h}�K��<�O�Y�q��^=�9\��U�������ɈFc�F�Ƕ�K��xY7������p@��Cդ4���.9ov��=�k��Y1�ǱD�ߒ��9�\����@�#���](���0K���˓�7p �G��%��!_�P�w�$���`�?�\%�ӳ�.�l���w���Xg���Ι��~p��5��B�읊�^�.����0�%�H��4�ϣ�g�B��m$4�s�����\9�EI�BW(++{�k1) �C��#�w|"_t�}x&���5��[u��?��j��浳Cw��"�#���A�� ��QU*$�d�wQˢ��<�亳$��Đ���z]5%�>��D�������������ފW�V�+�W�x��|&���r1�E�� ��VL�ƇgWsuᚐ��f:[�����76`�֭X�|��Z�I����U�� �*��짖�h[L[�j}����4t��*�%"�UB V��H��WX�i�&X,���#��Y��´�{ƒ��F._����gK��̂�,�ד�HO;X+�4:�%�y����r$'��Ff���T%��k��:k�bQp�'9ş�Tw.��9�9)1I�$�y$��*�E�1�уh2��tF����P��"��kO�f`4���(-�)�E�����22��,8�XT��4RY�%	�"�,�q	c���^3Q���^0��*O;6O���:`/�Eզ�~O�l�Vu��!���i��)�S<�_�I��w;�IH�L�f;wF!�v�&�Z"�©�G{ǒ7�Gs'f2���𸩅8���6Gn�-�o��9��hdA��uj7�en��E8�A()C�%E���G ϒ�� #�3�4���:���CEUr.z�����I>��W�AkѢ��4��DkH��;B��PrXN$�S^���ػ}��w��p@��\� �WB<�# X"g��JCW��]���Ss2�kr�����,�k4�\Nݕ˦���?}�Y��n�j%���w�f�j&�e��S�J����D�ֱ7�F)�;�`�[B2�����*��N� oW�YT�p��R���uH�D �N��%gR��`U;1�&���I�-T�����f�`7*ʚ�y�fTVV�������QDU�,�� `Y�O_J�$E2�*��`$I���(f�#�W9%��H$uA.���ȥ�$�<���렬4�D*�)�K���5�<�շ駝v5�!��Q��vɺ�����?��V0�+˼���
t����]��[�ǜ� ���ޅs���'�!9J$NN>-���J�*�[N�0 0�>78j�&U���0XXn���5���j��lЪ�{<�t9�����!�7��ׯ��o����f����������W5j�)��~��NR�d�h��@
e]�`���O��i^�F��sT]��i:���.����"B�ȅ|,_�N��?���[��qх�@"��W��ϛ���42��tg����F3�چr�����.[1�i��u{����?��vo� �V�x�ڈ�q�(Lx�����D����BK$�H*S��wr0L�EK��/]r	&�"�o_F��"%����y�I�4x���HtJߝ�</�Q��nہ��~���D���HV�yB��HN��������T�;�ύ��'?9�}�E�d�F��	�,�E�}� e�y{]U�\F���5�D꧳-8����oa�'.Y�p��Q[�����UL�>	��L�;�!������[���R+���������24�^��_��ZYxE���^|�Gm�%�ەBbB#�ch�e!7*�"�>��;�����()G]M�������v�$���/	=�iJN7L�����Ub��E�����m)������4͸زG&#�N�Vf�X���U�������Sr{�8�s(T���U4�h��@l�p��ң���/�M�V
2:ۉI�CA,���?����[�/�PI�G����o�꼏�Cwgө��*Zv��3b03��w�"�K3����)AXJ6����Ir���Ŗe��0z�2�}����<dy�x�xH�UcU���w=�$Iߩ�i|���S-�*6mڈ��{�?@lt��V�|��b�o�Q((G��e��������a����EI@6���
p88�d�9���D"���o=��U��> �ptˇښ fNm�{�?����h4��M�9<�'�8������vO�I=P���8: ���gK/�*�I�/��o,�{/A�14�2�co��@	�7B
�w����8q���c��hA,����>RQ�<Us{�ս�Ӣ����~�z�͟��{���[~Z�
�����I��k�3�4�i~��K--�d:��E��bb"�M�2�'��^uũo��~.Z�����!�y*��;/��b�~<��pAC�ґ3؊Ό�i$�,������a��J�%y��#���@!`�J�w���y���+]�m���u{Ƥ��1uZ+�|b�������1���(�uÚ�I��7^�,�ݹ|��m� V_d�����d%�1�*^6j�a�7�ۊ��ppzQzv����O(r�e���*!��ɗ��*hn��E矌�;$N���������9S"�`s��Ry%UJ7��D��A�k�h#�K���F	������8����c/b�q���1�9�g�=�h�\�����o�PW%���0}�]i�8-�KN�k�����C�܏�o�M_���h&[ .H�*qS��ϛ��*e�]Q5P���:R�e�1��I�U݉����*k����8Z�fW���b���Q}U��6ރ�� &��9	��\��)rwv�b�4�ve��a�������L�}�1�ކ���N�I@c]-j�1>6�*2�S�1:E��.���v������������W�<��C���|��|����I�߁�U���'����UEV!/��y���v���b�(ҩ�&�~�kxh�{�<'"��.]���58���� (aٯ��ҷz0/�����F!O-+����X>����c��){Nvu/R��Q]I��!_۹s�)�R���Ŵ�&H���*S4�\.���.�Ҍh,��D��mhn��[�or9��=buu����g���k�i�Ʋ��e�ʝq���q����"�H�Vg��*�`�"�T*I�)^�KyE��<D��~�ǘ�o첮��"|�}8�u�¸����z����~������&P�$=��1����3�	�aX��n���~�>�o���T��Okȓ��A�0�]A ��赲�����j^�L%�H&~[T�R��0�a�4�����߳y�]b
d�7���?��g�y��}���3O?�P�&��%ߑm�chB� "�&o�WZ�T&�8e����M�\,�5���n���mw;N:�C� b��47�iOL��J������^ WD�,���%��AJ%Ppo�Ҋ)��0�g
�D֚��z���#��y�f�I��J�M$�\_�Sz<�L�Vpp�����/P�5��\�GC�	�r����8����ûvw����ܐ���:�?�֜w.��&����ƢV��m�T��otIն��#Q�@Y3��^��
-�ݭ\��]��vC#ueQ%��зk7y���];�
<���7\�]�*� bg/	�g�<�]��'��L Q�g)��Iu��y"e�������mU��nLP����K8�U�<)32��)��!�&jAUU�Q�Y�ڟ������x���jj���{nJ�sW�bji�ڹs�.\�eK�% k�n���h�����}&b8c�|4�z2u����������,ǯ~��/}ܲ��%TUC�1c�sA�遻4�����8:^y]�Uy��w� ��gg֣��	T��x|������_��>��fh5J$�^Dɘ&bh!�[tA���N�*����8���ωN�����tw	B^����'x�{�`�^�p���Mo���j�,^���v�������>E)���ս#ڠ�."��G@��Y����m���ڴ����zOҹ~�w����_�r�cfE-�qsP�d!JB!,]~2�5�gb�.	�������Det=�xg<��E�9|?�	���j���v�e��[��7E�j�REˑ�fPᤊ�j���b�;ؿQ1��Ѐ`�6�;-R[��ji~VC�ZϞ�=�b�E��s��mI���h>_��z�q���~y�f��w_Q&��EX���	⦉!j�y�w��~�@���xq���J��B�dOZ��/~t�x�3�Q�9���ͯ"��Be�/]�����vuCaET� ��#��o�
ɧ�C��7��ڢ��'������G�~�.(��Vq�w���/�@�#��ЮT���������Lߝ��A>#��ؙ�0���%���6���#{�=bnuRV>7�2~������M	𺩂(����y�Uj�f�6�h=���߽��v�����Y�҇�����AJ̇��Z466��1�;wnǴ9�G
j�WK.\����>�١���D�$*��xW͝s�<ںsZ��ލ��W@W�v�Gcp���Y}ɴijX;"��=�'n��<3\q�Gp�'?�G׭��<�1g�N�\k\"��;G~2~v-p.?�'z��f�B�H#�tu�\���ܒ	��r&G�ɢ���L���y�xF����sC�qLki\��\����*9�o=��;6\��LD"1Fޖ�n�fa^x�g���C'�l��(�"a��x	�{}��r�͠i�4P9�M��8#PO���Ķ'֠�Z^���=?|kq_�Vy�l����*���e����'�<�T���4�񒥕��5��yf�:Q̔Q� ��v!CSD���Y|L���2��A���R�����ϙ�(���p��Y2Ɗ�OC�<��ر����1���憆�/��W�*�y�I��ς����<�<�3oj:���}�nhy��w!*����AW|O���THe�/�=8��7q��Ӑ�/�ߺ	��^����_[�q]�R���xx�9̝?��u��s�G�}��7����]��[��xZˎ���뎜�8e�Z�h6�ڠSJ��К�duk�Tn�Ù�5C����-0BQ�S���x���$�r�R����
GH�3HS��U��*�����v �0������dXz�b�9Іꪘ�:��������ի��k�6��݇��t���R޹Z�|�;֏�Sp�j�ǐ�1�8�o�,���?��ޏ�,=N���S�{�!�z�%~p�4L���x�s��[����;f�|��ύ��/�,��2ev���K*�Z`7u�=�`�m�D�~�`?��
�:X~�'��Lu���}T-�{$�R���UE���h4�D:_���B�c_2d�u��� �r���{�"�y������؏�T%���vm}j͓dJ�/0����s����N�l�|�8��VVP_V�)��%9ǽ�,-]s}_������@ޣn�\����b�ƍ��t��u| W�u �	<���W�?��/�	�;4���"#X���	F⦏.ǯ�o<`0�M���88&UP���g��_yy��X�s��#��բ�]\YV*�%H�d��I2�|��E_VJ8�[KC������[�N��P?,�Ħ76�-��}����k�{${�]w!��@v���]���x;�d���}����gל�ƀv�x����sq�>�O�n�[Q4��������Zi$5��;�ژ��Q�毞����m.�p8R�Q��̢�2C������Q�!c)J��M׮r0����p���.�P�0
j*Hk��n.��~�O�ɇ���*�޺�FD�Fq���c��wvka��b�����D���!~�ٗ�C��^52/�}HY�c�|��W�#'\��Eո�����H�wbv����t�BN��,w9�A\eq����'p�}}��_����2L�R���P����?&�%�}��*�M	�}���w�!�q4�e�UŌ�cޢ��Pd�߇�U�(����}���	�?���'u��cY�0;i���cI=���(�T9"�[��t���ݻ� ޾��v4�b�(��L�f�e=�:gR�3g�{�?��ZMmY%R瞏<I�����ǣ&T��S�ɻ���X�w��ٳ���iooG&���t���6���Q�����mW�q���eQ����^�_��|�1o޼���}��E᠊!��T<���F̟��O��ï\�W�Y�f���d��1@&Yd��1@&Yd��1@&Yd��1@&Yd��1@&Y�?�͕�UP��    IEND�B`�PK
     eO�Z�IQ�H� H� /   images/a05d3615-68b8-4f26-98d6-1aedf7f6d878.png�PNG

   IHDR    �   �T9   	pHYs  �  ��+  ��IDATx��y�\wu��\s�y�,k�lK�-� c��? �uB @��n�{�^�������t��u:Ƀ� cc�8�x��³$��,]MW���C���޿SuU�Z26���ǫ\�N�sꜪ�����ۃ
�0�0�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a�a�9�8`�af,�a����a�a���a.A|ߗ�)���B�P���J���0�{ ����@a��Ŗ�����r��������`?�5�0�,����N�W�������iZ��z����ҳ�|��D"��a��s	1�߿|tr�s���Q�T�d2���{�?p���ѡ�J6�}���)�0�,���o���r�Z�POO�jU�T�uatx����mKW,sS��\o�$IE`��5aq�0��m��gδ�Z�J-������N�R<����v��=22RD����0�,�azz�xc���P���ƛޖ+����4X�}p��q��7����nKO���p8��$
�a�%,������~���N���yrl�s��+���"555������ٳ��}�ۮ޾�����SI�>n6�0�s�@^ ���LM�<����=p���믽N�,��L&#B4��Y�f�'�����G�����0�.`q�0���_���O?�[(����r�
8v��>�&�-mm�-d2((v����a���a.!��{h쇮�z��v�ڵdrr���ѣ�U�VI����b�

P�_y���>~�6Ӳ?====�ۜ�
�üSX0�%�����=;�$
��7�|����pgg�433�d����=�vǮ���3�C�P��f�a���a.E�!��o~j���[l�L�ڵk���_���aX�x	��g`rdL>����˷n�T>�'��K(,r�0�+`q�0� 4E��n��������
�R��C�گ��r9뺰a�z8z��42<M65�_�jտ<5X�H� �0����a.Qj��W]]��K��r�����Ύ�XGG�l,Z�����'N��6��^O�3���Y���?`��`q�0�0h�4��g&�r�С��ǎ��áX,&���B�P�&&&BG��v�u*�JcR��3q��a.����)^{�5;�3�ec�m���j�V��֬^�bQ	���Z�?t˝C�g�QP̼��\W�,	`�}���ĩ��^qŕO�\*���������-�_~���a��+��*��g�Z�f횛GFF�6�^��>E��|�i�=�t��f�)Y��p
��aq�0 *r�F�����O�8�r���m���ɞ�)���͛���#����MM���ݝ�'''���tc�|2sfo�[,˺�Z��EQRUuPӴ��z'�9�t0�`aq�0�&����t:��jV���߿���I�D"���
}=����8}��X8�A��"%0�ܜ<͹\n�U�nnFQpY"��9�#�c��y��m+��n3�E�f���a���r���'�� ���7���~�5׀�H�b�2p\K)r����ݴ�MS��ər�l!C��߈F���lB��ڎ���@UU߻�4�2�=����q\3�a(,fQKo��k��;/�Z�u�\{�T5�m��v�
��B7���+.8a�nދ�.|�,+���wM"!���
��L�R����p��Y��8`�l�#?:|�p�i[+���W�\)�E���Q��t{>_���*��Ln7U�@@�!K2�!�hZ�_�l�fڲ�	|}�Yp�8`��Lqr�J��M�f�099����CC�.i�&]u�U�
%#�0(�*)�"D =� -�s/|��8��,�
����)`fA��a(���ɱ3g~���O�I�ǩӧ;.[�B�m[���b��h�%E�a�1��s}N�쁿���O��{��9��,0�``q�0��KO_�e�c����Z]�������)�|ŀ'��y@x�ބ�A�=M��Վ��Y(�p�����a,fa�ߴi��KO$���uv@"��R��,) 
���Nh
b�tN,4�Nz���u�ӦiNR $�l`����Y�DK�ܒ�7o�VJF"�$��A�l��jb��Q�����I���=�&�$t�ԋ��#�ju�q�Gq�)��0�>,f���:�N��ˊ�E��ׅc�fߗd2�� �\|���g ��S>	|V�Z�B�!��Z�"a������f�K���FI�J����߬����Mh詎�䐁o�6|�&	�c�#��}�����\�P������\ڰ8`�f�X,�D��m;�Qej�1��n��3p�}�Iel���:5��܄���;����e'X 0̥��Y �AVL�\�#�O���Y|�j��뢠3@4�=_4����q]�������Q۶Ǫ��p�wpd�K�p�8�s5�[Ѽ/�Q������9���y��ϧ�����ɟ]�:�ׇ�N�P�1\/��s���a+�8/S$Y�gУq*�h�v��B�`��hX�e;h��Z)����S�D�|��\R�8`��YlŀR�������!���	i|o��|�P4� �J����(�+��4.����҂��,J(��>7�Q����+A4U��9q���_�B��O*~�{n�뺷ض�U�����0sI��a�H$�f�Xڅ��OQ��>��yq��xPh ��|�0_0ԧ*(������J�eY���3(B����r��\�8`�^�Jk����x+ǹ�v�����Ms��������&4�CC�@��A6
=�oe�a����(�r�5E�uY�J�&I�hOo��L��M'�/ˡq�����RE�!����m�\.�p�0sQ��aTW �ϸ���y�qqOc���8�B����Wy.�H����]߻��g�u�ه�W�a�����	���#�[��[�{�'�u[�=�ι���[5��^�z��Z���y'��
��MӜ���ZE��(aq�0*]���UV�k�NG���&Y���n�68����d(�w�����qD����j��(L]���b��0',f�R� ��d�Xf��y�qq$x��ޮ:ⅶkܶ1てj����{}T �X,ڱX�Ǹ�Is���a6e-��]{��x]�z4�[�$JA����.�/.T5�͈J��k(��`�;���MMM��7ib�������Q~��/�phE�ݥ+��i
�@A�2躮��+�4�<����yu�K���`�x|ڃ�������r�/����g��0,f�S�?�,�Ǖ�WU�8�o�m,�BA���(�}�`hl����4�]�y�������xy�1����ɑa~��8`��hpM4�of��ߗ,���ֿG��0��l+���c �>ض='v  ����ynm��ϛ�|��|��a�r��Eɕ7>��ݕr���Ͽ4���Y��q����	U�*0���>������L����Rp�(dr�׻5��Am�s�������iv�$R)UEQ�Ȓ���������t:W��F^3B�nLƓͧ��O��L{GW������ӕij�͵��J /����yoaq�0��8�����3�R�r����#�rE�Ѿ��a�1�V�5��*��1�uj��`VC#�י�ڲ,P4U��׮]�����{��}wr,�y 9z(l{�p��(�jF��ɐ�G���Htd����=�7�<9�޾����apX,0�o��Y����cp0k�#��?���N�ON��km�X���?�E�Qa���
TiYUE���&J����k�<[
N4#����ʦg`떭��'���Q<&ϰM,��_U4ח4K��vX�z8�?v��T,���G���@wg�Xϲ��^:8�bE����ms�$ü{X0���N��g�LF}������gϞ�K��z�f�öݶb)�������[o��L
>$�@�MSg�dy������.Կ�B�R1!
��I�X�=�̧�3�w�^(JT>	PH�l�>(��)P�"�}q��\�j�u]�:3tf�8:�H�ɦ����S?��g���+�[���m����a.q������`����-���wMLL,��J/.��K���j�Ҧ)jҶ���h`}%��}�1i�������xL�"�N�#O1�Q?����<�;�q�zV���P(��*B�x��p���3����8z�$(�g�Y���B̊Fb��U�Y�ͪ�W������bq��"��F�N�'�"bG^K&�wv���w~4һqe��k�)�P`���a.A� ��n:p�`����ok�F�7��ٕ�Je)�4�8��c;�e<�" בh��� �-�< _��W@�Chl}�90���۶)�Iz���|S��0?�1v��2�TCx(Ц�+�-|��
��c����F��2Z��>�Q�+���PJ|�mEQu躱f:����������p�T��7����{�����yۦ��M�*��0saq�0	����<ff���R�Rq"�J!659��=�tb||�����.,im�h���	�1W�#zڶ^�@���1M�22�U��R	�=
۷oU�E�D�N��yεan|��i�0���8��%���72���>�� ������
D�(T�.�V	TY��b�pI���a�D %��V<�'u���^�Y�W���Ux���O��b���v�����+�w�cgW�X3y�5+˸>m��N�a(,�wL-PP<N�)�T+��v��X�Xnʤ3�\6+�*�b�/�Jm�|��j�=8:�r�-W���M�eEhXMF��zH�sf�1P�"�����T3�a����ˠ*:\��*0�*�b(��{p.��x���������x>�J��1��d�e0t<�H4
�]w�9s}�Qp�*'�~����Y�$�*:�O�k��b�(>,!�$Y�D
�,�QUU��Uh/ds˓���:2����斖�Ͽ�����W�=p`bfӦN����+,�HMh���J>�)�܌��/^NNOdZ�Lrb|��b�ڊ�\K�XjuL����}�˄�Q�uBh�YQ4)�U�T|�|Գ��QxN2��xVE�40MsN�CZ�(�� mB��?ǻm��(.p�n�q�툔ƹ1�ԹPm����gI���b�"� ��ڶX����;�ؿ?4%bP�V _.B<���5�/�dA���9!O�Lr�t��@"��-P6�G!611�k��`e>_�ahp���w^�d�%˖}��7�-j.,[��
�>��ü�P�����1:ZR���н?y�9�IwOO�:��T[�Xn�V�N�r��i���q��vÎ禍�+�窾�ҳ��XW�?�t>Yמ5Y׫�
S(�j�p�v�aժ"����+>0�4�wl������~z�����]��7�S>�e��	��8��q���>E�Z��	ρ$����j�H���?��?���I�h<��mUA�h�^|���`n�%(��~�c���,K�7%
I�Y���b���	w�������N�<z�С}�]��~��cG�_�%������	���@���q����F����?읙ʬH�g�Ke44�.˲�M�jv]7����8a��T�wd]�4\�纒C��vJ��PEc&Ӵ@�u�!a��< �0����Ā��{~�?E�hov��D�ׁ2r�|����/�#�(�b?7���7���
����H�F��P�`9�8� ������+����������T*�$�(jtm�{iv�z�sf>�x)\q>T"�P�
ϊ(��Ir�\
����IF�����m�|qpld��=/�z�����OO�^�Vb��,dX0̻�����MO�F�����\��*�έ*��+�k�eU[Ӣ��
���9.�G��8��GE��/�A�U��L����퀋�Y%��	����;��P��%90�$l���>� j�D�PB�q]Q��R)����r���0�{��կ~U��M�U��ޮ���,t~��H�j�!�2���]�m:p�m�é�A�� 33I&�Z1g��ll� Iv���et�D �{W$�P6F,�/5�r�!k�)I(�4�zPmɑ���^^���㓩}/��煍���{饃c;vl� �,@X0��PL�ӑ����ӧ�7���X<16�%�/l�Z�R�v�Mӌ����<ϑ|r��άAT�"˵�THH�Q�d5�'(�-o�*!5M	Z)S5"_RE0!�m���ڲ�B��ߒV(��؎%�hz��I"��VEݡ����@#,�+�g���������g��c�D�2��m��G��;;o b�������2�~E�$����)����*��4�N����c���ۣ	C�< �H���<�WM$���3@ъ�f�s�߇�S(���sS(g�+䄩�I+�]5[3�j�m�k��ʭo�y�����_|���¶mW�رe��͜��,X0�<�=���/�>����S���^115�ɬV.3��b�b5SQ!�qu�����y���P!�"�00�´��� 9��f�$QP�k)�@)X�X|�rA#AQ�����P۷/l8}��@1V�
h��p*"��rac���M��ǟ|֮_W\q�a;��W��|t]���˵�<d�g:�;���	^�q�@�B��h���1��p�Cc�Rׄp<�������o01>��hӪ�?m��!�C�0�*� :N��ǎ�A7T
[������Q$�o��IU!�h�����[VJ�Q<If�q�Ո���K������MG�ϼ�kס=�]w͑aߟ��E�EsI��ajPa��L&���cǏYy�����c���ʆR�؋>��@㡋�;*%�F���|`(�3��ED�����hZ�|��ʂ����9(M,ׂ�$�Z��E��#v?�{�����?�.$J-eq�O��]����j (� ���-�SY���?���X�d��D��A���u�z�m�ߎ�O��<B��h��д�iZB8��9�������s����N�ڣx)�NQEVB�hq Y�cR�#yKW�o48*�OFa����#�lQF����x"�����.������a�Z���ry�L*us���W6�]��͛��I`�K���z@�ٳ��?��G��422���-�1-��X,�H��5U���a���k�
�b�.QF@��G�pd�g�.@)���z:a��! "����G�	NCϠZ��'R�%:����uP�lց4�3]׶�2��O64;���=����k_�Y}6f��5�0��eatϥ:J��s����A��L>�룔CD�\?I� ����J���F�t�7���Y
�
���Z��:��!(�����Bpn{��,-!M��=��OB�Ѷ�k��M�q��Wh��1H�tPtX��B�p�%a��Hy�����w���g��9�窫֥k��撂��o���`6���ϵl�*�No)W*K�i��+?5��@B�fٳ)��T�;0;�f���y�l����{�za�Yٟ5�AL�$�	#������0�s��8?�k�( �yhA�HJ�͞��!bD�(��W^ރ�}�b�vA˅�u���_������
�8n�!���g�@�����ct�@p}��O@�����C���%!À�U�2kͣ�`��V��i�8�����bʄD�n���!/�{ �`UM���9�E瘌G�T)KN�l�pn�<99�慗^�x���������cGV������os�0!,��d�O��h���^r���fRS�s���R�ԍ7��iV)�PRq�Ǹ���l?
���8��r�fH6�n|���Xw�i������O�����?w��)���v��3�l&���~|�K�4%�p�"KA�������2X-��:�kqO?�8\�b�y�P(�D�^�TA#���P���e��9N��\�>�
�7C���{T�� �}����/�Lz^|�e�¢_D�PD!��Y��7J�9[1��C(l�QP�e�h����A�b�@A�a%,�8�A^��G�� Rׂ\���CXā8�)�U7i��_S�VV�3�kO��y���<��y��̥�f�CS##`�����5�����\5���ʢ�UIKyݱl�^+@����Oƀ *���`����s�z/��X���˱���{Pw��s�{�'�a�����Q��W{-��{��0u &+j�|�e��p�$P��є<1M����b=C�g�@��o��r�y333�T���������|Ci;��@�Q�A)��Na�9�Ba����կ����#G�Vȗ!��x~�H��oצrPp�A��-'����s���s�A��Q�p��.*���N#��PE1�P�ExT��S�/��Y.�Z�7���=��={>���ھ}� ���A����f���I�ƞy��%{��_sj���B��r�\\.W���h�]��H����>$�f��A}��ڵ�B�TC]۴��9��~-Q���S�c	eC�`��	����6�C��h�f=� a�w_��O����'�1RĜ�^��"�h(tF�Z�őoEb����r z� {����_��?��ŋkM��N\H�c�k5/ʹs��AD�����EJh�R�d�@�2��[��������߆b����A��F��"�rD삅�����9A�bѼ��i@�<�p�=�� ��bP$���Ȯ��z�Y(��R��� ���D"1��PO�>ٞln��jUW}�_��a��-��r����;������aq�,8(��ԩt��gw_��k/_svdt�������k�V�0��j4��-�T�Y����Q��f�����WRɠ�ѣ�@Z^�m4;Z'�������@BW4H
�	/�7���TaL1� ����T�ǥ�*%��a��$ȭ=�W�e<L��?q����Y����C*�R�Tq�h5|V4J�-Q�@��Lqd.�8q~�!��~^mk됳�4O�m�
ޮ0ҬGe��������I���*9�s�\[(�@T$��\.7\w}�n����=X�h�:m�YAQ(�#j8t�����w�D�	�޶������"���V��jMϚ��H؃R�(Ĕ�W�T*����6K���n�U-�p��l��ɗ_|u����3�����TC�"���`����g�?~��e��vxx��\6we�\�T+aJ��xj���ԩξO���1d�E�M ��^�hnoY��:��t7Yֽ �'զ�Z�Y_*��6�F�D��N �H����Z��r��pc/�)�d��*�IV�h�
��U|��--<N�r���2���G��LU�|Yu\S��C�\���Q�'\/��ƣ�$�82�*���T��g.55����?��><_=v��=��H�,2ꁏ�쌹M��ޔ��r��1�Y�q[��<t='Rig�����ю��>|+�>5{�|C|_MI�a*(�(2�f��������N"p?���@b�T.@��鐔�IS���`jN�&T�}8d��J(^��uܠO��k�6���ߞ���V���u�cz}#�Μx�����׮]2�����fA01�G�ӟ/~��Wn��*W7U��b�Q�mQ5��W�H��Ws�����_��Ǒ�"��~E	��y��A����\z�Z ����BR- P�\?�J#�x(V� �"Db�Zp��ÆL�>���h�0��e\���D��U�d�Pȷ턌�/��*�Ȭ�)�~,󋉢���rY�UcR%Z�����FU�]W�ѵᙾ�z����ѷxqxj&�t5����ζ��7~j�U���������$l�Q�\����^���3��0�=��x^E���8�O�]w��)���x��7�ﲈb��2�T�ihjjq9\�4	�@l�ۢ_��X��]'͜,�W$i��(�^%]x(2^�������lU�%
�pmoQ��7�}�������~���pW�T��`q�\�P��������������O~�Z)o-��}�B����BU�Dq��\~О��A���sN�� �M�Q�?(X�#�-4k�`BGt�skA��۟�����i���ȣi�-N�R!赨`XE{4���jŪ��$�L��=~!�;��躨}��Q�?��_��ըST�ď��_}]X�#G�H�j��f��J�ӌ�J�T��G>���������x^j��-�)�AT;Դ��&�|i�S �@�Dź�o��P��(� ��
@����1JX�PP�ҥ��;?�>�LMM�o��Q<x�g�Q���<��B1��R�Ez$y'DG
�tqb��8Ӵ�g�~G�D��/x�/�¸O_�Q?a
Y�M󅸠�J�xB���JUA�8[._��=?{�E�O<<44�Ғ%K�_�{��s�Q+o�����������������ƶ�K�n�4C�dD�!a�D|�hhd�g��A��J�6d����p��mhI ����IRP�>I�����%�I<��	C"b�*�khZ.��'�onjy��s���ֱ?��g��W��}��"��4���zH|]@� 9�̩=�wUn����E���������X^  �|��է�m^v��j"k�^�Z�;D���xG��{&�	~�BZ[��hJ�,��*XK0��.���B�jA�Ԧ��v��`^Q^ڲu!"Qb�D�a��@>_�!�e[����-��DX��K���(b�����R.��NO?�s��O�x��<�20��	�%y
>���+�nس�����m�Ym[V�q,���Z��h�a��=�0<*l�(��0ƞ�\a0[���jufk4�B&h$K�Ĕ �M��
�!"�3���w2�3�I�g��pKy1��Gc�Z�	�a��4����D�iWgk뫋W,?��������4'�������o`����t�����e�����e%VdH�.���-�#�|	�S��R-�VtH�RC���r0�	�B�Y�	7�FHgf`���� �~E�!��bV-�E��k�l��j����E�E�q�H��=�oL�^_��BH0">!B�!SӦ	�����b(�`h(�~�T�����QI4Ғ�R�Q�hR�`G+VeS�,7O�R���y�̙�+K�6�$�E`~�8`.R)?���O�ڽ�����?��f6y�ߒ��2��pT]�J�$"��0QC��< 
��R�57�*�"���wj8�r�uA@�r/��!1@��6��e'��´�6��'�E �L����P��dss���Jɲt$o�ݷ�gOO���ɮd���o��q��?����������{���h�7��Q�,��J33�,Ղ���Jsl�ыs���S��_+*����.+�(loi��n���'���~H6���B!_���$�6<Rc"���LĨ�!�m�l��b�=�**_JjKA�.�E�U�𷌻� 5Ҥ�K�&���Bq5bb�T(�@��>AҠ�ۀ��B��4_*|Ҵ�%�ӹ��n���x�3�����aq�\���Q�}�o��7o9���L���\.�XV5$��Q���i�������v�FA��&X����؃���"�*��C���u� !ewk�pBAjE�Ӄ����'u(2��+̺�ɕL��.��B,�1�E"�#�D�)ꌮ��Q ��hɢW�-��Hk_k��k�����hy��''�3��"����{TU��z���;�;7���P6��p�R$�|�E6	���)p�h$��?�}�m�����hSgO���*"�0�=-����h8h�q�^�*�\�������~;��,���%y�MOA�P�b�ԕ��(Vb�5��"�!�{CQ�EJf�v�Lu%�\���bW)�U��j�fs��ڻ�urb�k��|���X���‹�9p`"�/����W�������ǭjue�R�;���t͓/�?�����!k ��J`|��)r�Q�ߩ��E�cIt*$sF��*��Ǔ�PlO	'Ƨ�  �@Gt��FA� ߝ�y
JyJa�@��M�c"���B)�0�;�ڟ\�n�e��N�A����VZ����{�qQ ��G�����Q��Huό�/@��T���[������5n�7�� ?9��[���"C���wͺ��?	?���0x��vt�)�1�b
��u�MS
���JE��AmI	���j'mU/�Y���G�ñ)V�g����A��c�C"pQ��e��+D̄���,��z	a�钂?#�Hd�N��-����x��͝��,������]�?��;&&&�ڌƶ(�M�%o�
����\j�d:`��0�AM����O�=�f�TE�u*���e��3�lK��baHă�d2)�����Af�u�E8�o
���4W�ɦf ���oh|b��FK��O$�n�S($��t�<ӽ��卛7�����x㍮t��-�@�v��yptt�h�ۓM�$QuH�Y��<�$�ZNC�9�K�l*�X�X��k��8/��������p�n����V9R�ѹ;n��������B6�CTKb�!��BaP�K�׌6�Ēq�.�H��G�8Ma�*e!--����U˦	���&~�[�"�b���@!�Mf��k����ɢN��RKQp~򹝿hϗ��ʾ�xq2+q�[��sQA.遁L�������w~2�/|o�K*�r�����֩����oǱE����D�]2|ZW��6mP�F�e1@�r!4�Ѧ&HD#xS82<~�x��n���Z����(�8P�b:����I��H�z/P"{H�E�zKs����D&��M�Z��_\�t��.[zjˇ>�_(7��n����K_3-�>�=�Р���VI

I�δ^Itj��|�[cje+�3�S��*�`�uES+j\���L*���18s��~m���o���e4��ۇ�a O���N
	��{:;�W�Q*	�IB�zo��us{+�RWd0T�Am�z�J�n����O(WPp&� 7'�ukj�D���$*����[�"��l6���-�w��E���c�(5q�.��o�Ey^}���Ǟx|������Mss�TmF��j
�bޖ�J0�o��,5N1J��63�Q��uZ�>�@��|5@Gk�XF���itK7���q4�i�z��i*���ֆ�aH(/��ffҢ�yL|M^g�x�K6�MCקp�C]]]/�Z�b禵k�mߞ[�7�;6e�>�|%ި��gP�u�m��F�%(��[�qnan$��i��M34�;������k��?�y:sΞ=+�4� ��UMa���	�0�hTą��"<?�"���G�L,�g�g2����"���,SLC�3M'Qf�ZUA΁���zkio=���ɐ��T���*���W��ײ#3��K��;��any�����m����Cu&''#߿����~m�S�K�dW�4�j�DM~tQ�>�"H��4�o�x#��Q��m
%:R��2�� ��:���0mM�D��(Pd�0p���	Q�+�X�ǣ����d�ZZq��(sLƁK�F|���

���h����k��� ���֬[��UW[�}]���`����Q�M��24�7���om�tn:�Nc���x޺,ض��<��o�o��߫��>������o�Q��h�wR-ѫ�
D�d�P�		9H7��lTJs�,!(���c4�,^?�lJx��Z�h����k��)\i*$��B �,�R)(�K��� ��<�a��Ѝ����|�)[�߇Ǻ���y�aq��^�i�Çϴ?��/�<|讱�����b:�([�M"ؐ��m��_�j)v<�zȊ���" �J�����������XBx�V�,�Trȥf`jfF�S�Q]kK�H3L4š��]��(��摋Ŝ��g�@PZ����h�PL�<\/g����z{^X�l�έ[�8�#�~���������C�m=��<�YK!%�!p�@ú�k�+᭍���A ��A�OC�[7�rIu�HF#q�Ƹ}�v��=��?��?
���f��h���|��2q�^�(1�%�9wIp��Z���X$
�x��:���C0�Ud����S$�@�H���,6��rU?�~ҥ FEdWě�Rl�����V!_��i�ų+x���1-����h����?�Q,~x���Xƙ�{���	�_�b�ҧ�}���#�*�JWP�D�H����61�K鉸\�/�⨝*�ջ'J���R�o��B����� Qmr�8J=pto�HnbbB��R*:
��!F#?��Ǜ����]#���M4tL3S8��S	�H����� Q�e�9����V<z���;/�X����>x/X��;3trh�6��Ԍ?Q����|��0����*+�g���oXQR��Pp
�M�ͧ>�)�?v�~�9���MO��� �P�K4̎Y��U�dSb*���j�B-�mk4�@�alj����J �#195�x��~S���n)`U����9�c�Lq����G��0���Y-�EE�H��I�T���车U�����5H	���ݗ��yaq��^���w����}{^��������2E�B2U����pТ�J�VU�򫢙MtHq
u�U�B�� 4W��6h~D��FnY>2p
�PP� $j�4D\/�A��M��557���/j#PQ�RID��(�<xS�D,m�-~<�ú>�D�.Z���[�z���݃�n�-�O#�)��b��c��u��(��VZNn6l��l�N�A�՞ˁ���Wj�"�7M�U�a_L|�K_����0008[�PZ�ق---҆����L{S���c�G����orrriT�]���}=�DE
e6��kp��A���B1��,�(b�P���1��)Q�Q1���E�`�z��G�iV��~ʐ��@8��q$&�4�RU%��ڕ�f>�п>-�$^e���W�8`~����������w7?v�+�t��|�؆F\��w(���tC�n{�X���V��"����h�d ��T8���MUՃ&9$
h�`bj�SS����J�bF�$Ba!D�MM�l�GK��|jDF#�J�:�\FtdD1 �j���X46���utt<�n�ڟ_���S=[{�>�lٲ���؛���_R*�-�H�� ����_����A��x=D��^S�B��������+��TV����<�z�b�
������Ѳd�kP�Vn���Rg{������B�����%�+��(����L:
�L
r�?�4�?;x'MS��2SL���SC.BTJtA��N�B:�Ϥ�x�7@�Ϥs"��,r�U*E�q�m����_��B�\*~�����d~cX0�3h���7��>���o:t��=�ru{�Zm�TCҍ +�R�(�����q���U�C�)�V�_��� ����zb�6�H���C
B��w
"�M5��TD4�7�HD���n-�{�5��Y&����)���J,b@K"�F�6B��X��u�.n˦��_��ʴĩes #�>���Ǥ��h	4�78��.j�,�g14"F��[c�?_|B=��\�c����J�B�p���'��<p��P��W�-F��׮�[o�.�|tvv�`��HV�2+����E��S#���Ã){jq$֒���D��x=����*W�05=->kzb�[�`E�dsi�ΒA��f൙�r�ik��r!�G!
�~bA*ff&hU�
e���@\x2�K:�*õ��}����}k�7���;���/~�g����Α�;|_Z�#�D$�$/(2S���R*�r��`�m���*�b9U�S<Lr+2$��%D`���(L�S�k@�k�ǥTE�#)*t�����FH$�Ќ�Z���FL�]~vpH|��b$��M�����'�蛫��xt��5/,޸q�F���������D�%O��4���	�1ly�R���w�A8�v���yQ�P
�FS`�=w�G�ݯ�.�_����[Dzbooo���	W�s��:�Wo�;��3����JQ�]�4�D�K����o
��j�S��a��P.W�U[k���A�X�X+�����#�F�MiDs��l�w��j7-I!1E�{N�X*^�ƛ��O�����f͚0̯	���<��S�=���KOOo�+*�J���C�Q$����W�V�T,���4E��l��Z�#Q��v�W�
�)�#�ֆq�f���a�HMC�Z
B�$#�����(���Ơ���DZZ[EZ#��IHЃ��m����ɸ��r�p�Dww��׮~~�Ƶ��o�R���\��@��,?��vX�?Gc��1�������Wm,����=�'�V,��~.���_������Uk׉��E��i�&�K%�U �V8	��/����涎�.Ӫh��A�j$%�Q`$arr
�S3�T�3�NCgg't���ؗH8.�_z���c��Z_��������6Ҷ�r���N���8.�[��~r|d䆗_��W�����y���uaq��V9y�7����޵��/�R�����Eh�d2)n�� u��f9�b��Y+Xt��)�P49��8�
�<����tZ�Q���*��#>2 T'!�Bkst�����o��m8$*�Q.;M%P��4>���CKS���`�9���⥽O^}��=�V��K�]Ɓ_�P�{Nf�3Ϣ�nſ�������lj�AO���=ۊ�����z[�����H �s�=��栫�zz{�Qi����"�S�+��J�H4��g�ݚ������`(���*^��/�]�3�����@�e5��/����
�J-���G��8�\A���k�>�)�[�8�CA�O�I�%�vԞ#���k�Ϻy��o8�iW��n.���:�8`~k���=������_����z^��ky�b�i���(R���ܰc�J��"�%"PYY�r�D�#o�F0�k[�O�ѠO��ii��4G�Ũ1R$�H7W�p�����6Q렊�L�.5�ނ"��ɝ�ױ�����DN��5���˯|��[N��^]������&����p܎C����.6*1(`T� 4l7oGs5���m�C�
��3�0�@ ��iPEF�4&ZZaђ%B�E|@�I��>*�p�O�*�JEZ�ti�=���|��+sz,�LLNNJ	���8������)zp�x�ҹ�Q,dr������.���Y�,]��#�K� ITM[�%U�L4��n��5�MK��<�Yʰ0��Hu���Yv����-��uos	�}ü[X0�9T���ё�'�������1��?����PHr$#y�%q��*JQ�����s�7r����Φ�&�b\��!5(n�Q[[sRx�xs�75�͸Z�;D�"��e17LE�r���Fhom���ݜ���45������M��-7ޘ�)�����O�ZRz�Ԋ��{А�p��g��{n���ȉF�*ivu���M�N��sx]R�B0eЈ_�J�I���Y��n���O������泹�h�c�T�h?�{hʀRjQH��3�xPnPab���������C�P@�x��I��J�I����D"	==}�#QM=*f��K޴���$��Ԗ�?�󹝠��7�|��@`�,����0xꩧo~}ϛd:�v�v�B��7���F��V��L�M�7c���be9(��	$����bDA�VQD}�q�_q��1T�8��\/� 1��mCA�ln�ވC8"�$�͋N}cg��G1A�͉����R�e�$��g/߸���1��~��K��~ń�q���5�ؠ������~�B!0���!����\i�����B5,���۔Q��x�eW�Ċ��յH��G�7��Q�X�u�O�����3ӯ��{H�B�����zH

 �bz���:��@�}���$�q(��(N�X�x�;�6L�8��ʒ	E��Ŵm{�����"�g����Ԥ�4-��{.
˒�1�,�ʕוn{����d��,����{��=����gO>���{�o\ۊ�R"2�կ��J���aP�g�%W���=t����uP0hF�&��HoJK,�3�T�i]�Q���X�JI��koȝ�d�r���t|�ː�Q�t&��#��Ql����M$�S!#�ڢE�Ol�nǋ7~�F�|g󞂣�bz,�G��9��_��~���[2]`6�^��ܶ�� ��ߵg�����[�(6 �pT��긌�rR;o�>�uG�����`Q��jń�D�����<�?16���-�K�Ñ=��c������#(X�,_!�FF��3<�91U@�eہ\>#�=���բ�MoC���P�-Q�Qx҂΍P)�xܦ�.�l�J�"㹷ONx����?OK���Z7G̯���q����{����O��Cײ��Ts<�Cx��(�J��TZ��+%�e� �y1� +AT��A9��0A�4!��9q���1�j1���D%��S��h��f\���~�
~�%����������)lP�i��������Gn����5k2<���A��'S��g��V'�0@Q������*	�F�T��Σ�u�<ႧxѽSt�đ<^+����zA�B�L��<>���� ����0��4����d�+6o���g������r�L�$w9�-Qq���ĝ�؆<Y�P���x����!Ը�L4�߄g��R��Q�+��"��Jr^Tdlk�f�~V|o%�&Ź���"�k)f�����/��7��O�8���f~,���]�N&��ɿ�:8p���Ry�m���V����M�Z)��xT/��[i�&�\��%Fs"��V��n����A_��M��5E��4"�Ij����!a�N�b=}"�Х�
|�r���FD&B&�7Ԟ�Vh�F��*���xp�5W=�t�Ɓ��a?��54��N����Q4�[\�]��M����S�l_	��RC����/�Y���fcY��3��P+�$I��	�Ul>�܉���Oe3��;v�9;��'?y�4HjDV���TiBrŜ�	�ðQ��:�'�	eR3щQ�	c:ƪZ���f!��x�����ق��6(����Q �D�䂛w�tL�-T-�+��k��g���3w�noo~
>�6�8`~cv�������x��?3+�ͺ�������H�A>�e�i޶~3�%i�R^0w�:��>yHDP�"y
��R�!M!��)��*�QUCWEg<��mjk���KD�!Eo�h��f'�'`fz*��ՏE"^S4��C�+֯���mW��eǎ	�;ZZZr�t�5K�~�9^;.j���_�]#���Ku��w�9(���z�g���p�}�/���5U\t]OLM�����O]q��ɟ�|�P4_�*4���d⵬�A�hQ�و�؅��6���6I��Z*G��[j �u����H�¨悸��d�6m�򐸅���!1B��1-�N�H�X�|������ӹ����-ZT�� ,�_
><x�t���<��cG�|I���8ĉ�-�qӍ��@:=#F�d��P,�"E��d�k�4����0���΁�Q�WX<HtP�c]�7���"M!�uuAK[+(�.�f2i��LJ�<�����4c��YUU����k~���z�n�b1�B͡��x�1��7�.���DqQ��[�����{'�`�ƿ�S�u�͕��_%�����(v���0>K�x���_�ⵧN�znlb��d�2-1l���#!�����D !e��	�DCN��Rx���(�Si���H݃fh:����B^T�	jb*�+�Z�&j!���<ω����=\~��D���cj������;�����?�����f�Q�)W��Ǫ�*n���'ρ)��l�� Ӝ��i):�JےV��t�t���t��4��p(x��iZA��+ ���Ǡ���{{!����BXP ��� ��g�ÑT3��ڛZ*��nkn~bǎm?��w�.�Nv�/�@����4����mh�/C��{��*���5~�[P��h�����ނ�b>t͒'³qmR)�U�/������[��֞l���"]VTJ7�������8��M�~�a4�4��dG
��z��k{x��-���~NE6M���M����,�!�~��\x���NR�EV�8M0+���N7���]�fz��S��qNqd�����ԩ��'~���ǎ�Q�T�RӴX(�(�F:T7 ��S	Ԅ�~c��r��94�#A��(r����g����D4(K[�ѫ8
��3��wQēI�E��''�a||\D{��ш����D�����_}�U/�������q���ڦ3��gM���� �F��,T�^��?j����ԯ��؄�)�:�����F��hFA�xݫ��r�֓��?��Gٗ��C�X�C!� �y�c�"Ж*zRZ$�
u�1�LԲ�����	l
F��M�8��I�ſQ4��j~-�!/E.�#����U��MkEE~�/_yi0ٓH�M �̃��9}:�|쑟}��7���'yW�m7��%��Ho�(���%ciO7��/�_��=7z#W(b��<�t�bh�5�7=�g1��H������Hih]�����"����X*��atd�3)��]�ns"���_[����[o�q皫��qJ���cccx�����Pr�׹��9N0� I 	�Y$MQ��Dk�D�lY�]�ػ��>gw��d���=��dJ)J$�� &�D�����9TW������`8����<�驪����w�w-�����f�<M���=�)s��@��W��4�s�/�5�i����$ЪHh�=놡'���UÃ�����oӨ�s\�jq3��
3�c2p`Wm(
GX�, Z�	8S�MW��X׉Qk��*�-W�x־+�a7ʺ5h���Vh��oA)��aҚ%E�M}��_8xp��+<.ONx��x���j׮]_w]�JM�B�d�#zWR���&&&��N���	x�
hDj!_�����,�!��1���z�)=!<��Q�5�̤�I����C���Q�7�F��x�SCP.����x4f��*�g6m��Om����e�޴��Lh@z�{��x��!������?Wja��F�������4�A��sE�٩����0��j|��!i�W+e���m�׿���\����I+�+o�M��rV�X��@#*��@����yg�6�� W�1@C���w�#��ڠ6O�[��s,bA5?� �,��5551�N�J�y] ]�l˽��ɓ[_z驱c��K���'3����������#G�QU������8a�2s@E�F<��'�D�k��o'��=-�q0�T��q�5R��E�A@��)�`.Ԕ2MV��k;���Np�A����gs028 ��)0�{�#`�E#�ϯkJ�[�q�/.[š��fo��y*�x<_(^�,WrLK���*`�Y�7���2W�!g��0�y�F�<���s�T��\���y�Y�*�j����}�+����������g��ѐ$
+�%��q�Dj�47 �A`��A�_g�4�ltԁV�Z[�!� 8�녊}��]�m4^\S�h��T��K�]�Y�UR�Zշi���c��]9������O�IPq�����e��F6��Z7�H{k�g@!MPm�a��ZkOtL�G@�&̱v��O���K����yJl�z@�\c�|,��2��Q!�'���M�&����(>N� =>��B�E�"�{��Z���MOn��a�2���h4���(F�ڶ���jܬ�4ڳyQ ���#&�@Ñ�ㆁX��<Mot�R��ܰqÖ�\n���/5�Q��P.�[}��hh�� 0�z���z�E��x�M�%���?_ E����TQ�$#�f��b��LhGCl�T�2���E��y\{-�c��Ύ]'{{��L�'��<9A)>��k�v����Sãף��Rȟ��EY�r�����L�ͤ'QШ�n���d
�,�,���@�X��Ǔ$��&�C�R��-)Ik55CKk+�tG�i`Njb��FO�SթF�M��զd|_s"��[?�O_~����}r�Ax�l�f��w)����s�ϰ�UCp.���Pcu�BX���Ԛ0�� ;DB�����n�n|,��^|��Z�X:���c��������Z�C����˯�`Rˮ�9�>���B���{���j,8�����A\���g�U8W Ө�'e6�E��z��'n}ᵗN���/��q��x2��"�_y�ͅ/��ҝ�L���Z� �4Ԉ����P�qǍT$�
��,m��1���8 �0�����C!Vk�HE��ӊ���������l��%H���Xj�
��MNS,VD}��w��p��ǖ�[����>yR� T�um=��~����S9S���ɹx�g*2�y�3������t�8lud�����drխp˭�j�����������p����w,���"eHӘr��p�fh|��Rn"�n�Z#0N�6I��4�T��EAv��H$�p�¬e���s��D,x��6p���Zu`ߡ���}e��^o�x�O�#G�۞{���LM�o/JݡP@��l�+ f���$�i��%�D���q�z��>�N0-s���>f�} �e�F ��5�	�$���%���\���k�.d&3lp�Tz
ˁ�d�s>Yپ��e^s���-_�<�|b%�e��^���;�Z����Ň$�I�?��/�)�1!Ζ������1QQ$W���B�~��u�&�|�X�/^�h˧o�퀪i���Z �^1�(W*��a���y��b�p�bm���X�Q"�C��PR:a�1�imj�A��B��B�F���F���Ǉp�my	�4(ҸSCЁ�'��~�+/�xtq��!��/z���'g��a����?\;1>�y]3�P�ȑH���?�Q��9fƞ�U���V'@����e�ުH�� ���R���(� K��,(�t���fhi�fT~�`��l� #c)��Qↅ�椃Ǧ�>��+._q߭���jOO���>�B5"ccc�B��$>O!��|.:q;�v����\�Ϻ��sKF�|RԂ��gy�9�d�-�� ���/k��ַd�7�x��o��_�j��d�W����E��
���N1��29����g�AAD���Ã�e�ch�M���}~�EH�,0�&]g�����.%����S�#
��`,���O=~��1��{��x2�P:���d�}_�2�@�%Ʌ���\.���0�E���Zk��h^("I�H��R�hF*$�� �0 ���%�Æ�2kii���X*�66W���4�� ��0��O:II�D�ϯY��g�m�����U�B���v]�i�&ovl�"A3#�(�٨�2��ώ�9����H�k��H��.��$|��4D��ժ��O�/]�f�pM�}BӠ_:������dv��r���s+u2 x�dкe������LjS��]� C��G�<��X+$p��Q���3
eZ?T��P�a�c9��+�4h�3�')+�p��}��}�ҕ/ⵎz酋W<p������S�/���[��ac���vww�}���LMM@���{6�|hc�y8�	OS_Ԧ0����P�Eh A�Yޔ��:�a�GD%K�	�J TQ4�&�����(۶5%�ONE��'֮���oڼ����&s�T�vE��2�~q�G�9��p6��ٌ��s�������x�2?�P�6D��٧�]��9�2:l�ܲ��o�X.߷h͢�^x�e4�[�#7��-K�m��tH�AQ�#1	p�N��'�@�����1Xй $EdŊ�|�Rdb����pMj�ȁI�RsS���8j�9�Q9��g^��ݷ�><�xrQ�<9Mhf�Ν';_z���i��)�R��6%��
J�w�z�8X�����eT\�H�&z%T@�q�"��S�F�� �H@��>f�y�hDԨ>4-��.�H�|�0�Aҙ<>vʙ���[�3,�c������+7n��M��p� ������_�N���~J�J)�]�]$����8���-����ѧGl�N�	���]�D�?���&���4Z�qE���M$����_:���w���{���s�;��SA��D�ӅRi���~��8N�����n�I�@�/�HH6ہ�w�>3S�
�a#p�AC��ń0�1(�� #� �Bu?<��6*"h��E��j+ʟ����\��^��A.B���'�ɡ���o^iK��~�P�w�C!Vc " ��>�L@Mln�˭ԙ��N���x<Q'[ӣr�� u'P������ĺ�uk��0������/���!5>	c�	6�Avl��f2�|�]�7ݷb��}<v�>R��/pm�v|dnA���$���4���}v����}�{�s����Z�A#��
������g��_��O�V�t�}nY��$���������WG�+�aގ׸�X)Gx�f$ctMAOE���&����$�pj���L��F��"�j�Z4/�cdd�Db�&���m�+��� e��OC��b�|�������{��'�x���i!��x|�?o��r���dV+��fYĀ�lt1�}Jcǭ�:�n��0� ��C
���P�4��-@��FU���ԕ�J*�Rg>��@���b&�'3�8�G��OK�Ɵ\�ڇ�ذa/�	\ B��b��/��UQ�Ÿ��0չ���i\��|�0_+#��}�
���p���9��z��Ӳ8|����/_��R&�7��ƽ��?���/�?�\.��oUl�Ƕ������u}Ӝ ���A[�\mD:�h�`늀:q ���P��10q}R���:l?���+
���,71>����[o�X���3y�.2���'L(��«o-޵g�g-��dF����#jVRn�t�΀X���x	$��&RBTkP*Uj�PA��u�P� *��p��B�Q�c���@<�V����A5m������L������cQ'�S����V�]��W]��kk�[. �T*M��}����-%��F�|�$���LN�s-8�-�sPd`�ɐ��5
q�k��}�e��[/����Ͽ���z׷�]�ƽ�0�瞓�!�t|X(j����V��m����"sr�E��"z��@��^$c�����N�\,�لSA�Xd!S�WY��͟���I~�����7����!�<"��K<p�	�#�tp��oo.
7�����<u @� d��V|\-�i����+V���:X� ��1��\4�:jԲ�4m�K<47ǡ��A[;�bq��,�k튙���ɦ���Qߓ��Z��5��G`��\@��W�W��ތ���i���y=�����>ϙ"���F�5�,j@i�:K�Q�o�*Y0-kQ[[�/[���w��g��o������!��}����&�|6{�e7���J��9�
�"E ��cP]��{&�P�Aj�h{<akZ�x��AVÌ�ҁ�nu]ר$�i:�j�r�;���{i/q����F<p�	����'oH��>�ƽ�D�� T63a&''Q�TXg�H<�|M�V(�6Q�6QXmA�'�FbD�ց���zOlZ#�O�<
���B[G7��M`sd�yM����
Eh��lY��D$��M׮�ﲵ�y5�d�Y�s�E���pB���H�4@i��fG�&�*��Ԩ7`y~b=�Ghm@ ��Ѹ/Y����֯\�F`�&�X�=�ޫ��W��;V�eW��7R'�cY>�vj  �Qv��Q��"}S���>�AD��b4�
	 ��a�^ai�bEeQ:�(Q<�Ʃ[�e�]'O���k������=�x������u�ݹ�NK7ע�
F#�!*����t��E��Ex��V�R�a�u�Z�H�RĀQ��CL���2P����h$B`��]��;�B��N���8��
��noMN�«�7���m�7�z{=`p��$\��`#��
H�d��"'���L���Ff���]�ـ�N��|��L��qjsl�e��m�T4C[�������d�A|Q�"P�׻� UFR#i��Ԫ��f��t��CAF�L�H��zQp��=�``����E��em��P B�{����a�� K����_"~C��ܿ�-;w�<���O.
���E.�������۹��1R��i,ɼ�B����8��b$��*�Uu�!�1r�A1~EfǓ¢��Xl<3!�4*�dS,��d[Xhr�*L�O���(��+����Ӂ����W^z�m7l9�y�V���,d���ك��B|��%}p.sf�	ӄD��5��X�_��.]��x�� Fm^�k���S�Y�v]*;�����zz�����`��U��\�\wk�Q���C�����X.A<�L.�
y��,1�O>Z����l��a$ _�LS�ӽ2�S��~��'�߸{�;�⵶����/8����|��5�_(�*=�H\�P#)�b����&i��T�:���F��jh�r�B �ʶ7�X�b0~�<]ţ�!Ԯ����NT�2SB�Ccp��10�\`N�-YhN�__���t�U�r���.���T+�-�^��w�S��e;	|6�����F~v��iE�g�7��쀘}��=�vl���kk��G�����N��65ⷬhZO4�}��i�7o?3�'�{��;��|��G�c��թlzm�ZI�M��!���>��4BA?�߂�����6=��h�u�Ba
j���,������j@ׯ���;x�Э�{�0��8xr��.by��񣇏܄�be�P�����R��j�qMU�ӊ��>M\����AY�QkPm��J'Ќ��� &�T��Z���Z�;�tyTZ6�� �ɳ��9���5�\�a�C뮾��Doo<����zQ&<	�v���v;����m�L7Լo�L�s��M3��Di��g��L3�Ck�~T���d�i�W\:|�=�<٨? ���V���_������ş��|[&ғm�y),��Z$�N���:��#pN�F�\_����V�&���L���S��H:�'�����~͞=�_���y�H�x��"��I7�m�Ϯ���܈ʸ��|f�яQ�(����X�Ljdݨ�\���L��Q#g���~{1�N`yU�*�h��$tu�@K["1��x/Sp�����A΍E�Z4ܹf�ʟ^u�u/���UI_$�ϒ���x�)��6i��e�u�h8y�FV<s*c�)q�9>��3�Yy��@��b:-�@��?fl�hm�h�kJe�B��>��/X�����V�!x�{�'�����w����������x2���X.���C�0G ��,�E�y��<[�D�������>�@��
"X�׹%Z�d�~�UuAŒ��]�oߚ=x+#��-8��ڡ�}���C��"X�޼H�����A�R	�Ji�WS/2`@��6�̈́F�4E
(bШ3�Bc�"G�	G#�����e
A�R�t6'O�bʀk[��ζ�=���f��g=`p�	U��s3����"��W�9[L��z���%|\l� ��{��9SsF��S&�v8\[a�u�^��?��������H��:v���屩��߶>���J��j~���&JP+$����"(�+�u/� ��Y:�R�D�D�Ih][��e���ٿ�5����|�x��"��å��{��5c.�p0�D�c�~
A�"�0c0T3���h[U���R.�|�sD�BdITo@�	)�1R�x1����4�)�hbۨUqphғc��ez8�;ҳ���n�ܯ��Y�O.J��N���/u�C�ao�m��W��D���u�҇�3q
�)}Ј ������������'S�N�h�iS(���+W������?����N���v���hJ5,�N<�
�>CӸ(�M215R:!
2�NM��b���t�"E��e\��
�-1`/ID-R4�88�o�[{�Sk�7���\dB��G}y��x�:�r��Ѱ�
�k�z���F�t�U�5�Ivd�x"^�1�HWP�1@0#7�����:ēͬ8�fΧ&�a|t*�3x�Z�t�/���ǖ�Y>�)��[�)�cN�y��c�����D�Y� ?��~��C�=O��s��3�G�=�ZS�'�2�Cl��L��jnn���V��;�y��f_���sx۱�,ٱ���/�spX�O�1(6~W�"�.s �>�k��e�N#x�8����KjcV8��bS����|}êeD���'�x��"���x�V�v�E�O��"�Z�>�M\��D26��7ڜ�
�Z%}���G*b���(�@�eO+���������c�ɤs08x��YU�2�c7�4M.ho~���nxl�-cޠOH�9��q��+��n�F�q�qsdf�����������\���B�4�3	�Y� �OT/@��8�h�W�/��j1_��$H�)ĉ��S~���}��`×}��|>r��h}A`�fԒ^4Y��u.�Cl�#��@�B�MsX7ݫ$ɬ8�49ɲ쾣G�^y���Nܗ�@��)8��2���O�����I�V_( �B�уC/~r������A ��+�j �,IQ��d��E`U��^F-g�͘�H_J<��l.聖�%ӆ�L��� �� ��N��/�77�yӍ7�r�u��X�<�)\WA�Sp���� ���bͣ=�Q�0̉g;v���4�s� �y�s ��O��7y���S
���#���X��X�yu��e��t��k�̔������#��p�L�G���T��bl�a�:�cZ�t]E������bȌ=C<�d����"	�H�O��o:v<5�Z��Ё�������O.8���E$��ڷ�З|��� 9�શ�X�B��A�P�JYC���Kl���|�R��*h�Z��T��A����1�5���Q[:.~& r��`ɢHDc �2;��T����\Ƀ���D$\Y����-�7�|�ƍoyEN��%�x<_*�^��#��z3n�EP�3/E��1��ϔ�=���5�[��l�i�M��cp2�a.6G*44�VP����D��r�9��f�ڕ��K��Z��\޺����l�[_�ֶ�����T*_�Kj%�߃#zR��|���@�AH�lSkS3s�&��JF�e��8����4�\�W�ڱw�ƵW���f��N<pp���'�\[�T6����ēWb�v�b� ���?R+#�?Efu�Rqzv���eI�h��/���;/��B��8�rF7�0�6���	T:UW���2�P$�h!Eٽv͚�ؼ��6o¢'�H8���rO�����V4xm"��9�y&/�\230�K=�|����1��\ a�m4����MBzr�#��|i����������������Z���w���]�l6�DC�����*�*�"�&7R��-���a!���i��e<	��@N��k��O�gE�e0t=1��^ut���x�w��N<pp�ȑ#C�ǎ���N ^	(l@R�R�tf��M��"�4� $@�U(�Ҍ^/�`�&�qHě�@m�o1�7J%�V��mmn���E �B`	��eH��T:���ۖIď�߰�W��ly�g��"x��Y$���r�G-Co�l�N�\����?�y�}g��G~���G�4�gjc<S-B�wJ�Qka4�Ы_�`A�W7�Y7���qbM<���}�������>�X��o��F�kP��W���>$ޒ`@�D,�
"���^�J��E?�`�ڝ�3|Dشw׾��}��)҅&8�����]���*\�A��Q��&.NA6�� /�,�w�O��7Q-�U�7p���7A��`$^DH��Mg�Mֹ�;6�)<�l�Ύnhj���t.'��app ABױ����W�z�n���{�/��
=9�焼�}����.nZ�/��c�
�������T8Wn�����T8[���1ä�9��W����t�UW�G p�N/0��a�9�:�d&�D�4�U*�0�I�yf���>#���q$�)�8LӨ�%��@��
*Ky۵���z/w
<����P�#Cm'�q\��I
F���f�y�Nd���P�|
�$6��W�\.��?K�ȒZZ���$�!ϸ�yQ �4�	�XS$=����D% &'���*@�W��X(�_���7W_�����Wz��|����j����k��n��m[D��4�f`�ӽp��;���3y�s�\ �\j�įp��ęכy����:~��
�;	�x-�{������������뷧����玺��Ԉ��+W
�.򌟄:���X)�P�M���Ȓ�� ۟�e� 6� �@#�	4�,JW��%x��7��\��J����봪�֧(�uA�A�T�B�Ċ�C�����
��EHQ�#AH$��W���aS��e��l���A4���vX�`D�#���346�FF!�M��L��BeAg۞��|𺥽��O<�R'H�p�s�f.���}��:�Ϭ9��0�0wZ�!O:�Z���4����(�O��l�r}ꩬ�m6p������z�o��oK��Ͻ��S�_��S�cc��i�W�9@�^EС(~�wj���0Ȣ����L�	_�Im�Nmb#�Z��Ɂ-�N��3Ey����B^�\�?L_qq�H����͒��E!1��jԩh���<�s����� _��C���T���h�!�LBKK��(2��&z:�K�0���,vw�Cׂn�$�@?�/©�1HONA�Xpީ����j���nܼ�un�����#	�Jw�=��꣮�-��rn��}-B���C�QCP����\|3�f�|$K3�͸�y� x���Y��!d�	�7�T�`膄�/[���Ս�u%Ϟ |���������-�rR�c�}�J�J �-p�H�9�Tf�}rm�*E�〦�H!�
GX�hC��F'�&6�����x�i/=x���: ���
�2Ș
ZW?�;B-�#��T�,X���~W��l�?lC�B+]���������SCB�=��U]��v(���U+ h��0K9F��/�2Ќ}r�X��%Z[; �H��XT/�Z�,Ӭ�jM�	�����A�)	.�B��iH�M�Z*��ٞH\zɲǯ�j�k���2x��o!\W.�Jo������v�D#�Y����9�g�g�8Gc��9[�`."���X?p��s��H��0SĎq���ߚe���T,3�W��{��޼l��������km���s}닅��"P�;' P�=��5#�ԉ��ڧ{ � �tF6_�J�򒑁��'&�'��\0⁃߳�����鴢=�JT�d�L!��*q��'M����-�6���v�23�W%Y)�~Iw}����"������,��<H>��vnp�V�X,��Ɲ��L�C'��NB��Ate��-9���T̳9��Cs��A3�9P!%�T���1D����Z�Z�w�T������b!��E�\ڻ�śn�ԯ�m�0�y�|jeK��s�k-F`�D�لF����!���-%0��h��+g��W�����^\-����I�@uR����c������R�Bf�{ ��<�$����)���}�����Vz*���������Y4��
4��"�B�r���	Tt*j�����H��Ҵ�P�O��)5>����^�}��Ura�~OB<08�_ߑ�t��2]F9��d2]�i$�K*���Yn3(h�̛� ��8�iAr�k㚴]�'��ٶ����,t�q4N����@�T��b��o�h[I?%���7ѹ��a�T�P.�Y��Ԅ A�u�:�
D�"Q�m C�����Ĩ���м��d,Z���{ 
�ɋP(�܄	���X��"{t�~��M����ī3����6�q&�G4�(�p#��H}̴�s:g)N�����{NZ��{m�;ꛦ� � ���e4'���/[�"���~w�O�=�"� ����o�ɷ��w�@h���㉗������~4M��*G���9�4��:Y����(����NI�x|����>��o�x���\�̅O�x��w,�P�����魌�_ng3�����@[�璢�[m�l]�C��U@ϝc���4��Z�5�S��L�$�	 8MP���y�P�Qഊ
��B*�$���~�v�BZ��D)�<��<�i\3��h��!F9N��X�G�U0Ћ1��P�)���V�\�1�����0�
Y�b5��_����oڰa7����C{�
W������Ռk�J��g;�zڠ�v�8���CfF����BDԗ>�(�x�$�.�]5�����w�����=�af ��n�/��/��B�J��V��ţQ���@���H�� 5(U*�un�e��Ԝ�s�TSG[��G�.?�pE�{>�u!}���#��!�����>x��N*���[$iQ$nA��7
EAW+\��r��k�7&Ʋ�� ��\�B
��~��(l�&8GS9
E�$�")��)Q|�ӯџs�T�۶ E7�A�l�
�,*��ã�ީ���ˠ�K��
>T�,�18��Y���$,Z��1!�x�2�7�����bv
x�2c��ЪK�o��-o5��{u��N��/���W�
�l�c��i�!i�+���Ε��#��랉ifN�_�y��jUAmqɂ�fs�c����; ����m�Y%��ٵ�_��w�^X,��A�	 ��uK*&R-Rc���d�?
�'!��t�4�~v׎=���H�'�X����,�`$�J��~�p����e�f�t�E�:�7�ɂ^*sh�Y'�&H��%��@,r�#�m�I샄8�CgA�e�LW�*��8Q��)�i���s��	Tx����� Z,��ףN"9��v��@$�
�Z�&^��hCU����&����![5 �W��dNUKP@eQ�]��*@( ��n]m��U(��=f�%H��C)_ ь��ڒ�Go��<޵|y<��w(�`pJ0�'+���]�O�\� A`;gE2_t�\x>��¼��\������K3� ��� _�z��o�
��1�sh�)[�jo�s�0������|6�嶎��'�Զ�1��q �}G���C����zQJ!���CGE�|6'u�u�ڶ���ǟT�KݷdI��iO�_����$��0!s���#vmv�r�uI�\>߬�r��2}�؈�݀T�C�!�1��A�R��V��Z����f���B'�"�^���#�2�CbC4�s���}~_�� Cb�^�)퀨?dh"\*����e����I�8ԩSF�4�Q��aq4#����0Z)�`��F��g����牜�Ao��ZEud�϶&b/^��G7�x�0|�}_¨�נN�
*�?��w�-�)�q�]��C�=u���:f�͖���)jl\���!0R'�2��9��&I�5�W��fs���st��-xrtl�S��O�B�&Y�9��ܔF%�؈i�`�N�f��l;%3���>|�x`p``�����<x�|�`>:~��MՓ÷��?���1fb�Su*�&�
�휃�����l&34D�h����.H>ƅsM�r-�t8�uD�w�2��:�)�c���:�Ԓ���7DĀ$'#�/�G�)�(����Ѡ#p�����׈�#�ɘ ��(z 2�~A�1�!��^;��LT58�C�*�CQhW� ��0�ʂ4�'�P)V\0]-��۰vͯo����'|��1�U�;t�uׁs-��ܔzv|���ޠ��N���{�(��L�7]��@}4��i�;_(��������g�2���f�l�xW4|�Wl��ѣ�mjn�mźUS���/�,�l���������d��\,mQ��$��R�y@t�4���
�q@��؆���R�ѱ/��?pr`��#G���s������P�O�x��\|B�����{Go�������Q��Ld'3,4�+W�Vd0�>��t86>
�3iȠ���:t�]N�9��[�S���4LS3����5˲tt*
����\��*�"u$�D�����r\��*Z����k�U5���b,�I�G�a�JID�a�4CS8�|E��Bo D�������D���A;Y-C�A�E-���� 2��TGG@ql*M�jiy��n������V
{]7�ԛV����>]��54���NN���>�����MZA����4��Ն�q�Aם��p."��3z0� q����d8�����!�ce�"��|Q���뚕�����,v֡f��_������l����Z�e�c���P]�(�P
�����Rɦ(cn��c&�MWh�����T��w�|���*xo;��O�x��jO����̾��Z�Z�j_V�
�ǹ��@��n�	�ã0����Y�
"m׽�F�j�z_Sh�'L��>�Ғ��'�m��X"at�uV�[:�D���uI470��ʪˊ\W:�����x�ٴ��ˆ�Ǐ���d4Db8$U�:4� �b���P�t"P�����Bw46�/�0%\��2O�eH�E���8*�	�d�K�`�� ,4+�h���77�~�g���K�lI}���]7�o�|��G_��5�t�&�-�n���x���tg������=���V�y�/���3hԞ/�
�</܍�u#Hrj�Bje�����f���~�/�a��i���3�{�}�-�@��3C&�ֺX/�l��;��,�()��e�vK��cMo��b�T��~��7��yۇ�o�m۶L����˥�%Yh-V����	T0M���(�P���T��ZMB$�rEgsW�UR�1Xڷ�;u�T��g���S/U�ᄊ������|D!`0�}����o��/��격S#r�sA� ͋�+v���b2��VX�tI�'*f�`"���ӽ�Poߢ��}���:{��ŉ
�'��U<��$Yg>cK�t�Ĥ�Գ��P?�i�2��e0��90U�H��Pp�@p�*�������.�B� ��d�ij�a���]������ ��%���XZ���tZ;V�����7n\��*�[1}>�ۮ��O?x�7��I��_�H�`�v�1����|�N��?��s��C���ˁ'��������^��,���V��7�-�q��#a.΄9�a�����:�<������+<j�'p��.Y\t~7;�wں�������*Y���&Ƴ�@��4>�rL����� �HL*R�#�x�|���_x9�h��п�'=�x��>���d^�~9�ܵ��>�fK]'�U�*��+O�����F�Df��\M�ɧ�~�o\ժ��F��%oܲ��S+�-+\r��o�e��;9t�nۋMTS��6��@7������	6T�vs�R$�8��
yہ	W�}#�aqs+����&����!e2�C4� �J�yH��Бl��C]q����p��tho�>I����_�B���/���#�_�}�|4���U�4����aqJ �ߪ������S����m��Nz����z����ﳵ����Ġ��-2+��@r�	���ؘ��5���#�a�󁂙�j��Q��s:ǻD#ݒL�o����_��߽�;�ϡ� ������-��[�q' EuUQd�jEec��e����-d�YF�D���ʍ���B��"������Jv<���T�'@<p�!�Z�Ww\b���P�Bq<�z��q�۞2\((~�}�0�YE.f���A���T<{���7�^w���>��S�^{m��2&T��k���U}E$����,߁X�'�Di��#`(䋀 I��E��۠.K����JT��)8V�CW:}�&	qh��!" �@ �錆	FހD$Dߦ)����j������z�nwhh,(��!E*<��`�����z�p޺�O�,E���͙F��D�4;��?�Oq��%���G�����/���x�xr�H=��^�G��r�iZ�+��&8�W,���٬���5�h�i���ps��L���<3�;�=~ �p�ŷŢ�Ou�v������s�?�łc򄴏�"��\�u%�R2T�H���3p@у`}�#�BF�`���QI��%'��藏?2y�u�^�w>��Bȫ���u���S��eN��V�9��E�H�6�=��8(�ڢ��5�(�w�H�ŵ7�}���ĪU���o�?42��p�E6��B4��� 8�4�U�Ё��k,�`�,j���.��Z�S�0LUr0�V �@р�.H��0��Á\�X�h���fh�x�8�'�b��u�/��I��L�ck�=z�`b�7ZV�|�ݳgZZr��^=�<�m�~���W��������[�|�۟���B�='V���M�J�uq���������K���]���_�ێ�~����>ߤ䃻���Sӛ��]��<.��ʧ��0���I_̪>����5}���MhDj�YSf�`�}�'���`/m����f؃۶m{w�֭�fK�g"���L6}=�h�Rb�X�#zQڀ:��
)z�G�L���B�kaɒ%,�@���q?~~��];�������y��x����+�����wS�t��tb��8>!�ШZ�(Lh:l:	�:o��O.�B9���W����|��o�����Ï����S�����"*-�{UWY��P��M��D�\��D/#�C�����+A	G � ��;�'��&�a�E	x�W�a�d�|���DBvoD1:�>=.ܠ�"����l3( �v�v\s�ĩ���o^�bWSߒ]����ѡ~���(k�,�ߖ���g�>����?�͊�y�����$e`���u�;���S���s�,Ǧ�RȨ�?�,�P����?�o;8����Y�伐z�b.$�_S�k��*�~��g�Noml�>W���ƾsdZ<���>��{����,���j�l�O�.���  JҺ�֦���������\�\-�Ǝ�r��h�� ��d��b���"/Tc�`x%�@��$�Ρt�za�(�a�̪����_����k�y��<���U<pp�����{7*��]f*ݗ>%-��07
�}�$L�ɭJ`(�@�.ko���'�����7n�<έX�;�Q;�+����Tmy ��ɦ҉�X�Jm�҂�^hZ�\f4�===����tr�h��Nq�\�cҙ��!��� Gb��WpT���Vt�p�����%��m*��Ŵ�[$�5�q�0zfA�!��.f�m���uC'�n<Ւx�m��W��_ީ,_���V�\#	�]���D��v��T�����G�ٰc�X`gnl���}_�Z���4.f���x;�FE�sEjW@P ��@%�Z��ج�2n�R���a����<��X�/�p�H�� ����:-�n���8�y�ȏ�ܙ�~3y��l�g\��}3��| d��2�z��Q�Y5��s9��l�hmz�駟����9��;�t�:q*��0tc��V}8�pl8��sRĀ"lH:�c(�P*Ո��G�D�D��P($�?��cOO��]^!�y*88���'��0��br��+<��vux��!H�&p��kf�X)<��[n~��_�➦��*��C����T^����<��!(���c H
踽��>�²K��TU�P)�
���l�$Ƞ
t�����0+2
F� ��@�)	&y����v�
��.:�����}�m�_�ͥ;v\P��IA�
��'
\De�q�R��C�%SS��Gv��\v�W�{��dNB"Q��oEi���u�ᾩb���~_.g��sOr܇�D��`�#�_i�w]]��x�yI@�H2A�9�'Fu��`�f�)x �)�aT����
�}EJ��3�ડ����~� @���0�$�=���CUW_�k�:��\6-0�sg��\DL3S	����f�<�^f�u9q¢X<��j���<����=�ܓ��G���FCO������=�t����C{k[���t]�$p�cC� �x6�$������<1>66�R�oA��w'88�����zK���Zu8t�H���a�z;�' eih\S��a�R���o��C�o�+/95�)��SS�y��`Kd_=�L�Ɇ6�Z-��S$X�d13��ã`p�Kr��� 4���6�а�`��z-�H&����D�/�����m�������Ӿo�����o�z}��;��2�ɭ�f_���bR@�aaS"�j����.��|�w�ܿg��+�_��W$E�P�n�M��e�����K/��VUW)��(��?��܃��S��'���|ĝ�����>;^���R���sL��ī�zxT�:����0��Έ���5�DAϔ!2�q�\~�h˾���m�/+����8���|�w�R������d��/��`8-\��Y��:�.�ɠ��~�(�\��߾��4�9�sL�j��ԂB^���p8��:J�ⱷ���Ŭ1��L���Mu��p0�
e>����M��B}B ��4�:u
t�X
����c)�l<������_y�-jo��y��x����ӫ#��-�щ�a�4�9	�h%��� �LX�l�駾�����a���ǟ���[�jy�O���@T�"�u�J�1�ybXF�g#����fV� �(���&�(.���$l\��x��}p/��9(P8]p����Hi||R�tuw���G�>�-�������Z�^=�{��{�ygga��G�}���T��ɩ����pG�T	E^�q���ȭ��Ė��SK^���l^v�5O��^�:~�A��P��C���t�ftA���>^����x�[t]�A��MN����������N��|��w��{�p��6;��`��W���v�ABԉ�Q1�+0���O�g�e6�ҭW���w�����JI�E���?��G��/�^�y#�l��_Sl_��[qĘ�ȣ%c�0�q�?s�ځ�j��?�������t�!����#�@�u�J�]��]U�*�쳝7�Jّ@x@���,Ӿ²,?�P�"�Z�W���E*I��M��e2�d��i`l����¸~7��������c��@�G⁃y�E�N4����剌@�"o�p�*¾�a�d�Vdq���������7?���[��$��'Ƨ:���B�R�S�3�r�,��
ˣ�a�1P�]v�%
`rlD�ExT"��򈊬@��	Z;; ����Y	C��
�CHe�\�1撅��¥}Rz2��Z�����/�y:_������|�[�����u���:�=?tr���}k�lq}�^�jZ<&ۜ9�
$���H����O����w��{޷l�A��#�	X�����/˂�ϻ��Upm���r[�\�Y�������Ó/;�,Y�A���O�S>i�dI�a��T�M�v "��f�
L\)�������CŇ���9Vg�r�5�4S���do�LV�o�������+-v4������ێ���K1�?�m����Jfe�~�1[8"�6��HA���AM��`J����X����B�t��Xxv4���2>�\�T)�U���,B����	*��j.kf�ZQ7g�TxH���L��wPf�H~���A�����պ�B�dE"=#T�Z{������/o�F��-�'�x�`~���2.Wޘ�ٶ��u����M�����E%ը�Z���m��ڷqK��~�c� �R��xA�@�A"�ި$�\ UXЫX�$-Z}��`�CǊ�X��.qP��8$[[ ��&�e�<3E"�3y�:r�Df��-�{Z����q��CG����_��Yy�=�[�����ԉ��_K����c;w\U��QYuG%)$�ʜ���Um�ˏ5�5���il�ž붼���f���Fx?)l�w��^����*���$b�-�߷h��.:#�o>ֵ�� ��s�N��Ez���h���#�r���B���]r�᧿�$�A�`���j�X�@��ש{����� ,��AF���銠��%cj�����,?� ��!u���i�
�g�������f)"�M;lD>��!�smM�-�����R��'یѭ��qO$h�U���UU@o��tT �k�D|�P,L��d�
��6tM�Ћ�ST����L۩��������G*ޥ��^�u��:|��z��cx��x��x�`>	[c�˝���R&+q� Ղ�,LK�hk3}����}�Ͼ�kɒ%���"�B:1:6q�OQ�iq� ���@� -fT��`��ِ�|�P=*�g���$�!%"�8$�[!��������+~(�(�8�a�ڟ�������_3�M�p���ݭ�2uc����M��W���w����rZ=dH���:��o�f���:�gύ�\e�5K	��b"�o�����C�����������o���3ӓ��A� B`�Hʢ	�"�`9�-�Z���s��1�~k��W�r���-�J$DS")fR ID"��A���9T��{�����1 �S��h��UU����M�]��?N4���nX1�%L�@߅G�������oV�*�NB�͘��8p������L��:rp��у����hy�T�<Q�-0=���B�j��9 (� k]��1��@
���I�A �}��x.
kԔ��7�hWk���鑻���2+��=�ih��>(��U�]�J�	C3�p,eI��ǆ����ٌ� g�η�>ּg?��LdAh ���@Y`�˵Q��k׮=/��W��U�o��oO�>X� J"���H�� �&2$+�7�k�$	���'m��5fX�V)s,���*Si#�%=����w���#������GMp��F�>G,V��d�)��:.��]�# Ɉ���[�e'_�r�G^���۪c���SF�X��LE+h���*�:*q�7����nªuk�F��β�M�4,<��L�������-����d'�0�˱}��ʋ��t���׮���^�'V^�a�_�׿�m۾���.�j@����񞺡������B�_Qн& ���N�o���_��ͽ/<�{t��O΍��Դj�$�I��u�_���_ꪱA��$N�u�A����lI��E�@�18��a9����Z.���&���xz����D���xC����KV�xzj<<Af��r3DQe����I�;�T���[d.g�V�c?�/ro^P��5,U�������/�u?������יm�X?#yQ_-q.~�m���-������¯������<�L��HS�Dߎ[�*��q�뎎�����Q52�k�*�����=%3����� ��;�y�I@�μtoj4�������v��ͯ��w׮]�Y��I��!Mp������K�|e�W�GeE��i8Z��2.���>��ĝ������'/�����Te.'���-��M�֠P.A�V���zڠ�/A+��hi�BCE���<�a?�X��:���7s�Y�0=�'��5��[��#�=����G�u�xl��=����Nly��ϬYs�ꖞ����h_<��[���������ǟl$Bϋ��ao߾�/�|���+;^����+���+�e�Z�xkW��n�z�ˀ:���O����ȑX� UT4�oCm����m;��~�iZ.�o��[�(z�57p��\�o��}�Y8�;v��Tm.��B�/#p |��$H�s\�!�9�B ,�3��*9�)m8?>�x6�[�����[WϞ����?����}? �i��\���YaSM���~��[����NN�e����}�_e�fL�\ߓ@����(W��e�QJb>�uכ�'�N#8(��h'bX��JJ$C�ޣ�&KJ�(�V���T*�r(��mbD	��\����8t����<�ӧ
ccޓ=�bYrs���	�i�RڭV�Њ�����DL�§��fڼ�9��S��>z����o�(q�#G<����+�r��F�a���ێ�6���+ AX�Y5|�4}b$ү$L(ϊ6zk[�Z�8��y�M��s�����1�`޼�/_��W\���ꪕ�^x������7��ŭZ��E�8}�TKgO��<��?���u���׆���g)"��9���:>r�%�ݵ�kk�2)Z(Wd�"�ĀC@cZs�;8qM3 �Q�L�$F�R�b '�\�ZH�S鶎4�{kt��aI7X�I8�m3��;��/|�q�a��("4K�Y�J��g��������3���Z�2�K	|��7e�S�Xh�B�i�D����ޡla�ο��������,qP^~G�Q�Ǧi�CppZ�2):��ϥ�i߸���R�����N#l,I��~��L��*z��[��:g�3����'��Gϋ4L�#�N
<����g�Hj��q�U4Y��'Bp@!K� �{5�*�h.T�@�4�8�a�Dр)�\&�V�5][8zz��m۞;���ϽG���xo�	�1X�¾��v���X�%T:��G�Y��Dh��rt�v*Sv}�k�.�p�D*��bqy,���䊌�@���T́m�,�0��
�V,�{� �+�1n��Ъf=�qҙ$������*�ɩL�N�Q�@�\��c+V.}nن�o+˻���-[>����T�{���/['r���G���Hr���������]e���7b<,;���>O��ǖ����n��u���EI�~�]�%*\ʻ"��|WN�1�)�U�����p��X�h1�t�ph�~^5(����P��C���%���������0d2�P�T��h���dy�c���x^�>\԰��s�7�i�麮�VG)� y�@`���"^��T1���1��_�����=���F����|�U/�m�����r�N^���-�I��3������� a�ѥѷ�C�*u���9�Y�^��3����>^7a��Tp�m�����c �
��f'Ƣ�!˴�i9m�gi-�����w�GF����g;�#ѥb[�ƙ"
~oK
MR)5��,�&�3�0=����j�̺9����C1f��<n �M�ū^zu����9T�4��]�����/ϯ��ФH2�\�Z/C�5�u���M�<�pK�^��E٘m;��D�eG��*A�M$=Z��/f.�*� �s|=D�	E� �JB[W��4(�a�r�"8�RHǲP��y�������N	M6,�l޼����K/+��_���Prdd��s�+��޿��m�(ܞ'.�7zp4]��e8����o���%e�H���)J�%��]��jY�]��@�J]"�\��ST���F-��_u�(<�����I���- 1"��j�|n|��ÿ>�8��Ơ�c.�1�c� uv�E^ Y*V �$^�2 c%a��lN</A&;U- Y���IX�w�k-.^VO���{������6��G���Fs��h�J���t��D��R��vȀk A_�g�g2 ���h�}��9��N%���I�hM�y	D�\\o�C\!��{!��[ \�֋/��B���<��LW���)��u��$Ͱ !GX��r(A�r��+@�<��%)����*d2�Tj�8Y�B1��D*Q�7�����9�#�<�����틞��_4���>���\�P�X��¬k�d�g���?��2]sAR�R�f�p�ڱ�i��rI���U�+H@��@��~����a�ҥ�obG�cHX@�Nj��Vd��4��w���1J���Q9}�(��n�"h٪��Ss;)���{��'lӊ���u��u+�Z���XƲ��~���$-���O=]�u�������x,u�Q�[1���B�f��^��P��A���'eK#0�74 �}LH�F�Y7���K��Dbh��`�0-X=4|�]���<��6�.D{2 ���&��H���� J�E���� )	?�`��'%* 6O��J�u�O��O?~PT~����p��A�x���/�R�gF����-���x~�ip�;(���m뗍�S�+:�$�sR���ڢ�O����x}�<��EQ��b�����A��כ����B����I�r��\��8����2�C%�4���3�����(�J�ӣ�,,QM�_9�o��<��*���um��������~*o<��\���e'��V�V�ţ�5�9bD�����j�Q�%��=�,�hI3����ǻ$Qn��-�)B�𻥑P��J��� ޗ���YJwO�e:AVb05]���4��2���5
��=��_�s�ƍ�)��ᆏ�^}u�C<x�ݻ#+�-](�tF'�F[�[���O+񈔼��+pw{:��4αO�С��,� 3�	@�$	B0�LF�c�0�����T>�D��jLXb���"����$b	�Px��h,	�r^:x*"-�x"VA�I��g�3���%G��Œ0�|�$`B�g��,��3O��-���IJ��?^*~���^=�ǿ}?�{�j�"|�����x	�aTR���.��T�����Ϙ|�P�ab �_�7�>3��cv)�/�;=��g���TH?��Lrl.�D��o�%�x�������S=O�u�ĉ^#�X� E��~�qг!�@{��kĔ�C��g�����7�O�N����b,�@��ǽު���/m~��es'p
��a4��Y�6�yp$�i�@��+�hL\�h��T���M��ܺK����\y�y�1}h:Z���Ȳ�$�@��{
h�UQ�SY"�$��L�z���x�k�L`(�g:�{P���;66�|��8�4y�ٿ|٢W�5w���e�-�l��^7�]�v~y��P8��B>��{��?���}�S�\v�:I�[H���T�'Z� rp�<��fV���p��/~�įe
/ب�5H�#̓@J\�%^&cica��x,��0'���� ���_c�Q�z��mݐ��B���3D�(�d�H��
6��0F= �% ��11P!�|Ay�:8�d��J���xt���_�4]�w�@����˚L�ފ�r]�?2�����ރ39
��:�le/4N�N� <~��g���� $(
��!�S�=<Q\�C��u����r9gӿm:���/M�l!�(���$��Z ���g<��gs �A>?��Rggg Tv�����Q�r9¼�ý)��9S�ӟ��S��J���<����C4u��t������0V.��!��R2aqe��;w��E[�y�Rt��+K��ϊ�1���H!Zo�Ç2�I֡�����zL��L$Si��/�06:5��=<�kjәtj�����_�җ�/���=���Pya��{�+�?��ǿ|ņ+�eVEP�o���e˖�C��d�P���'A2>�B�~����b�1�M�5�"�g�p?A��]����yP(_M�t ��q�zd<~qO|⊵p��)͎�*)�B�#`��P
1��@�N�}PC�����qa?� `���ʖ������C�!��n��V��渨���yRN��l!ۍ_r
_�*av2 �3ig���x��s�&�:�>6�/a�A��� �x�FnQx�`��:}��.��	D�����x�V6l;��8�0�? �j��=h� K*{����Z[[X�p���%��z��(��!A�_�`Ep����=��{��4=jv4����[���^����F�s�2���������(�h�=w���Qo߾��]�Iֲeٱ݌��*�GIX8�M^*�DD������(��2�4���~�dZ�oN/H�(k���z����˰���嫖n�"3���BV��+~
��z���~�w~'y��o�4m+�(Wq&Լ�ի/���tX xļ�'^��~|�0X�4ǳ�/yEt���eR3A�U�2��;Vcm��2ȩ�G%�Yeг\�d>8������� ��R,Z:��ӱs"�JN~,�ߠ��3�8�,�#^2�Hxۖ����z�O�^�rl` ������ǽ�#F�H��}�։J���ܳ�o�9sޮ��)_��ɋ3����}B�?ԡ���zg�>��?I��9�݁��vuw+~���$����+�==G��)v~�e�\C��#�w���&L��}N��Lk
��3��*F��ِ`Tx��a�׽�ҋ�{z�Sh��{��&88�0E16Y����$ص�Pɤ��"�B������M��ȗ7mzp�M�_�8n��.t�y�3U�|�B�F�	 �P�Ş�8�/�Qi3�ݐx�,֗H�ٿK�LMM�����n/���{�,\��_�ڻ
�lܸ�y���Z���~�E�+V,���[o�V�N��謪�n$d���98A�Bx���O�#�B�<���������J,�@M^�0v}!Y)ט�£�6�T�e[�JAe�ǚ(y��d�[���0��b����I0�RJ���G��s��y��^�"k��(�I���<x3�H�;�51�V佋{�L4ݧ��.@�Z��E��q\{��=��s� �i�
�0����Ɉ��A�U?�E�=�3y:n���"�<:�/y.�T~u��ֺ�:� 8(��i�����0��צ�+�,�A	��gi?Ӿ����"(N�T���"~�����g
�aLN�>��Η(9q;�l�|�F �|�R	T��Ŏ�^�u������Zgv�8'OB��\Z4�;z��,p#��ֱ�Wrc���S�;v�r��ct�DZ��4m*bDQ��jV�@��k�e�uJ:�R&?[��v�o
3��*��PIu��YV���,���K����w���F��j�Y��]w�:��縸G�<?�
��ٍ�Ȓ�&��� �VO�(*$^�2Mj�@����P�콙�4~�,Y9�y|���1p�*�Kf�Q�E�p�,�|�|6~�����D.��>�,Gd�x�j��b4j"���$3�#`|J[��X/���눧!Q����NE=�j`�[���4Ǉj� �s���
%�^��&�����\����g{�.��p�3��=�����</6��<�p�����V�(�Z����ӷ�bv��ғ���;��x@�k���<�{�i�̀aB"���q��8��	�@���Eֵт��.8x� ��%E#p��[��� ��V�:	�OÊz��۱m�M/.XJ�F�9.���T:w��?�9�&��Ι��^~����5-z2?ͼ�	�*�(*)9��%W�h����N�T�T�r�����t��I�A�]�}K���ϟ���Y<�����=V"q�Ѣ-U�0>>ʒ/]��j�J���c���o��.��,�oѲ����]�����k"�\��k���������!��B�hp�L��K�*�[R�^e��8.����K�������cɀ�����nZ�CA�E�]�$�_<�.�S�߀�������렊����(�]j��H��ær-*���@�R΃c2*��!"'�(����%C�N-kZE�� B���ż^]�����$ߵ~�2�=·�p68�{�*��{����	���uC���W|�?MS�_FCbUGg�jhZ*�����_�Ahkoˊ7&	�M!;�'��g���>2L?\�@�c3� ]��F����������(�sR�c��Q<tMM�n�����h�<� �	�/����"D�'�WwvGn���jY*%"�--`��wq�-���(�k!����%1��j}zQk���0�ݟULӞ��|��8;mHڀK�,a���D��5�|� Bk*��$Z��{*�Fajr߯�O�tL�����j �v��6m�����ڜ�sow=�����s������z|�x~��� ����c��W$9�<J4�e�JTd� b(߽ʟe���u��|M��P�I<h�r'4�2�����jػ� ����H���"k��H*�bq0)�öX�Kʺ�A^Lg,C��D4�C:*�?�d~�Ei���7�����Q0��/���35���[:�-
��1��3=	���_A����P��{[j�ݘ�s��a> �3����9IܢE""�/�=�R���c����~�cm=mS�X�c{%��_�,���.��aGX�v�_�����gD4J	�T"L����Aͫ�ccz�)Ϊ������W>|��-[vPr��&a�?~���tO��"����Զ�F˱b�Pw|���ȥ=Gc��cOҵjW�6�r�Y�-�ag��S�O��GaB�T˟�eC�7����FN��Q��	h�9�&�jC�L�ZjmK�>o���~+j�M�n����j���N{G�'uCog�P�R�s�uviˮ<t\K�-���'�ì|Aj�x�X�AD0Ѩ�]��1^��H()��%^a�����S�!�o�OÊ�n���>���98���>�[�YR"�u\6g��<0e.�Ikx<(Z�ڐ�&�"�R��yq�7��������^7qm�L������F��� }�]�z f'��j��hx�]����>��	p��~?�������Q�Z���o����q ��szAQq�3��G&&'+��V� �H�(���]Z�W��&V!��(j GN��VѠ� 5D�L�"=cIȲ�k�/o�z��^����@�o<8��jS �^���U%ʒӈ��]�3!O��"
t1�eS��ֲ�UӢ ��EM��p]KB��x^�ի����Ƨ�^H ���FI#mRJD�qOJe��h[h�����遡%/�l[9�n����|G�#��%˖�O�]]��5;���V4�7`�Z�=��Ap����av�xhM�qѨ�Z*d!�J`]��Ae��L�x��\H���L:�BY�E�g@8	t� �	��\҉Z[�p嚅 ET����>��.��2��h5<FA!l{�'�TK���W�xn�/�:�>�!�rq�"��6��
/
�~����xj��x�����?pfE�L���G�B`0��C�%=����U4@��.\�r��s2��xD$\���4�E�?v�\��t�R���{����y�����'�N����%(g��pg��ע}ؚna�a����n`觼)
7��L�K!1je�so._�����ڋ��E�{����xp��rq��DB��ق��m��X�?;�0O�x��[������ާ�<���d�0Ҳ$�̢p=��O�r��u*�L����d2�B
�<Y��P�D�"XF�Ӵb5�J���w�Wo1�k����q[i]�r����U(��p�s��'��b*�*	�����T��0�� ���-����B�yP��#P"!$S. o��M*�������P�g�P�"��C�dѐ�'ׯgA�2�xrӧa�`'|�����R�!��@��p$O���D\Kxm�XId/̪���L��>D��:'�m!�Ns|�G:��t���^�W@ G�U��N���������-���]�0���A��0�r{� }.�8	���c��%ܛh0�r�B����i��5q����d[�mH<�4���{�	(��P�#�R���I�L�1���s/ޏ�0`��Qq��l��j#���/-߽{�G7�8��g��xw�	pģ�.b���%�Bqy�2�IkX&8�`��ENen2R4���W�jU���V�(^7E>z+ ա֬�T�m|��@����m8ڜx�`@=��\s�
�:us�מ���`w�Ȼ͡�F��a�"^W%.ar�g�9V��?w.Z3���Ჸ���rvFP8����a����B<�'A$s���E�\Ф�q��J�*uYD���e/`f�FJV�|	�9�3Jd��ֵ"Dc	(�X�d���;�����>?Q��DP���2P.�D�����6��{�g� �˵Բ�ņ����b���k=]��i\�m���ރ�pf���U3���r����xH�l`�ٌ�a5���a���e�)�p� �MDN�E�������0-�s%!{�ݝE�,�(;�yB�A��iޡ�"FXu�JE���7gDf@�����P
�ʍ�q/�0�4x]3�Q���3�؂��i�~��Mp�kRV�|�V��Z���瘈t�ik�2s9��-8TB2Z����f(o�E������'��M�L����k~�	r!R��6�QY��u�$D�^e���VhmK�A�gB9_�|v��V��,Z��]S�⹬|!7<::�/��(<���#�+ep�<��L&��d=q~��P �oy��g=�b�2ǐ�)����2���Q�!����17&	UV�����*N��l�b��	����)(���5��`�IK�χ��]On����
u�=���" �|�|?��\�Zi>�7G`����ޅ�Ҹ/ws�� .
\s'�1�aͶ:p�ލ/S��� �?�N6<�߮� �E��<|��^�X>�я��l��'��4�)��Ji��Ḑ�8��	��+�P��:墈�=���RI�go[�d,���
~6�88[�g�4G2X%�e���Й��F��U�4I7-<h�7*ޗ+�,Y��!�TK#�!��X�k�>��'�|}74K?���2�Xb���ަn@B� ���Yq��UXEE��~ZP�(K��y�j֔R�x!�
|�Rox)a��Y.���A�N��"y��@��~�0*I�@��soKED���H����T���vݩ9��[���8�v���a|��|Q<| �z��r�Z����l>��娺fz<;_�bRTe�?Ԑ�*��!���g;q���cU'3{�0<Vɠ��'D�SO�ٽS�Z
e�J4���V�Z"�oI%!�����G^���'
'�f���%Z���N���ET _�C������Ci� �2Z�	3� ��Q�������9�,O�Z��R���ZγNs\� �����]��u�&�I��oP#��# 3�0���z�g�L��%�R",�%J�&��Y����C��l�K��:���[X���K�A&�ƈ��b��G��AJ���AC]e)	PQ�F�w��I�H�.�D��}�$Z��Xde%��C��`��D"
����P��CT�｣j"�f�\�8Ν�7��O�,ta����0��ϥX�3�G�Q����Lݼz�k/�p$�{xA[[��}Mp�CV�%p������H��D��pC�N����]�<��ȷ�K�J%r��?��"d��L�a^2,�Z�� �В��Qs!f!����"���Z��RL��M.1	��y��N�����:�0���rʏV��*s��~ڱ͸Y�.�Me?S"I�m)O�8ʡ� ��y;�!�5ʙp� �
1"��<
�x��d��I ��(`|׬̈́S<�d������~.K������	��"�AMC.��H,�<-5G�s��m;a���%�[���@$���P(W@Rc,�󷉈*�@?k�kh�w�hc!�tRU�]����n�I}y���9����sp���f��o��=B�9�ǖ�4xf�*r��dyğ!��\KTD�Hu��'��'��G}-p��������������F��,��y��z� �i�/1|�
W�(f�%�;u�T�������B.?b�4X�눍РN�G!���<�4Si,a�=SB,�Il�i�
��HƤ�b�z�����o��}��un&����7�"{���꣞g�"���a��Ív��0���{�X�h3]�A29"ض���*~��6��n)��7��2�b��մZ�%̓T2�tZ�Q�^5���R������J4߻`ɒ7n|�d<�+Z��/]���𺋿�l_�t�\����׶F����X9a�-2p!��Z~�T�
�l�;�7�Ie?щ��$�hdO�DG<�2�B�>�;e�[����}Xf 	2�o�D��t
�xA׉����g^����a�Z��>�������g�ND��K2�F�$�>���,�@��r-�z��Ȃtbjj��C���Y��04K�~�F�����e;���!�^�if���a��E�]A.PX��7#cBD^�P�����v����Z�RA��(�TZ�`>�F"�Mf(����9��y3|	J�����ͅ������yG�kОi��P�x�@�	a	����е)T�3�Y	�ꐽL�òl��MMF%x��r<�.�|V�ύ�h
C4Gj��C���
��[���a͚�Zhz����h�����X���ʲ(�.�	G�e��|�4�\Gȗ
I�g��[}�"��A�%�� t�Qf=�H @��E�6��h�-m��ni�3�Q�SZ�R�i��3>��o&�y_7����	�M�6�P.�M�I^�GDDDqF*k�h<�#�� 2VP���ą�g��갋��C�$�/�=:O5����,rɛ4yldr�TT� ��o�h��L
�{ބ�7kPvy�ا>�~�i��8F?-q~Y��D@P#��.�f� q˳-0��0��t�{���>�����=�9�l��k28����	�i��"T�7�K!x�Xc���E��ẤP�0��i�2y2�!��R�����g�g?�#3�rdJڣ�#A�}�}��O��q���0yݘ�ޱ�F��;��M@��Dq����=�P�xLyv�`ww��ji�����ڞ_� 5 MX	VG�<IE�S,�.ʙ1<wN�k��z5���`�D��D�X�91�2����+�K��7>1���W_�R{�����h���jp������bD����a"ArL��Y5Ì�N,�j�bܦ��\�˲�����3n4�b�LC�d�v�,cCG���4��8��f �����1W,@�\FeY�V�<�<�b���ǎ���a�ƍU��9+!�|��R<!�̪wYH�~ӽ��?�������Oe���}2+ q�p"�z8�:��.Jiִ�qX��s@qZ�pE�'^�\���fhM��֏��i?�m7��l�Y��c���o�x�!H��A]3�9Q⤆�QTb]�K,����,.W��˾�gϼ�]>�����&��� 0���1\{�z���x��Hp��:�P�e���G<%�o��m^I��,b�dk%�={����?o���R	�ZR���KЍI��;`�ETe�Qt��ĴXx-�\�_��k%4�p�^��ߧ��|��ɉ�ķe����v�ܫۖLWӨ�1��グ��	(86pA����ʒiQ��E��������t!{C�\�����c���	�TF�t!J�T���j�񞢶i�ٽcץ��&n�f���8�� (F-���X\��;�|��ߧ'�h3E�~}���R�Vo��u�B̵Z-#����������R�3!A�$L���g���p���fs,ȱL�V)����\�h�_��bD�U�G6=�;��z�s�A�u����A�E��3��P� �' 8�Z Y��pY����z!ZWp�ʜ�\?�~w�.��Ƚ"vCĒȲ�eT�:�j��i��pǧ~��l�wN�:�=��q�g!_���ų��5���7�t ��٫�� �i���Q�
h���8�/_�}�����o�,�Bs�Z��{@,�/H�T��浆n�GU�jY��9�IUU_����X�.O������k}/H��:v�"-]�5�����c�=�u����*�\�֣�(����_����K.a!��>
^�Y1,�͗��Uf�Ŗ� �߿��X,ފrd}�R{�0�;}��Ŝ9̣��2�;U��&�) `0�sz,@w��A��(zϋD�B&�y5�i�*�R�������A���O.0�_f�Y'����MNM^�c�+;P���O�	p�$Y�F#e���x�%��"%�\�.�%��3��=����.�5_T�"n�R$�J�6#��PP#"p-^�i�5B���QI��Xy_���5�|Œ�?^�P�p����s�R~!��6Y�x�y�,��̈́�ȏ���f
^fﻬ������)	Vb��]�c>��ۨ�&����=��"��f�������,)�\�j���P��_��s O����&�YO�k���_����=������|m�E�$Ƀ�����2ǎT��,p�$����E����o�-�ȱ��\2�r�����O��� �_;~<�V*�����u=�k��>�>����U���Y5�]ύ���)\9�����R�nZ��?��'p�.F��B�/�upm�"c<ǽ����S��CCs?��e���+��`�!W_�>}�g�Y$� �}%�1�xK�b�~�p?A��PHI�h���['�Aމcǎѱ|kkkz"�*����.�{{�<Z[_�:�J%�h|��r��-=��=��/1"3|J�2ꆛJ��}�}�VK��F�އF�Й� �*�ȳ����d]X�Q��U�Q��,C�|Ƕ7�^�z�4��2������qc�q38���#8�c`+�km��E�'A3�Hy�&_��jZ��-㼘OO!�m!8�C�������̒�ǣ,.���5٦�IJ��\������ի���׿��{tw�U�/�B��L&}YowGG{��{��/̈]���:?��!65�a�\�|?��=�gU������}��?FDD�O
�8v�^���zf?���,Y��%HԄ���t��L1�d6\�
��8����1��?�;�}�ݐ�W��7�A����A���
ʹi��
��܅iVґ(�)/"�r\$�Yt�����T��M��={��x"� ����&!�����9�®7��'�ٸX���o?�y[9���u�w���6`��g&��������r���P�.�c�9��{V�E�v���W/�N���57\��-�/,9|��*~��?s��p��K!��Ҡ(��~
;�{!Lt�3���ku�hX���@y9�7���+��	��k_}����|)ߊ�]=S����r��y�aHf�J=��I�Ǹ�[���mo�NL��Z��.Cl(��0-��`�m8C�5?ŭWc�q�/d��NƇ�{�kdd��W��}����@��GMp ��#�EA�㦱Ia�c�����}�(gxhF�W����x������!(qCsZ݃$Z�Ĉ��-��P�$�X��Ss:2mK$!�ja}֫�)Ъ5r�;�z�Йi۵p���k@�`��U�֮��7wm�V���]���])�f��Lv0��t	�2U1P�3�, ��ޗ�-�D�ENd=L�p}�E�W6	$��$��ܰ�X؈	������B� ���Ie�ĔI�I�Z����h�8�ppK��̌,��o톧�����}N櫐=x�mA,��b� �Q��W���`}�<	��= ��@���b��Y���Ǟ|��.Y��E���?��z�%�8�N�Ēf&GF�]G'&��xc���Uj��[���}?iM.[m=�yO���w��� ��\��6�-�����^��T)˻��:�fO����]��	#GJ�B}s�pH�{���q3dal���dT�Rc�I��`H�jl丌O��Goo7��g��!@E�7t�3����聣�����MEʸ�M��a����������G��9aYE��(WJU���עJ<]���:5����^5*�;����1H[{�_I����i��H$�<8����]�w���+�4*��y4�P�M\��7����F�[�ψ߅�=�1�u�a�"�R還�:"�-�~>�_IA��@)._C�O%�Z�����b�D�khuƦ t��%+W�~�u�}�]3���l�|�����}�ͷ>:��1P(�Rm�(c.Ԩͫ���'� ͑�8s[B�<Ga��V�uu�Dg⧡s��f���T��.Da���O ��_�������:��|$�H��]3*�ݭ���� ��
�d���/Y��'G��4�Y�	��A\p!��Y84���Q|&iX�hȊ �� S�@N��@M�Rdلn>�����w�Ge~4W�1����	��t��0�hgM3���X�TU4�*����k�۲�l�����G񞧚 ��3ɜ=٬y8�Ec�$(<o�'���'�Z�
�j��yG_o_������L� VI�@�\f���jf#�O���IAG~����L�Ń�Ld���=m�������]ϣ��E��[t�ȑ�xn'�Jh�T��НR�Y��\��k�0����a�C����.�9.������s?rtxu4%�o�~!���t�9"�q?�A��P�Tɋ�])�oz�7^����xϣ	p�����J��v���Z�_�,�Y�5TȼQ�����u���m���Z~�x��!��M4�~y��Vhҩs� ����Ɉc�uI��\���=�M�6�''k+�����5�"u	�'Y�ɋEݯ�&��
�x"�<F��BC+mr,��84J��� F�L.T�f	�h��4��O�HB��l��ℰ-�O"��\W�B��m�T+�W/[٩l6������X}�e(U-dq�S"��\�K��-W��,��Ǟ�����7m �^����Pr8Zkh]ť/����r��S��WOW��$���B���`���jB,��J�>m/ѤPѬ�Y7������^���a�����_h�7��*~7���RɈ��׆˯�ߵ�(^!���2�#�?�P���H�3W>[b#�p�)��P�\� 0K���CL٪"j���Z-�ѵ��Q2��2 ,r�ɜ,	�"���D
��^uⱘ9aOS��)�P�O�����Qh�d�k�Cp�[-bn��м��}�r�W''&wi�J���V�YȐx�zZ3�l��R���Ճ�L2EB�ǲ#�V��}�ccc'zzz��6�q4��?\9�h5M��"�k~��: L
�6L��F܎$�t<�R(�/�DU*����R�h�9�X|��.	�ꎰ,d;UMGE\f�ױM���wv�m��|����Ad�&���l�R��V-�$�3���>.��BK"
ab���}ܝ��0��Ha��mk}�� �gʵx?��U4��,�Z�=�6ͳy�IOδ����7���tn*��d�
Gd�Q�W�f�S�VX�r%._'&s���xLO�x4��`�ܫ��A�����y�p��ص������5��u�U���/����H��j<G�X�%��T�(�u�3J�~�en�XA�B�ZCA�6�P��MZ㜖�j&���>u~�p���{���9��xu���	3\�����q�*cN�BC�q��ߒ����Ѡ�
�U�o��=�Lf�����lm�ry������T,��b9��4L"��R)o||����W�?�����DItf�/f���`	����~%t��kG��?J9��`�F�[�~k,�nyV��+p^q���{@@�-t��q��v�Q���X�5���T�	^ʓ��o�e��qh��4���."��ӯ1�h�$as�%�jn�.�<G����R+#\��tRk�W#_*�j�ì�g؈�ⓩx��Q)Y)�fH��+���f�y�w��]Uu��ؿ�r����Y�z�����W�-?eKgU�u��2-�DP#3աaX��K@��Zk#x`�ܯ/�8�Ne�ތ�/���% ��>���6@�S���X�5F�X�@k2Z0[��٩	hoo����C��K���	�"�p��$��;Q)�����S���.�/�����*<��S�)�6w��+a��!X��_���pߣO����;�:$P���;t��e -�p�gn�����_���HT�DT@0O�1_�5�.�W�=5��Z��X���{@r������M���t;��U�7-�\���Ћ�����t���	T�5
j�
����ַ�������>���n�K�HШK)�����G� ^I��z�^�G����֬��K��1�(�=3�YA�-�d�$j�,��� �Ȟ�(�h�]������˽��^�T˝�d2](�8����l�QCS��X,2���.P��b֥۶�vj��vtp��7}4��?<܀\������Zᙺ`�����fՒK��|n�FF()�%҈z�8Q����sjmͰ�9u�鬦���sH&bl�4�z]gT��
D�Gd�Ȳ%�G��Ē��w�Ks���o��}��k7?6ܡW+����q�L��B���9=�nia�!4�c�5�B$D]�h�9V7�@�g�`���˒�B
��mI��,����6���f���� B��� A�!�� vF���N��ɓ��S$�B� 2^{�[!=w9l�sߺ꜈ ��T��Cù�������!?��x�@^A�o�a�ͲeK`��^H�g�x�-P�Y���$
�hV� ;��k_���L���'_�����`��S�H�B��,�A�Eϊ:��ӓ-1>���������/{�����q��A�¤���ZPQ�R��ə�X�TV!h��2G��~{�1�쳔��y�f�������F�g�h 1��LO1��9������y�^Z�zu�a�b1�5�3_&����l��#A�����e��X�I�j��t��yjj�#�h4Q�u�����d�0��A�@�hP.�Y����䡦���SW�>�:�tn�ټ���p�X��zn�Cu�aROX��yv�]�<�>x g� �s��R�@�����H1=ڐT�Dɑ>���DsL Ҧ�B�D��6V�Zw]�.���h��� 6н��+zޡ����8p�dv�S���+/]W_��#�pT�BGK���EOD0�+��H��@�� ,o��L(����#Qj" t,�Jxܬ<��6����=��F�k،!Q�b��ʺ
"Χ-��T{t�w�����7���3���h� >�2��yp4���-�;��8�~k;ز>�߂�y����_���NZ���'Ylv@Ea\�������w��!�̃SA��zh��|�o�衝pj�N�3g�1F��=ᛛ6�ީ		V���X��X���`�9�j��w"{���R۝��4zj
����+8U�9C�L�W��n� 4rdVj���ݻ�g��0�ر�g-D0����!�v�&'���[�b��`��YM�f��L��ቋ�ㅾ�~�_��"�
o������9���g�B����c�.8b��6�E�v�T��ַ�c���c����2m��Rmʕ"Bk���m��K��K^�e������U����޷f��� 
�f���Mp�/�˞��j��D�:�Q�.1� �A��;32�� �NF�+R�VNh���?ψ�2Hs&w:�3F�P�<�����]R�xhkka���Ҕ�W����(��-7���}
Z�޷�����_�V奛ͺ����|�X�-_	m��K�"$SQ���M~j��z�k�h�P��A83�d�vA�)�N@��Y����;ҝ=O��C 4B	Lԗ.Q8��I(Q��$%v�ӌx&k��y-p�����ex��0YwQ/'��w(HFDa� T���ptI��O���N(������]&@��x�g`ǖ�೟��(L�K0���]�����`,;	C]m𕍷��m[�Ň7���X�-���0L����ɏß���w���((	-@����xA��x{���������=w���DӃ��cY�Q��u�
�aw���a� ����B�ྲe��ԓ�p�#�B4�ۛK���Q�����O�Sс�~�:�2�X,����1R$"��-��Z��T�SkI�P5	C$A���"�b�X�2�23���LAP?a�k$%2&�Yc�O6:����t2�j�R�VW�����	"��0`�
A���L�1�7��U@�L���j��##��Ǝm�Ӟ��xW�	���=R�D>o�+
QƁC~X��u#��!�ۋ�$n0��C�\�W�Ǉ�z�N��Y�u[��zM�c� 	�[,y���<D�oy��R�#q��W _(�nT@�,I��+/;���}���>�������mG��^4^u���ŋ/#?���+��`��(�x�����e���gO�!*ys���P���k�	\�\��N� ��?@pʳ�6�A������ɥ�i�*���Щ=^c��IH�3��@�t��g@`�.��S9��ӯB��QZ�ʪA�y�N����V��Go�m���T��8��,Z�.�{w�{�d	�[_ۆ�����?{lݻ��Sp���p�՗���^���R���=
�>�4pr�wu�5:���J�5:'�%0��M`�a��t��(�r_Wߢ��J�{�G���l&)~x傔��Q��j��j�s�g�h��.��kٶ,�4���<U~�c�a�Sm�(���Z��c��~�Z�sw}>���'ɪ�jtX(<&7��G���?)�z�yGy\�e��єk�jĄS����y�J�"��A:��r����=�#UE�)�`�5/�H2�,��5K�{"�3P�tB*��m���َ9�&ג��p�v�X��b���mo�^e�E--�x^����~N�����}`Ǌ�;��@�	�	��hYQ2��h),�NbAS�TaS� ��sD�4'�����^Ψ(W�D�jZL�S����
�ȏ\�d	�d=P#�� e�u���lC�u�������ƍ�kb�?����#W�~��O���S��(t�G�a݂x}�v��",_:?ȈF-L$�y=��q��+U�!��<�\����/e�8։6�Y]����߳�3çF6��A腾�H,&
���D�z=qZT_O���<Ԕ�1<=�t!� B`߃mNC*����0,EK����`��.hO��e�R�җ� >�8�:	V�Y�t�f��O~�� $;;�T� _�/���#���O���9�񫮂C;�Bu�4|�w�O?�(ģ*�?|~�OBw&G�O�箻>�����}�9|�@+���jZ�q����Q���K�85����ѣ
|~��M�������9Z�C�V�ɲ�%�.�-i�3>�FݬT��S���-[�?;�����W��)��b�T2;{��k��ƻr�՝CCCh�{\�T|ϛ�
�	]J�Fy��b�$�Bǖ��>�'_I'���h����O���0����h�cM�XY1/�X���
�"܇.+�~Ϛ;#����ֽ��{"�μ^�i�TYY�s(a����=�� @�3����Z�V@�dV2I��Z}ᑃ�W%�A�����MNVuI˨<mO������d�,�D�!뀍L�3U�>�r�x<�!hq��:+3"�1��{4M�������P<��X)�_���¶��=��{���:�߷x�	��o�%Y���N$�=�a��&]�A�E�����_@:y3�Zo������A
7uը07'��M�qlL����T��r��g�=��*�t��:�r��9K$!@B����ܹs����3�޷�]��{g<�1&'��A �(����V�su�t�T:o￪���6s��մ����	���������S�6Q8X�|����	�~�������1�P��(,�d�}T2�6;�{���#�4���zz�6{\տ��k��?N�Ӝ`%=�i\a'�R����T�uk�ŉ�=��Eh.;b���pι�0�����ػw֮^��+������~_��|p��:�S���k�~�!���ek�Ɯ�Ȅ�8�~]|�͙#�F}��mx3�,���|{��Jn��6)O<���A�� R^2��n�f��~���&n�_��π�{�i-��<�[,gS�]�b�YK�B1��g:�v�UMun>gݚA��~�g�stww��~���NS/��R7����x��/����&�I��5�����K��P,�F�rFC�K;;;�E&"%I�y��W�-M���mW�U��S[�+�Gd���W�
��C���\gʩ�����<R��x�>8��lw.x�e~�|�(�
�hh���C����'�����a��jK�|� 焣i<����]!ʶU�����h�#���=Ε�1�X�N�F��
Z������z^�F./�AYo!���і�`�ژ×0���~�p��r�|"vM_8q�X�Pc�й�xφmR��|��x�9�:s��[R1cz\�.$h5�t�̙%A��S����$D%�����^�� @e�:>��*���I�U5a'��y��E$��5����|t��~,�3���ك�E+�x�\t�E!�\0	��(�(f�^�����`_'V.^HF��L��ph��y�^rb� �B�Q>r�d���z�����6�����BV]�%�t5b�qA�[��J�p�U�a��Y�$""�{��gq�W��熕���_�VP�v�ێ���������ڮ�HE���@�˧�맷n�<q�y����}7���"ſ�`gF�☜�c��w�\&��\�X�0ȓc>�v�54�K�����fO;���S�͘>ód���&��#�x�JlTV 첽`�P��q+�B ���8��J��q�h�P-;ٖ�"����x��-Ƨ �E��Y]g�S2x�0�����5�'�����A�׷+c�����f�6L&��@UtA�g�xV`E *ك�%tSt:�y���;s�E�(�VL�/0&�Ae�r޼f��x6�*%�3��Լ�����AWL���{K�M% �"�0k����1� ����<T�.�׷�}B>��XIV$�����]��`d�I
�d3�)P�1����?����y�߰����u�]�1�'.)K�6�?]�P*p!�K�*�N�'��76ឫ.%@�����6ȌY��g�|ˌ2,.$(��轶$[���Y���D�GTS���2�NE��#sE��x�0<�����B�v�#�+���Ɓvtuu�q�b\��L|��C�=�3�(��}�����������F/��Dc1̜1��b	E�Ӛ�t�B��CJs��5��18����W�@45�ǟ݈�����}^��"#����k1�m&2�r�~��C,EGK�|���M�ށ�������ljD`�:\��m��Ϟ���(���i�t��CÉ�������~哓]_�Q�ⰀS,�v�wO��:ٯ�m��;JYdu�O�N��d2�-^��U����t��W�>��s�żh�c�q�d�F@���pNib�A2��ЁZ��&�f2B!��S����Z�3Y��&8jg�Q8T��L�Х��,WE�����"˿?K�G�.Ӱ+����cz"�Q���/�646N�XV)/�k���%[EhM�Q��t����`�t�>L�/4&�Ae�ա��iI��	%K%o��Z���e��ʶG�:K�je�f��`����H���!�������{���3)2E�Xb_��d�5��rk_yϰ|�h_�/:w���jjG[g����)���7�Z��M�R����5�+����9��-��ņ�T��b<DS�,�Ǝ��׷�뗬�Ss���8d���ӧA�3��3B�]�t�_�Z�9q�i/�0p�*���̀e�~f�V�� <�UQ؄lA0_�z�`:r�4�uj�w���>���k@�Ņ#��D�?m��'��E�G��ޜ�x繈(�~豧�t�"�`�b�J�߽��>�͝	�X��y6V_z��8�g_}y����FFW�L�a"�+�7��+p��wb��n�锉�X����\�"@��[?�Y#��kC
�|  ��IDAT��Ȟ��8t 7^}	=��ɴ��֮��K���9�L� c*��c/X���G�o�5����O��Ψ,E�(=�J�fD�ᵴ�O�3K4Ukt�=n�Į�F�#5
�3ӬS�#:�*"5�:��b��݂������!��XDI��6�׊`"e���V�'S�����
~�1�S�T��Z�d<�9�D��?�B�kt]?�Ρ�T�r����i&Q��*]Xh��$c�̻#{ƾ=�f���'�ؘ̾����+I���s^t�e!�����Y��8-Ǽ�e���1��H��-��s�R��3�L���� Y�3r�
^��.{�P�"o�$�I���������j|�?Kh��F�h��d��;��15m�cJ�c"Ev��Cs!�6#�v;2f���tvOF�al���U�-��j���9F�[���UD�E:���\�D�,��B
�%�۠��j�S§ �' �Ӡ�T�:��_�QDUH��Xf[���:Wqw�P,��dt���)2��X��(fOi�Q2°��HDG��{��;n�s�>�=ݝ�	��s���>|�O_�fG<»�o�p2�[�Oxc�lݽ9I��"�l��.��u��Fʲ��#���G�(X��~�u;�;�\��Z��/~���W`��b���ԩ�him���3��6O<�"do3��6b��(���hl��p,�(���w�'����������W�'�WhT\)9��	gb�T�F6������
�r �u;F:�b�H�I��fV�d6Czmdl�=�8>ܾ��9��v��V(��:��T0�Z6+�߹���Yh�\�[:��ߧڇO
U����O��h5���� ��o�&�W�|ŚD2)�D�A^�Css��l�x�$Sq��a�;�۬�dI�:�v,�D�01����$8�d�����R��T�{�YX"�/H������ޗqJ��!��d�`%�b�`�޽�T,V�Ig]�"���*�)�9	�&Z �5�4a4���o�(�5%�s���<,i$���x6�c��9K��>��K%Y'��B:���p�
fQ�D�/{5� y/]��8�#��6�v��g��mPM�>8�t��<�W�@N��#A�6)�f����	�L��� �v�B�;�?�x2.�k����v�"�5H�'<���عg/����>|+�,BWG/��Bc�G���e�t��0��o�N��2��淰��7�|�|�(�Ʈ�� c�A<���	�p���g������$�I����v;]��)�5�K�#�-�ǿzW�9�~��x�_~��� g>�]t.��"��9��~^��D́�c��%0�]Ggo?Zf��u`���8�x?��r��Z���뼋������/�������5:	�Z�3��P����r��)p��.�LpVn��;���]?��fWO��9{�렣�?������;�����f��.�G>W�e;[�v���:�m�d~;3�@���zR��Ԛ���@��~���t�'���|�x0��mG�����,@�;��r6���t-%#��L��`0x^���/b|�1	>��9�IR�&���<�XUw�ީ섍tV��^hQ��༬��T����b��d�-k����������N%G螅�L�7R�jdEm~�j0�B��jcjhC#�?�������7������vݕ�7.����
�J�n�H_jNER
�Q���x�5A6�M�*����u�Xb������
�"N�I�q�ܐ�9ZS�?��F�έ�����)�t7�<�gds"[�U�l��o��oOT�VհU���, EӸh��؊��l���I�8��!k�a��q�iKQ�%)�rB��t^YԶ��N�sj:]��w�}\����=�{�E�� 7��-�C���szq�w���#����n�	�dͼ�W4�5��l�K� 9:����mƾ�^�;���>� >��@sS,],���2�Yh�� M��t��va����'~��p�M����h�ނ_>�N�̩MR�C�ǳɅGz����g_���=7?m��'�Wgp덗��(6���E�V%{�`�k��a��s@ÿs;\�߯�}z�F1_Y� �Ɋ߿���"]��kE=9���Қc �_��T���]�-[������k�:*]%�05���Wv��ƆwG���n�'W�� �息�S�OΤ�����s�.r`��)gt�M���չ��)2Y��9�$8�6~���L[/���� ԭL�R�&��9`�q[�2�n#��f&�
�O8�rg�Q��QU�Z 6�,sŲ�+����92`@�/�3��=:�AfW��j:�vfX������"�Y�54zOVq,�+�ܕ��$$���&A����S�&Wu�u����䈹��C��G��-�\��gLE(��[��Pg����A��g2pV�%�ӥ.��d
�@�0Uy��^��w���V�*���p�L��΋P���h��G�;���1m6'"hv���� Ok�Y!���'�dut�9͍�!B��{�n����d���ñ� j��@�l��|���{u�(qB.�S �Ʀ&���G\t�h�Mk�jב- J����-X�%�ફ��{�ih\o��<��������1<0��&��+�&`�a�p�Wc��7 P���+���`����3	f�[��l���?8w����~��s���y���F09�*�ۘ�MN���JK"�=A�n�;	8[����؆��ó�>�]���/&�2�f.�s��Dss3֜�Z8}^'l�]��� ]U'��m���#��`S~���
�鋂{[!0� 8���?J��{?��=����'o2@୅֖&!=��\We�,Lt:ʚ2Ţ�nh������9����$88e�l^�~,�-�)�f��z�"J����mF�T�2l�-cf}��ц��Ǘ^��(E�3�K:\.3����Y�X���m�H��-r�f6_f��-rٺ���x"���=_�������f�eãw��YO�%��{�#��@�@�6Y2Z*E��S]/:�b.��ӹ4ܞzx�>���W߅��p����8����jk
\=�%���(BW(r!E���H9���l9�ʭ��R�01�e�"9�ё�����Dϱ��Q�&�Zf�`g/����k�#���@�[���c��.289��j�(F�B���8J�-X�Y3�'�>��H�7o�J���[��7�yG&&p�u7�ŏ>�K[wc޼e����CEptSf��U�G<a���(j*&���V�"����C(���m���}V�Vǁ݈1%�F*��4���PdL��|%$���_ހ�N[��k�,��n�h8����Χ��ĕ��C�e��]����wg�����'/jt�cr��2dBP{R��J����%��[��+��� ��\6o%����}��w�}W:v�G�9�
��<��XC<\~����k˚2Ry�XiKZ`/U�Q�|JF��-�S��N�m�޹�l�GT�<��c���vw<_��UG�(H\�%p0mj\NdJ��MCdQYΜ�rrl#�
M,no?ě���s�Ipp���BN�)�t>cؤB�ZDS^(
��m�lB������BYa��@08�
gX�g�}��lz&�����V������|�B�C��s������Q<y+�L�!��B��� ��V�����}e�`9U�	Q� A�O]U�������r���2��.(�E��kQ&���( WB]�4��x��]B�`�6�t-�Z� )�(F4��6���&:8�cV�4�}���Y����#��u̰���->���N�O77R�><���cp4� ����}�49eࢨJr�`�eS��!r��e��l�Tg�q6��c����3�E斛�<���w�����.�dЎ�N��m!cӑ�j��fф���y�1����]�(d,�	�D�|�Sq�<n�Ƈ!:�<MPwo��1��n��2,�ފ7^}	�pC����X��Bq~�Я���Xa>4��kW����~�ܵu>7:���T:�y�a,xW�9�xұ���y�v��p��G,k�B`���+0r9�Ù�6.,�+��V�rE� V���oFf�H�]]]�###�55uw6����C��,���s�=��ʫ��`RYϠZR�6��w�U��AU��Ԃ�j&�*Y�*V<U�d����VH����\R�j��9�t���D�3��)��:�v]l/����A�k����
����c}��cmmҿ�8���c�2�~^��p��KeM�d���t�fX��U����r�{��P�<��D&2_�}�,Ɩ�?t��7-E��f��Ҷ����I��E뼗�+���3�tA�����cMG7���\DH#�}$_�V[W�!iP.���rT�dY����?Op�j�3oA��N�h���ҝn�X�F�����#Y�G��Ǵ	/��B�7��S����Ln�I2I#+�@$Ԫ�dr�l,���92�Pq�0GB1���,[��_�l���㬅�?֍D6�~���uS�3Ǽ0tf2�|�qQxǝ_GK�BD"�tK��p%zF���ko��mx�9̜?W�tŒ�X�l��+�1l-5�8w�B\~�9�esؾ�%��M���pf�qW9��"&8�`"����wc������9{��V~��#�9ډko��x�mz~����[o���ǅ��|��#�_q:���c�118��Ӧ�A�m�� n�t-�@��^����wDC�����?EO5���W4�ә�s�$5*�iܐ��VX�Z���N�Y.��م8�������d��Z�b�ķȩ��b1�y<���3N�m�ގ�˗���DS>���-31C,3KyT����)]�f���z��GHX�~+)r������`ᑅf���N��u@	+s�4�&�g
��\n8�.�%,+ӖmgwUY��׏��.����'�����$8����v=T,����������j��0�?����X�3r�'�"��)�����L���WDO��9ƫh�y��)��,���	�����H�f�7tRe폍�aW{�u,��6o�`,��)�o�H]J�I����P��x�H����&��yk�	JJ��Iӿ�}҈$᠈�Ȳ��ϔ��@�ظm7�\�\��i3I1�n�C���t}��cӦM��[0�hjj�9�� �k2��}��5�`CC��:���^5`���.Y��u">DEL-�Ĺ0���,UӀ���I�/8:8��{7�*�x<��d��$\X�x1�[wa_G/�5u�� �X^<ܵ>�"���<��(�;�"�񵫱�����1:<���a��� G�05ԏ���$�홧���}�'pt����ݷ���pӵWa���?1��n�:"�w�v�˼<G鹸�j�ڦ���r
g������
��7�xN_-�.9R2��.<�@��o�`������?�͆⾤�a�G�L��G�by�i:_��ݙdr�����f�R(�u�h��v�l�~��;L��<��3��=s�x����hL]�l9���Z�'0̒м]ʼ�UY&���*���8���DQ����座�IY{��|
�:��e�U�H�R�Z�������O(J�C�/1`�V__/j�xm'�	Q{�[��MbSʤLd=�hd�p�T:��I΃?>&���GAW	J��eX�\���i�r �T�CY�'%#WEפ\Zv�c��p�`�2Ol�F�b0�B���G��łh�̙e�ϋ��Ud3�1M�*�9�N$���7�oW$�By��H�s���ƃ��k`v3)�jȓ�a=V�؊%:;xKAtP,��QG o0��H3;�`D��\d��Xi�_?v��b��b�h��Ӛ��	�! �%��юx��'1|b�"���nr�hs��"s��I|������m��<��V445c��%p9�).��py*���u #[Hҳ�4ܭ�06Ѕ|2�#�<���`ђE��e���~C�j�-�e�"	�A�g��|��)P�!��%�ľ�b��hin���q��`㫯�{psH��>�v�jd���}�����]((&V]r	^b�]���õ_���8���&�kkk"o%r&�D:W��.�
�dy#����ރ��1Q � @��Q�Ι��֞)�sǞC�K��������Q��ar�ݴ��|w�L��%n�[r���R4"F`48zf&�9GS���_~���ֆ�sg�*5=e*b�(2yY,@'�T�����X�����{N�W7��]Q�O A����ҍ9]�2��?��6�Q�X��t�f��0�*��x,)���:��*�%�������-�6��s���l���69����^l{w��)���E��4�*�ee�%�Η��)Rf���6M��;)_,��D:�Iƾp�����K]���|�ǡ�e����D��K��Ȧ�`�E�����cb���~:��$�K�d2][JE���[sZ�U:R2���L�1_P(�6�V��탤��(�j�����Q�Ί��cYI�Y5��%��d�����E.^r��T�p�z�-�r�eP<5�(2oj���x���)����Ͻ�;o�躡�\.�C�8�r9����T�.���w��G$/c9T���9�ba�yHO���z�Ysf��	�ma	#�4j�g G�*�ڵ��yJ �CEʲ�7^���lE��A���+��qa"Dm���j�����Ĵ:/� �7���"G��a�N��j�x(�w�|816��=CR�y��iz��{D�Ú+��@w/.��zd#!�w��!F��128D��O ֎��n��L�7�=�+�[���Q�܆�X
s������1}J=���r������u�\�D2�����`�^�;��zf�$}� xr�i��7�8�N�Sr4Y?���#[u;!���Ӧ�͟�P+gC˝V��[���5L�Ľ~lO
�by	��H���]�vቧ�!�\{�H�E���w{�����R��#�Vt1G1Nvbb��֯��nw����tfi\�)����Z�/ծ$����BvG�`��/r,W��G"^L��?:&��o�ۑ*)V��J��W�	�Hծ�D���	Oh4����4�v�NNM��vۂ�t ��p���,��x<R�L;����M�;��U�'�s�q�)t���&R�ܩ���i2e56�ǋt6#�t��oͤcu����K�󬺃��ئ�xd��[;�cK' B��d���JBV����ӫ�h)�ŧ�d�ʭ��%E�4òI�t���Y$���q]*d���ݸA�a���x�}x��0J��Ԛ�	�v����p�_G���h���d0�0IC����G2k�s�8v��p\B��cM�^�@������̙���I�%�yZ+�r�-����#�-�Y;�c'��;�p�k0k�l��G^�+[w"h9�nlA��`$#)��udr�H��O�s��3�L���"LN۠�{��M��y1o�6���hA,��p&�mo���ο�\B2Y+� ֑�Q�4��7�E~x/����^�hm¾�;q��A����X$*�V��&�ݬ�h�?����0�e
Κ���}p�68t��}86D�$����]z	��`��@{�7w�3Q��,���� �+9�g���o�lSnVUm���5����My��: A�.i�Y���|���k���ݷ�|G ��C�X�d9�<t�M��)�XKB�� Re��d� ���Dحl��V�zj����� ������pkCKw,���W�0%�q�P��P��O�\��`��k%8�.�S�~v�B��c���
��$����෇�mʒ�H7GP���Kr�̜&{��6g���XT�V.J����ټ7�Ԣ|o�4�G�CJ$�.U��~�W�"�l�L$�x�O�ĹH�@�1v̌�	Lp��C�F���H�ƍ��9�xq�{���sܯ[�C3����&���灷d�@�����]��I�D� ��=L�j�E���!�%�E��*�߳��E����0��ǒظ�Ch?E�v$"<��>6L2�
�����0u�\��,�����z��I����N$KEo��DH��6ŏ���H:*hX��J4ST.ۊX�d�(���
N��
�����Qa�J%i�^c+��AD^�"���`R�bolB�Hї�D:aP�X���1� ����p�ܩH��X������O
q&n�䭫��>�9�΀��c��>�v���0�����`�Gcˎ]�46(�p��/���7b<��Dv��&�OM@�?���]�nX�G7>�ںV\|͍��헐O�qƙg���APT��)u��sˌ8���ph��Zf��2_�{۞K�tt#�@�:�^X�_��@�MUum�jS]l�I��˵S
��
\n������y�q���ۋGϿ���ׇT�6��=�K�
+q6U�6ӱ�ul��L�"��iδ��2_$�*�
�@]�c]���v{+�}�TR|g���/�6��$�$Z�]�_��*Fʘ:0xb�(�:�I��?8&��o��Z=g��Q�2��^��U��꾙X@B��zEU,s�Z0̼gl4���З
��bY����툪y�<)#]�vT
ު���� ���ϓ���}�\�X7i<ͱ�sw,��W������yS�*ML�����כcm�,}��gYޚ�� ,h�@����f�*�PN3ʜ�Pʊ�=���Dw����E��a"��ӯ���W_��w�<�(l�x� g�d�	���z�@39��t�8��� c��tDv��M۱�x��w*6.Z���#x�p;�w߽�V4@(&�himD{o�.���/B��0N�;�=�Е�j�1�l�r,f�Ј�j���X~�5�X�v�c��{�btoE��\�۶mC6�A�@BA��Z�p�5wxx�v|��;��q��o�^D��hkkAM]-�{:�&ÿd�y��SO��+/E���k�>��ga��G���!8=�'���]G)��y�g�B8��'@�_s�e�,̘֊����bř���pѪ�Ec�#�zW��>f>�ʫ9�M��ܐ�N8dY�˄@LDV6I��� �����d�3��49\&>ڳg~�����#���?��Ұ;ݢ��M���iy�BpT���'?Wy* ��(j�e��/r1?�����?�����d�L%�ve�qZ{l�jj������#�I�}������N�,'�Pf09~��5�~�Ii�&TR��F&R���.���s:��
d�9'UѸ�9���`�;��S�?{8EG�P�u�2g�_�����9a�%Uy������RZ���"{#�F�&&�܋�������л��Fr�Xx���K�%�L�?�DV _��j*���hc�NQq+�$�2)�%!\�}�I%���Os���Pt K���������&�v�7��3O�E�L�(H�"U�c����/n����q���GS�J*n�����s�@�bJ��,�c��L������W^�F�.]ÅSVa$Ƃ�F�׿�|�?���z��S�S�R�4Ni���i�����Aъ�I��B<���̚ ��G�T�7�aժE�'�;}�,,�7Kp00\(A"��� �Ӹ�2g��E���O��o|?��N<���O��[gk3>>zSjk�����C�Xr�\~�Uxw�vD���`G���Ώ� �Q|s��&�3N[��{��e�����`󛯠��J�f.�����n�O�������U��9�k��vĲ^\$IL���(�z
�f6J��U�s
�sK�;E�!�I	P�#lW���B��oo¯~���Qw�]HQ��Bjn�rEJ�*�|*�aUG�T1&'�a��O�=�O5�3��0�pxt�b�u��Q[|�|mv�ܵ���.�����1�p�;�-�F[�T��]�L�����RhUŪ/T�m+��e�!���s_|�JV��6G8��/��19���f���x���2��m�� >G�<Α�ep�>�)Um�*TD��EHα��T�ɐb_$��?�ӝ���a�"��m'���q�jS�9y�7H�C�-C�1u��h�&HV����S� 
'�X	�((Dց A����Ru���`,�?����o�o~�<�$l�z:�M�(����1l�u
9B��Ӛ��8�7��C�mE���:6�N�_�l��A|p���n��
̛ۊ�Ӆ&�#}�������=��'���[��\����D�B�,"k��(ߢ���p��aG��L�7]��M��ֻG"<�dt s�N%g������	� u1J&�4�S�y)"Jgrt��x��q����W_��w�D>���"��`������K����/�����p���x(���)b~��!���n4zk���'�����^yg���f�����8���Q��>z��=�2�Z���u
B��p�ek%��G];;W��{/ͩ��+a�0�+M� |祐��v�RُL#1��pԸ���|���eJe���E!x��Є��<��Cؼ����`��	Վl��BV(����\�_� ��|s�@Qlsr��U�[)��9M���}��O��3�nhl��W�o�5G�����=S�Jb{�t�UpP���x=�N�Tj�����+����̚��qL����$�{��0��8#�jA[ d�r���:#G��[��UN�C�H��P҅/��q"�v��o`�fY�h4e�BiZT��햜.,f�'��`O�(��y�Nl�@���جP02e�ƍ� �>����7���?�s�ݕ���_Hg��y��3Hd��Y�P��Ȳ��bD^�2D��HN�Č}�H�r}��p#�R&Q��i�U�q��Af鸁Z?����Q�o�~��|���{��'^�N���l��Z�>p��вr&6����hB�" �t�d��~M����Ǘ5?|-:vw���~��:���q�	���⒋/�O7�
G�$sE��n���$Kt<�KAft�ǻ�b���;�ཷ_��sQX�﾿y#��D.�%Z=�/\�����C���p�=�F�p��Ӝ��sIS��ܣ�ƥ�܎�]�NHB�RI%5u�x��7����\�G�}	G�1}�LLm�xi�n��Z��i,Uý�x��'��2ܦ�ih�6�H{?>$R�M5^����n*�ǡn\�j%�ٔ���ѥ;�+�z���a�$�09�꣩�i�Ɠ�DQ)�LSn����e�LB1��<��'��t����dԞ�.Zz�hg��ۀ懙'`�1����ۇUYIʗi�+���Qne<�\[I�S�NY6��_8j������_�|5]ɴ�T�3n.@�-<��r:tA�$(�S���R*���+&��l&S?26�<1n��gL���~�?EX7��e�d�m�yq�M���[0h��쁙/�Jm�*їK���q����V�l^��8�9�((*-x���+���mB�P&`�șWs�z��tY���hJ���:�石d��?a����M&��<���U���`�	dZ��K�p����eҌ���.Q��E!��J������K����'�p�"�	%��Ko��ǽ��6|�a2�~d�Q��x�Eذ�#��Շ��9�>2l��(t�2�����d:=�z+�B��O�����_?���\�����-$�I�$�F���=��,fm��p���"|'�;[2�m��8�C%�9�D��ƃ�N�0<8����E����j��U�s�	��%tT��4������#xk�S������;xl�st�TD�1!��?8�'7����]oD�vX*sͧ�%0��"[ 4����͈Ҝ���}�z��q�����^44��Q��(91�i���>�}�\
9���ݷoI{���?y����h����$@�+�?��km Ϙ懹Baa�*NU$[�,ɎB._8�7����	r[��?\Bvmnkk����r��H,do昡��[\'�0��O�T>��A�l�L���rJU_8s�C�i��榏���9�YN����d�4�9�.A���@�4`�l�H�B�3246#+���1���c|�P�>����f	�� #Q�6�vF���h���^�I+�]"t��2��`0�I���=������lE�|H���{j�<$����ɼ���6��i���L��A���op4X�j�_�'U���ՙ�~o�K�,}���|�]��Z��ˬ�V�B.���Yl��a�"�'K�
O�	�$������%�26vo���GCx����w�����-<��o�1b8��u�⺫���x~�N8��(� �.�)��54"O�su��k@&���Q����U�B�@V# A�O�y&Jt=g<��+�����F�T.A���,'mSL��:���Nҥ168�|�@��=&�z{Σ�{���HY~�#�b��{��K0;*�
*V�d#�Q�
��,�D�BVܻth�^܈����{�߆{��!��,d��Hx�Բ\��K`�0EZ��r�K��g7oFJ��K�቟��=���w:�T�>k��fHF?ڼdq�2MNW��
v��>p�}������b�[�E����,eh.t&p\�B���bm.��'si�SՊ�u�fO6��iK�-=���]�px����+������+U�Ѻ��z�r֠Z�]�V8�$�b��MQS����l���`����0��]W�d2)E�>����WAI���m$]�=�̜K�aRm���Ip���0].���d8뱻��[6DU�̑�C+�h<9G^�,��^=*�K�L�S`:-NYh�늋�J��!;�b�ʋ��pVks�XМ�����2����9aMc �'+�����|�[���r�]�X��=�:*�����2�y�n�<�� 9<�)�V-������Wʘ�R�$�����-�FЊ"��NR��	`0�c�<�[o���v"�Q\p�Z<��s8�?�9{��K)/�6��g����|�\����E��d.��ƀ�TGF�X�(an��H}�fl>�m�D��D���5���T�HǸx�u���[�D1Ć�^A�Z�a�L,$G�{lP<A��͐���k �$�|����t\E �ݣ�iS�1�R�N��N(b/">6�c�j=>�q��x��{O�q�57��qcb<$x�5�7\l�33�ث@?�M
�G��MoĻ��E��7��x���g�d�bù�B4��� z��M�gs���f�b�r����t�ν��x{W{!�4�N�zu�$%19���wP��S�m�r�R���4�$�g�"d�Zi�M��{J܌Q�m�F&�w�*�j�E�ᦈ���Xd8P�d�uZU`�[��bC.��{���������/mxpCp�Gۏ+�2�&�ޢ̊LnA(�V��Hg�|�(�̔l	�hmݝ]�_6����$8����7�v�1EO�LӬ)V*|K"�UD�/�cX2A΀#j��#A���Bc��Q���m�ly�DF@��H�ܭ�	ǹ"�TىZ�U��Piqd@P�t^�x8-X��x,� 64��ϒ�����K��֖}��ɘtaM]s}4��rd"-N������V�@�ʵ�>�r9�h��Z�>��l�~A�4���8��	lx�E|�֛�p�\<��386<��C�>#S�`7��8@I�[��̏��:�l&��*�2&����-<�y;�\4�(�@�mF$o��:�M��&Ph�s��ȩ[y̨�źų0���������������C���64���%s砉���c��-/SF���l*��+@�ݮ�{ĵ�|^t�t!��9]�k&����qإ�Uk�ݻn���~���4�iA�%vHt�l�횮���^�c$Eƴ���}/����=����"~�^}a�Z�=�X�p:�tb���u�0����k0�����A�p�eMe]G::���=dӟxG�Z��L� |UFe��2�E�C�/���K˽^����;��R��%h�U@���=E��k8�Ϡ�^-J,����(�����k����<�����?���e�In�\�m!��2���98�5��4L�Ś�G�fѯ�b���3�$8��A�|�WƊ�b�d��%<�D�pA�h�����@�(������J6O08�/ƾ�^�b1g�l��:��F�89�ExZEZ���r�@���٫r������2�z��L�9Q�e�#��7l�Y��/~�՗K��.����@y&E���	$d)f
��\��VEڵzP�u����Pv$I2
��89x�t��������ڌ=E}K+9C�"b��
b8��K�ɯh(dM��/��]*�ڄ�)Q'RrvYr��n�-�q�m�ٍ\,I�K7GL,���ջ�\��KW#>x͵���2�����6"<���wq�ʕ�in�ᯩ5\������_�/��e �E�#c���r`Ɯ9�D!C�K#��L��m�ᬋ/�w�y~�Uq]f>E_����$	�E}A��::��M^!�X$���sS�ePdk�)�7��{�p���X�h1"'F�T9�V�� +�0�; ���М^)��G��[�#<�UW'����3���=���vtΤ�bE�6��oQ1���U���=MdpL�XM��+�VS��F�P�M.w2ZI���s���O�M���7���Z�a�
gޤR���*~�Ȉڬ\>+��.��.�q���)�㺃�����������I�IJQ�d��3�s6��؏�IǼ�U�Z��^E�%ݡ��hlzhx��C��H[�f�IM�h���0b�·��R1\�T+���bS����1�|�X���?���a%��g��o�)�����囱�H�-���[��3��ܹ���Zќ/�܇�l&T�'��]  �
J�(��l�����!vd���S_7�� l��&+d�
F��k�%����9]/=�l:AQu�D�7��9��2�ȉ�\&���s�yF�]Q��+0Ƈ)��bzSb������Ai�߽�69��HW�� [�{��� �1���1�G���ƵN2^a:?S��+Mr�y��q��	M�9����9'�bs=-r{k$8��7��3��7�pv�{2��c&�As��
 �!�H�6��	
f��G���q�+0���G�7�X��xc�&t�oǺ�k�͗P�Ԉs�9Ǉ����Δ����002����B��b��17�+><�s�U��Ë�[_�As+vƪ���ƃ+Lè� #�5sR>[���P�%�[!:��Z�>	�9�bP.Z+ň�`YNx��?��G?�����*���i]��N��ϡ�u*�i�r��J��M>g3_��s�YC5��9&���uu�I]ՆL���$���'���I'��,(�b!�q�̤P.��6���%�ˆl�wtR����|�*C*��H��q/��4��W�[猁�[��rK�\�jиFB��y���ӳ�oo�_���w�����;��$��٥d���<�@ ��DN�T|ᬀL�I�%Q�(U��JCE鱌���3h�rTm�l0I�w��G�C��U�M`q'�Da#Oz�bCI���\4��daH�]���X,�چ)�*[�L&aw� ��幐a�E�H�R+�5�na+�x�I��tvw�7�<B������h�r�nnAgo��y���L*U�"Ƶ |�eeM�dL ݡAs���8���4z�{�l�b�h���)����
g���c�ۯ���_Ǣ��pt��d�]^�}^�A�{hjB�>�K ��BOE��e���ѻ�,Y���6�)\s�����!��í*P�H\3�G�����+�i�郏"C� g�s{�������P�f�챬7�HR��+;8�����=�߿)�L-�
�r���/&���.�q\�����Ŝ����6��6g�&i'���/Ď��h=���c.��+�XC��ɤtܝP坩h�`�<�ѨpՔ�%5cd���ar|��g46zS6��[L粲��y���g#�T���0ev.�tN�.9&EL>��C���@ 墟?7s`˗�S��*J/��roqY�H�LvD!��}6��N�fj^��"E�����p4:�D���$�4���i�A a���Y�|������t��P�D�A���d%\h���$��[�$�e-�o�ުV?��,s>�~�b���F��ȶX��PԂ l0�ɴh����\d��.��b8�:���q���ts��T?=g������%����Ȧ�ܡ �ٳp��4����/��Q(�m���,_�5W���#8���aw:�c�,6�I	�nQ,�AH%�P	��oe�X ������ٔ+���3faΌ����[,��9@��d/=�����kQ枠��š9]�R�*�bd2M (��]��B
C��hBl|� gb0y\����W��s`��U��{]c�Xuյ��U���h8�>M>���%˓��r���oH�	 �3	�ڃ�izɲ�{z���S �J��QU��U(뷈�n�u�>\�KAd�*��*u�K5r�����$K)_s͟��_����u�N�%l6)`���'E�$gy��MƩ
��.
9)g����F�A�dJ��1	~Ϙ:ujR��%+c(�/Qs���Ȼ�sJ�@Q���N"V�&+	���F�q��P��j+�����&�_I���EW:�Q�
�?�W�)z�"��bP�+F�E�c5d�"�)Gwq����� aÆ#�VAyk�Ǫ��gz��Q��2)�ru]��VEX��lVy���!� Qf9�r]�r�cy+�b�Lz&�T*]�x�E��.r��e�l*�"�ψ�Wl��v	��&��%��>̾h^{��e�=��:����v�q�'c20� H�A� (fR\QY+�SXYڵ]��]��~v�7��JT�I1' @"D��`r�=�s������4im-�E�氦0�N�����|'}�?�Uy��3�D��'/�Y_#r�H<	®5Aʦ�\���;����j�~�M<����<��˨��`��s/��۷o��m�D޽��v��)��ϧ��rF�.+���f��S�IF"��	�,�hBp���i��8l�s�<S�����	:��X�t6���
a�����i�Z�QE�+Ž۷��5�Hcs+�r���������+�q.�����^D(�A�����Z�����j�PH);���;�Lx��(-�f:Eێ\)��rѯ(�x$i���*l,�HV�Z�N(�Ȥ�n�p�e�Z���:�ua�ޠX�_�NV����RI9B6B�:Ym�|lp34Z5�/_��s��u\$�"
��yR���db>�a4��J
jy�?i�z�mhs~K���^d��<PBܧ�@�ZU*���*I#z|YL�~v��y�L��֛T���<�t�%�=�X� @N]*�e���tj�0x�y
e�"چ�Ҕ �������#Y��=h�C���cY�LGj�%�K����6������_�C��c��?�T�f3�¹��/��n��Q�&K��I�ܨ0O�,�,�yf5�|�y�E�{ B�����/����j�Ե)�)�*W�s�{.����+����� B��ެ���707؇��)�Ժ�~ݱU���퓿D<��uU�'��â�fX�j̎��f��n2����~7�|
[7m���e��O�`|r����	̑�]�P�8y���� ��u����W�p8P�F,G���� r�\����0���������W�I&E:DG
{������&R8w�2��S𴵣�&g⌯d�J�n��n��Z�����{Vu�ÜW/�n1cb��>�	��j�ef�|�Y�������S�B�P��֤� ��kV(+�D�%,$�\��*j͎3�S��vPR����'V���2C���N�2��D,B� �H�p4w.h�k^��܉Ĝ�T���s�h��TT�������ס��G��T��ݜV+���2\�M��Ui�T�j&����L��X���6�R�6 a�8�'� ~�466ĆGF�|�@B��`j5y`j�]�F�ǅƒ�o�Y��t &��d���\0�xxd��a?8�[2*'�TR)�r�{��z����(�3�4�5��2�r�#x��lZ��3[m����ǩ�8�'F;憇������&��o�Щ*��p�bw>"g��d�G��T�d���A�j�T:2R��P*��)�p�e��<��7�B�ԨVQ	-1�d�ИMP�-��j�`Hc�i݂c�hv��>� &{:��[����}�o�����<�ؾC�������~&D��:�E�&Q索��-���2�)N����G�=8�yu�醵�+���ra��p@�hq^�eu�N��,�@��<+����'z�[Z�İ.�rU��ő��G.s���gi�;���1::�I%�[i�nZ	cu;R�w�N �z��U��޴��:�1�,�u]B0A#�����:��d��Y��%M����OE�����[gz���%AW-�_2��&Z��5N��^���j��K��<�f�:��Ԫ��yy�kg�����O�;�>��x��p󅶣�^�&������F��ɝN��-���5E�� ����"$m�cg�,�3��T �F��6;�5:���=����~6W�qOD�&r�dʗ�b@�Yo��h�Io�s�����k��j���I&ӺT<�hvvʄ�'� �7�/';/��I䒫T}���\�LKd�2������tPL�jfd:C&�n����}�k�%�\�'���u5L'�O'���Cv"Ǧ��Ӳ����8N��5�,f�s�Mͳ#�9��G��"�� ��%��ON](�T���p�5�[��jW4)K�djy�^�&�� Z�8*B^�Q�S��Y����1ôѹ��KH$bp��EGC6�+�|ؓ&�Y9�-��@��>�I�^�x��;��}y�q�ٷ�o�8��f��0?��)��I�Z��4�a����p[�x��?���8�����h[Ԅe+�"	c�p,%���Qf<42oAI���J�S&�����"�����8�����`XD���@��{O$	i��=�'ńş�����-XJ��ѱ/<�5˚1��"@^��)%4:����^��=H#8w�������^���[[��u8�Յ+�(�o�N_�3�� 6'4t�V�c�t�l_��a�ed���m��ڥqtd�tmy��[Vl	�yӫ�{x���W��R�L��˗/�����0�ͭZ�Ve"p�U�D�/���AN����LC޹�\�ז�
�XL�Ŝ�n�566~��Ċ8�uq��1S�&2���bA� �3=�ie~K��/&��\�:��,%�/d���W��:�D>[d�:��#o����ϖ�"'�)�������9q�N%�����u��yF�6}��Ii�o7*/1Q�p��Ҳxut����d4��Z����*��2�(��sYM$i��?�l���8}d�ylkS�]s舘�3o���v���̓F)*9h	`iJi؍FE[��l.�.3�x���W�׫�F�Qe0�F�A�[T�|Z��D*E%'�Ij=y��!��E���b�	���c�9y�G�B���g` �y����ơg�Ic���F{5r�9�9�ʭ��,s��O��8t���a��������19I  ��@�ٳg�z�J���bt���c�ںBX%�j��9[n?t�\p�����a�����}"�c4j�\"C������{��=� �D^��NR�c3^��v��~���Q��޵�f	�n�	'.���V�?�	�X ��VXLU8u��7��au��2�`5i��a��u�����#�p��
n��1L%K���o�hb ��b)Xh�qw�60��S�a��Et>R�tၭĹ8x��VOB�X�|���i�n~�{@IhT�E9�.I׭ vA��ttt�./�|���M'������o��z~����ܔ\fG,��T�j�5Z�&k���׫ ���)O�'Lz.Np�����?���sP.�.�LI�sW�;�I�!?3%��G+��I� ~��I��5�����ḅbW)W��R"�%#�H���a���S���S�'��Vƺu�&��9�`vc�g+H�o�2 �D^Ұ'ʿ��Y� ����v�|�<,J0'��Ԧl�
<۵X�]Fn*3��^����֦�)�uR.���cPL��J�[&�b�s�^�$U��_��N{L�^��8����*�F.�K�H:�	�}+���B9F���(*j���ތ݋y�v�%�v5��sShkj�W������w��J���v���E祋P9���s�`��m��<x��wKe��܌d,�"+�F���_~7�[���A4�5b�;q�CH��wz�Hf�AP"WZ�*3.ʄO���{#f�+QG�U\c��/[�L<�wR�Gu���d��"����y�Zl�i.���������h���go\ׁ�d���v�v�ֶ5���R��,�:���@�������c��Ċ�:̒���
fU��/aN���^�Yg�L���[Q����ޛ6�E8��?	��ŰX�{����iQO�i���2��
%�]
�s��V�i��n��j���)l�;;;'/_��n./wО5�V� ��k
� G/����Z�Uf>ک���lS���k��c2�٠Kd��65;@�j�8G\$Mį�>�L1_q�
��=��J�/�\#��w��TW��~�B��yi*-�Q����h<&�Ag%pPf��p��R���g"4���7��(�w��k�����:6OT6>�kH�X�~R�ԨիDa"�TD�ߜ�33�>�����5|g����Q���ҏ^۟���l&�oME�I��ܳ��f�1�^�7�u�b����Q�hj%�dM(ɚ�H�i4��O$o�I��zZ�l&9�,���ҦX�t5.|��݈���{��Te�5R�D����8���)��ڈ��؃�_~��־р.�����(�8u�mx����ݻp�ͽذanٶ'�{��J����^X-&53P4�L
#�����5ԋ���Q[[���Q��#�sp������B�/���n-�X�=�i�&��񜏑�i��� �at|F�w��}v��}j7����
ED�6O�S�u\�p�o�L�}dVܰ#]K�1�`�c�A����{sᴘ�!s���ă�n��߁K����7��Ƴ�=�����w��� ������_��UHdNg�r��qI����>���!�W��R�<ٸqc��{]g������!=c�Dx?W�J�K@u�M��Ʉ�������nm��E��گ7#�TZ��\W :)L�TL��D�A�Z��q��(�,�d�)�rO�8�F��������Q�N+%eM�أ2P�;���SLck.	�`�Z�i��L���3���l,�h�S����$4��p����kۉޟ�V~�P�	�~�ĳ4�𐥔JEI
[�FF�k�<��GY�J�Q�cf�%��k�mz���V��}��Ku�u�OlY����߮�����ǧ��Yڸ�b�\�P���������U�ܗ˃�d�����琝����󸅼��ΣH����Z�He�X�~������z�;�પA4��OcQ���c�]8s����zz�e�&dSIQ8�[1=Y�L�+_��ɦ˼�~o�E/�����tw]gt���=�װ�Q��{5,�]����,Ak�����h������u�E�j4��J2��{������$�nX��>uzfB]B��K}�
kZ\G�7���������o~�;
'����_�v���-�5ȡ֪Gj�Z�	��|�N���	K�-É�����è��E>�G{�b�����Ybsa$�F0��m���[\<�)Ii�����@���>���uN����e2���}_�
}4�T���:���D�������+�O����Ϟ�0�Ӥۊj٠�r1��T�"j�u=�v�R�P���bQO���Z,�o�8��Rj����՚�'�c�;��5<��v��$b��Y�2�zdt��ZC�YU���eh�GZ��#�����Z����"Y~�IT~�7���	�e �F���Uf=�Z�U��eԩl��J_�����y\��Q�Kn�$��\���G�٤�}Ն����)VD����������i�����=�5o:�K�����sJ���{?R�q�����]2�]��#�42 kc-b�(�Wu��G��_}�G&�Y[� ��ӱ��_���av�
:vm�������QSӌ�ߏ��l�z�XÖ�z��Ί��8�)���[Yq�Gw4�+�����`JkVZ\��```�_P$��A�_C����E�dA �L0�x2��?�"�!x�6l\�db0)9xg���Ʊ��!ٝ�]�z�]��t�bR̔ȕ������qad�g/ᶻ�=����ٯ_A�-�r�D8O��W��l��:nܲ��5�����pW�zx�h�,B]M-B�i4�ߦ">�X\&����K�$E��Ng��޼xES �D a�@�d���=T__�=<8�)Nc2�e��1h����<�c,����r��w�8:9��D�f7�Sf�9�ȥ�1#�'�=)I�2�q��UX!j"�m��|NW�,�Xd���,,��6Bcc��V��M�B�6a�U���2<؆.{y��z+Lz�<���b��\:��p��ǩ�U8gW�a������D�C�S�����L��+(��M�3Cc,�e6l��F]RJ����eS3!}F�_b��|a�G�����'����wI�l�S���L���.�����i%��
v����<������MFj睻Q:k����b��ر�<��+����bu*�\��jB>F`vUv3|��ع�xg�14:%���.\D��������rWG�0��z_ʑ�2��V��V���䤸Ov�]����d�i�����2��7�.���W������%rJ�P'N����$:V�a��[�"<�I��HU��k��`� �9݉��)H�,v+����M{� 4�Hț'�a"�D��'ϜC�h!��:V�2aȤ������	�$�8zx�-��T�=0���U�PP��lHă���@/���0a<�#�'C�tXgs�����h�b�_Q�/��C>{Ӏa�k:1d�Sux��ƔY��[���{�\�(;l��uW�р���J�@v�������A���of2ޫ.^��h�u�jc�m���ZM���#ǄG�vE��O�e5�Ӫ<�U�O+0�S4��K�9��� �!����1W ������Vk��YP_쑕�dps���Ecs�R�.{�q��Fo�y���q����PzI���٬""�_`d,fd��p�ü 8��in'*�W�s�|N�	��k*�i::�+��V�8;;�dxb�e=�����a�/)��݉���{A�h^~��������L���	�p���KW�GϾ��6�EC����Zl�r�Ϳ�s���6�/u��C���h���`zz�?�wm߂��]��m�`z	><ީq��AO�bb^|!��Z1tFSn)%e��砯и��d���Qv�S�q����Y(Z���hA� �\��!���`�����K��8�-]��KW��7�R.A(2��kV���?����xq�QLu����|�CPV�6�&(Z�v���(��J�BO �|��g������O�\:�m%O������b�r\s��E�K�G>[��b/����\
��{�\�^���"�i?���t&��n�3[^;�S�F�ʝ[o8}f:�N�3��f�g�ON�	F#�ð����*��������ӗlh�.T��~Ģ�t�H�A뫫7��|�F9��^S��tf�Ď����k��P�m``��GQ&V]��%��+H%2E��H\(��ax��y�dj���ya����-���tF_�/�~[��?#555�w��z؟�ZAf��3)2��B���3ssj��$�M�M�H�a���g���\��
�����狀*s��"T�$�_����ee~�y��b9O�)��MD0?C2�&��澡����a�?p�����?[�Yrf��ek^�ت6���ɔt��Yܳ�F��Q<�� ��}+~���Ѳ|1���ƹ'p������8p�|y�5�$���1c�+4����c7c���b���!03��(R6�r��~=�|�������*��d�9Y(�
-7���t�0k"��ۇ�е�E����<�ƍ��݅��+c8v�;�paݍ�/Z���/1� �2�hu��\,�6!�3�%m !K�G�3�T��怺������FE�=�P*	)�����,A2S�\0�U��GO\�ADGP��H�i@��2S�B�#�E��v����s�868
2�p:��[�b����W��˚���I����d��贴��M����ِ?zyp`��+o�w�|��{b!�p�%�����X#�Y�M|�����eB6�Õ)�AG���u�d���됻'��:�/	xlKT��d%�L�u1�m��j���Ȭi�ĜN�1{�(|(��B>�`K䟗B��nZ��M��H�A'�jZ���hh㕘m�hnW5y��.2�<�РNgS����%�^�����D�5�G��Z]*Ѽ?T��N��A��jޯ�XCTf5�=kʹl����^](�=�����Z��K���0[�/t�n[�q�|_ﶈZ��)�z.����]صv5d2NϽ�:vlـ�����ygprrO<�B��tAo��H��.��$)��c^49�X�ny��^fE�ˎ_~i~���$T�)pe���ϊ�RU�rarN0�%�&W�cp�B��l�[�i��X,!F�S��ƬׇGy��U���N���0���1��D� �
k��ڡw�J�Vڟ�!�1A��$����䶣�}��n�t��p�v7��DA�
^���9���}������{��|5;yezA��7�`w�@^>�N�v��9DSi��fTW׈v�/���7�^����x�R[հ�;�\~�dWخըKyT����F���J�T�$9�Qb�H�t0��F�t]�T�7>Ok6�0L��J07�S�Z/&�23'�J{tE'i�jQ������2�y��I�L&뜝�i�M~�h굲r�ʂ�f	��z%�V���ވ4ׇ����Ot�P@��+�M&]0,`�MY ���f�������T&�.�J�r݁J䕙���+��Y8D}m�� �ȁF�4�b!��h,E�y�ǇUUrQ��$�R!/_%ҩx�֫�����٨\[��* ��	�0@�)���Qh�:)�.��ލ���-k�l���8`���5�/z{W�7����m oW����#�w��i�ټ��zڪ]x��gᴛpݷW�{�������9�?~E�N��8y!Z�Uu��9�����h���wj�j�U5���a�ޛ�Xm�P{%���Vڼ8��%C�yYA]*	��J;؆M����{'`��D���<�7nF��Oݍd�$�en\��a܏����㧐6ؠ��P��=b�4d�~UH�G/*�V��n��k�&324��ZAuM���ːtF�D��2���Nl�D�+!0l"���#gN�^��<7�3[���ъ_�~�T;7� �"���(�:�v�t�xV���ɬA��lZ]ݪ����FEZ�T�� S(��S2�Ԫ-Yc��d���(^;r(�����+�� �M2��R��Օ�˵�+��+g���P�/�YQ�t�X|����Ҟe�;�>�u1 ����͜N����+s-�I�*�ef�r��$�{<'����s�4ׄ]�!y���8� R[kM�쎉@ &4���v����t1/��$bq1v�lw8p�F��|��^h����ǽ	)��(ju�B!����|Ep%}mԀ�Q;R�]e����e�Ģ n�1����dJ�F�G�[���;�{$D���J��@<���m����=d�g&a6�08؏[Wߋ���_�ʅ�X�ڈ�j��L�y���B����N����*�dU�#šR�'o�D�E��� �G�.�M�[��v�id|�Ĩe]����N&X,�rjg��rOxP�N�'����S���&����E0�H'ϞC�݊�t�lݎ�~��x��8��M���=�4�٨J=�
��t��w�Ey�%���S1�z���I2��r���Y�5�����cP�h�𼊂$�t��!�*8��0�y���l�bVP0�Mf	�LԶ�B<S�L�.LbۺM�x�nێ];��x�f�j��4�q�F�UWB�ݎE�(�� �E�Rh���-�B&�����;뫫'���ZIJaA��$Rq�'N��A 4ψX�r/J�Ue�~b}U��K���z-�6�N�,Q��gp���L���J�S� 8K{�� -�y}�R)f*g�(0{I.�ټmPcA��8� RUU�sV9�ԣ*/m�6�Q�����K��H �N�M��Q��U�9�AJ�%]8n��l��[0�!�?�ƿOgH���<"fGO.���HYIU��Ҩ�9%��f�	�+���*�F'�Zu6�u���/�Ə�:�q�}��jM׺�=z�6���<�����.3�#����Sd�Ԉ�"�J#�j�/Ʈ��ƙG��Uxx�N�d��{�8�L.����gP�XK��Z�������7%֗ #O`,h��\���ث��rQ"�eYx?��_�tHg3���KX�bZ��^U�p<����cfro>�[�E�\8���7�[�z���/��d��(�S�	f��"����tNpa���ކX4��=)nN�X	 �
i�iiƽ[7 ���q��98]m�rd��L�H��i���VD��(�V��d�����}509�(�K����RՈ��={�r��e�u�֭]�w��qnh
Y�n��:RNZ��<�V[Q��a���H��S���R��X��:��͡X|����q[�ctmW�PRc�da^��g5�\�a1�U�G+Ɵ�/�J�S���Z�JT���*��:�漍�Ь�[�"N�>��i8Z��!�x�J�T�-Һ�k�ey~�N��h��r����TX��� >�0!�;��M=U(�ܛ/Ȑ*��9���=`yj�C���%
�Z�Z.$�{z�Z������C��*UF��4�t�*����O@����o)J$˅qPʇ�Ċ8T5��H��P��^�&MS�k�Fk�F됫�q���H�7��;V.�C۷����ؾa%�;�&Ot� �E��p�V\�x5u�����|�ڵ�bNw�E^,�8�W��K�b蛘���K����\4(�D�絑�,���W��5�pw�P0��V�X<"�-B����S�����I�y�=Xޱ
k7l�����I1�;N��.���\��f��A������,��Ȑ�̦Q pXJ%Q��	�h�\�2��<����������wގ�����}7,��}��ՆS��h"���o�Q3^���HX�n��;-b5{lp[\bz���(Z�l���o;��LF2콙<R� ���bh&��AL6��S����n3�\�F��p ڒ��U�\dy%��J�E&���F�lI{����7�z��ћn���Ha�'Yz{{��X������@�
*D]�(��Í���R�����5�[	XH�l��g���ao+�ot:9�����)���(��Y�k�|��$�AJ)���"�N��ŒE��rU���&GC�d4N'ҩmv��pH�@�_��!$�S)$�Q�s)�6�[�`4Co���d�jbbrQrv�s[��M����\֝�t��n�NU�`t�r��O�1�W�l�ԕ�z�h���lN)�1���t6���N,Q��nIZr]&��KH/}�5NKZѪ���$�7�.^���*�D������lĢ�Ka0�q��۱�Wp��q477��_�"��� ٪�k�m��RɴX#.$ܳg��{�S�m������7֙��V'<��	����m�&}>"��<�S!N��g&��1���gh��@(É���'���i�Z��5�P�&D	Xtv��}E.�y�. g���a`u �ʉ��@��Q�ۍH(J���5=F�Š�{Oך���"�F�C?��S���VF(���t�b��/��n�YZ��x��	T�4b�-;qd輸��mAS�m~�rI�{�",U���5tn�H�0�;H 6�=����cr ������)��^����g6�	r���k���Ԍ��nj]�0jt:���I$"�t��S� >��B9c.�i�j���$�j��-�e�#n�e�TﳱV�-��l�� ����Q���N&���g�����8`��hJ�.'q0�$����L��)�AU"{����1Y�+JɜL���5� >�8�em˸/L�$�S��s����M�¢pnvK�/�AoT�lwAep�r���ox|���`3�ȇE�z��`I!�E�-�N����I�g,1%h����UА�h��kԑ��h1p�4���`F^X��B��"z癷�)��n ��!2 ����]C#[��	����DV�~2�T��F$R9����Z|����_�����Y��X�;�ڌc�bxp�o`ld��������_ác#�E&Z`^5$ST�-�׿�g����Y���t"��!O�LTE�
�W5zT;�d����za�T���)y�z|A�� 3[��u���{0���'	��|A��C��@�ʗ<�w�	�ކ_�}F�Ƣ����{��$B��*���>��)�#G�HE¨��F��u-�"��I��:���'b&��y�*��	��L#�����C�б۶n���:a\�ƱL'����!I��� \u�x��ql��Fl��S8{�5�Ş{w�`R�B�];�~�,Ώɋ�B�7��l����i."2=��3�VD�aT{�Hɥ�0�	
}wE%f���A��Lz?���a�k��`F>��VcP嫱�R���\���r����l �E{3�L�Gק`�B��b��#����Xl��V�F�Q������M�W��X��X]�X�֜�D���C��9�6--s��HC��D�.O�Ϭ��������K���8�F��ҩ)���3<:9G�I�a��F���h�K�����ʚ�:�j�1==#�8�G���Pz{��C�h5�lI��VW$C�c�k"�OD�:
r�l�<�4��y�Z[�i���/�Ew�h�Zd9�0O/*���y:��|�:7�41�m���Ci�k��:W*���dfN�O�3|���O?���hiY�lK��DCM-��
[��&�zޗ�-%}��GQSS�'�z��^��?�i|�ч��|?��ߠ�,�6#����D�K�G2�wmjjB(���}8�'�]ʕɍT�_�d�z�{�/>Aל�C>@:�˽���׏�g΢H�~+�;w���v�z�>t]�Aߤ��	�F?V��g��V����l��diڼ:�sr���Vҩut_{�Q���\Sd���\�L���W�v����PR>��Q�HY��d�<7T��gϠc�RX[1���w����7����W�$��ĥ��x>�]մOuF���X�����0�	�vU9Ds�'ɨ�	��H����#~�g�T����4q�}>O�����E�^�։xق|\��b�B�PK���٢\&˅ߨ��K,���˔��2)OsT�ԹB�埛[��8���
GMCI�Qe���pZ�`��Z�bq�l�DN�C��_�,+:�:�Psp�,��(\���=��K]��q�#Ť�MF~%L\�愞c��hI�i]B��v2&:��7��()��.��x�;�>80ͅ�"��ɤ\C��LjT�ڦ����!��a�C�}N>~q�.*Jg#W�Vn3*�ZHr�9��n��ʦ��[�q��N��r-֟:ӹT��U��t
*�LS��ڇo}�3�e�*�}e?9?
n�uy@q,��Bg5��c%^9| u	O<��ye/�ѽ\�҈���%/�M�ɗ��W�x_��7����=4�l��6R���!ef��R�I>8n�''�p0G�5#��䵇�ȥ�q�t���?|
�[Z�ڲ-�61�+C�Q��ct: �ۋ��,$��W�c��F􌑱-j��I�4�� �w=��3�茴�$TQғ1.d0�s�n��,����*<�e47R�ۑ
L�?g��~�~�/_N��ӓ��'C��
;�n�['ϡ��L�3<;�5KZ�JGq��
�w��ͣE��~l�q-�k7�y�R�.�����v߁��[��O�Co���>)�̠qq#�c��\�� �*�@6�Z��G�#�-Be�"�-���ɡ|>��]=G[b��cJO��;���_\:�V�z�u
;B\?ÄCRi��kY�1�a��)�TF=��9�?X��D+u9�S��d�V�!W���R�(jP���-&B҈�m��.U�kZ�d|�����Ͷ�\&�K�*n���hIi�u�R�ʤ���NFIm�¨��l5!a4�Ky�}dlt����)�,�LIV��d\�v3f��ۓT�U"�
��
pE8��e ���dJ����1c�F�c�����z������������%��͞��Lb�ۂ;6��C�o��MB&c�R_��c��#�U�Ł%k:���A�������0fK����v��|�x���|
��*|��?ß��g��羀��,,t��l6���*��Z��:�%�{v�U�rV ����FG�RVc.���]����]�����r=�o�L�g��A��7:ǅ��l�{�/���$��:d#)��S�辫��z^vojiC$���\0FF�\"ŝ$M����� wlY���>4���q�\�ҏ$�щY��^=W�AC�F�V�������o����e��ڌ;Y2ZɈ'�`��AK�at:��|:,fP�U����7��Ka��aQt���[�͆�9<EcB4����%eۗ-�oz��}At��1YK߳�f��>�c�|:��ܲi���"��I�:��F�H�X�q�]^�0���g���r�teJc�n��ǝB�~�X"��es��P���`��#Gy�fsI��]����ʿ���Vd�&�+gK"r��H��Y B�ڜɪ*�P �M�&|
��%�d6Y��r:�Z-F�6yzRh�2���W��7�3�}`��(�}�����:��T�q+�C)��F�| +�Q*у
��DF��x���kT�2�;r�4�]��ճ���K�D&QMOw��l�Cm4�P#�c��ڃ[0�7�W�~w޺����5�O�
�--�}�}x���a�q��{����q�ݣ�k�-X۶'N�FӲ�����
���Ļ.q4/�����z�����(��0���&�*�-V2dȲ�,)G�<8В��b˦l޲�O�F���t_��b8x����H7޸���!X��$�V��b UB�?���t5M����Aͩ#0%%��C�Tь�R����i3#�A�I�&���Ix�&ql��`��/��_��X�h$�`,5��9_%f�ӗ���p:17>{c��~^;~B�$i�vVD��qe6ՑN�z�V~����dxKZ�5�aL"�aӦuH�&��Tx���1��g��0=�CkF:GQ��ʆ:��q���F�:��*DgC8�?�h"�q-��Z��H�w[�RA��&�H]y����yQ�T�1��ʼ�J'T�GEG �A-��29LrvS��m�v�c��*�C�W�
~����L+Q��c_fF,1��8�F����'x�w&�G�hK5��ר�ka�ۖ�2)N��A,��Y���w,P�;��:u�T�{��x�y�?0R��Y�A�Kg�{]�ڎ(:�$��(�R��d��ˇ�Jb��<��K%�:̠(r�j��6w�to�28��ϟhp`�����M�dv��ڡN�Chq�p�m[0>����o�q�2�ho�p�t�n��Ͽ�P<���B��W��?p=g��Dkt��Q�>H�ܪ��0.�s�A��^W��"1�藿�W>�%|�+�������e���]9��y�����R��L��J���[�j
�IP� ���u��h�C#���Л4ؽk��KO���ϼ��d�'gB(�=%���W���C�,t߸@_+r��K�مl������>�@����O��wppż��w�J�ü��Gy��͛���gM���}e�K�����kpe`��c��6ܷ�V�x�4��nw�ۗcvh�f19�D2��NFS�w߸���s�X�j9�� ��X�_��*���nZ����X�18=�E���La`Ƌ*�'�" �dN�h���D��P[�Z��umMCu�?�h�']�榍����R���2������7<�¼C��=�/#ͷ�!f�+��5����}�@��~�s^�+���.�GNU�%�VE��!SIT�*+�.�[�� )� �!��4�}Y R���D:�\I���LΦ���rI!3��Z+E ���Q�A��Y�6����O;GFo~w?��>�'�r�>�����RQ�B�k7����2����4�[\9(�>t������d���N ]��OП��J&�G��6�>�s%F��lcJ�gO��_��ݠ��,�T1�
2#��+ob�����a�J/��5�܅.��$~��t��x���p�,y��o@� �飇��[�����|g�/��+g���=��g>�_���8��F�꥽x��=��׿�_=��bM��*�[�f
�"�&"� ��(���ػ� \UNQHw��q��)^=��
{���Q56�ƾn�z�mص��x#�љ98�0��FS���b�A)���m�q�Bas�JoP�睁B{ĥU�m�Z��/=]!��.�do&F'��5;w�.^�C�ߏ��)R�Qh�5%�d�Hkzo&O��a	�͊��.�j��~���5�k�a_�
� F�F�FU;w܈B�����Ջ�W1_���o���	�X
t�N�_�	�{�e�G�����S�Q���:d��y��ń$G�\պ��&�]^TS��-#^���P� =3{��H�~1�5_�-RIe��
�1��S����cD���� ��nL�uFc�ɐ>��#h�R�8R$�qU����f���6G'�K�ߒp�!��n�l��Xr{>��������,��
�b		R��T�<5�(@c��d4"B%��X3=8[��zOI#i�I,M�C��̚�s�*�_*��J�A����Q.�l�9�S?�lc�ȑ�2��Z�gr�D"�>�׷,���'�g���S��.	Gc�zO�&�͉"<I�:�Eâ%��]��(�����#&�&�i��׾�8��������\�cIKy�4�ў ���ݻ���&�E�A��?�}��j�]�E�(�Ͻ�����?��~��$SXT�!@��� b$��i���2Y��4]!���?�>��?B��ǽw���l�a`Ā�
g.���}
'/b��x�wQ����������9b��TjR��rm�Ak@��4�I���΅�P���}���0j�8{�]�~�V����Ak6>:��y��1h�s�W��W}s$Ġ�CK8�ˋƛe˗���Lq�#d���_����_� ���gQ\�"ɻ�w���]w!�b��;�݉��:�MbhxV�[�n��)�W_�қn���������0<�1�� �s��zg�hSK�y��8Y@0��j�%�����@��\�/0$~t�bċg�k�e���^��)�haQ�B�X��}�eFd Z���#�`@D�\��c��|���S�G?�Z�4��R�������F��a+�kӲ�b\�'��8��Bz,���2����������#�)�P�2�r*�������Ay<���̆H�_�����i{>(��ҥ	��Y}z��弢R��vpQa��� ����u:�"zP"EZ��T �G��#��GD��*Lg��ƫ2�\���1�O�(+WBn�����D��5�M���R���>�>{��d���)lZ��}��d�����˗�Ʈ���g���Ģ	���с�'O�w�Fu��l��H?��w����o����~�v��~�n|�k_��?�	F�14�kb`����m���V���0Ʀ�`�7Û������m[����;�։�2��%�����c0ND�李rԢ@�=S(BG ������+�P>ϴ�*�`s�eh�qb.M)Kϗ��I�O��������p�,�����u�q��b==M��ب"���@���Ӫ�רD�;��0	��0=1���Ehk��Ha��{�jY�/?p/�>x�4�n7���N�.[�g��HG�v!�����ԷcŒ�~3x��AӒv����xu�s�&��޴��b^L�+Ĺ]́�]���j%���l%�~��GO�6޿�%�:q,�G.F���l�鰗	�*��<lN#�5bБ� OB4M�m�[�+��S
b��<p0u"�����'kӑ���^�T*�������� ����I5�����g��E���*��CJ���o�S�٧��:��,��	^A=�ː�,"�N!	�E��$�a2��x8L�Tj��>95���C{�-C�s��b4ڳ�\L�Q��o��^�앹�l�9�<�c^�7(����|�ε�����"��Ub�E� �����F�PK��?�l�	�k�Q.����=si����A.�.C�x$���9�����@؏7�#�ib���O��+�m�Z<����OBFT��w߅����F�@ߊ�9L�ԃ��ځ���_a��w`��u�=��T@���K���O?���'x��_b.��NqN*b���a�1H��'0K����h������7���>���Kx�ͣ(jB�2@lx��F����WyH	�g�>�o*��"&�ifE�{h�{����é��7�Æ�Kq��א��czx�|�~�n�U�~x��������! ��&A����T�2�vg2D�D@!�!���%����B�C=���ٍ_8��/wu�V����q�8��^�N ���[w@[���a<�˧�y�*ܳ�V�階t�a��{q���0��(���'��8�W�Eg���q��Ȓq:�]�9>��s�\�)ʡVI�� �I��dX�N��H�X�!��Tj>���!�+�8���F��|TZ����Y���!�� �gҪ4*O80]������N�^۾�OGً��hO���8�F��G��U5>�1��D,�;�J�dUyJ#�|2��J&O(�H4J�[
�v�U��Cs~�c`���]�}��>8���U�vcZV�h&���y>�jgA�eq�0�a�k��,d���,\��+#�5�CĆ������K��[:�ob��O8`�؆�W�s�tV����Vk\���kr��_H���ؼ|����GN�MF^�-������A�)X�i#��/����:
'yK;�u�t��^�V���'	{�Z���A]U-���G���C�����\Օ.�W�:u*��A�V�9!������x��s�̛7L���<��IƀA���Y9����9T��
w�]]2��̀�z�O�U�uN���Z�Z{���C���͟܇����s_�?�T1�]�x,-
�b����b�>z
�ь��G�
2�CGN
����Z��w~���%�)����Z�\D�i�Py���sZ��iB��sgJ8�:�W�]�-W\H�h��C����9s0�Ƕ�O��փ�.������L�Zg01��4��hv��\�d:w�Ã��q���͛��jr��z:P�7������}Ȅ�DBx䑭��uƇo����O�r�:�^�ǏƎ�cւx�V�:yC�Z��1�?�=���|���M \��%ȕ
uIA2_�wL��hjo"S2f�J�7�t��M[�A\���s��3�d5+g"9�`E�2�AjN*I6���mR�9�<�.��5���b�t6E��zM�br�]I������w$�ET��-e����ee[Z-z}�T�N��7�)p�F�۝���2��?�/�R}�Dޠ�	`����4�$�yY�N��𸽢�+��J"n<y�cm___wKK�[F5��O�T���^D��!B��J{b����|	Z���VY��W�,T��4fhq3�� |��+�\��g��rf"���L:�����z��AF��]l-����r�/	��v=�ou}S2_4p�Z����_;�;(�_:o!���#t"���E����M��khn�GF�{_ߋi��X�d]#�����s���װ�y�.^�����G�`ޜ��;>�o��s����[�G)�q�-p͘��G�"J�4��(�U�qֲ�p��8�5ȦTd"I$�Qcؽ��f�F�0�_:�HR�B@��]'v�vr�Г��S��r=�b3�]�������!���\�v+��}���$K���s������p���D�WM�#hd����m�I ���a$�iV�"�K��(��E��nv:�F�8��-@�m���s�0Z����\�{6���C����o�g>�7��:t��c��Ch�97|�J{�{����k����|�q���d�ї��p�@'X?1	�h���.U�\������syc��E a�_x;�_�8t�!�LՓ=�%bt:�:�3r�I��A��J#g
*bLlx��L���)��l���iy͞Le\F�q}��RI��_�qUlb��Lp�L.:I�L���(bd2���[c
��Q�1�y�%Iћ��EM���x�d%#�:Z�D12Ѝ��dTM���NQV*��d����w�hg'��%8�I���7j0�h�b�O�;ӢXI�U��Ş�-�3펕m���/m��d-BEB�ۓ�t��V������o����"}v�/��k�N�$(���.٦��������8-�>���pxq��;��7}�ο����O��Y��j����������-���ۿ�?����� �͟���V��as��lG;������ي�x2#�d�J�h����^�#۷CcZ3�9#�(J*�����f�����Qr�/��@,}��?��A��i���0�b��H�C0���y��˼5@NSM =�$M�� ��n,�=3Z�V���hh$��b�ldE��b3.<,�uZ�4o½9�,,��kz#"�$�6�VT� ���Ż�U�'ػ�V�Z�i�� ��ю�p�Gqɚx��ݢcal܏����Ⱦ|��+q��^=.ZfWݰ��p5��u�J<��QtMDQ���d�F^:?r LN�B-�Z(%3����
FY�,��0X6?~���3���Ri���m��~PG}}�|�h�4-��U��do�f��е��B6�;��5	� b{�[
l� T�+Λ�x�T���k�Νt�a�!���VT��l*�J�v�M�����i���S5oS�������z}���j�`6��:#M4V�˩�P�l��pj��AmBx�#��H��1:>:�tGGˤv�[NL�i�(�1�J%���&�E�t$T��0-�r;c�а���5�$C�,p�3-ˌfz��
����c`iS��ˤ��p(4�����y+W��_,-�$�����Ѓ�|Q}����M��-o(���D�|hn��l��'0�v��(jx�W{�ѥ���~l<{��+��O<��?�i<��SX�z-j�.t�ߏݯ�u�U�i;���a��s�+.A�D
'G08\��p����0��	���������og�\��>u3��!���G�d���m$��ۼ�	F��_�L�Ձ` ,�XL��d�� �����\,
}:C̏��n��Fl���&��<-��n��ǰ뙝�5s���#���	Vm�����9^&���2����p8-� �bޤJ*�	��hW"�B^H�"�?����C�2�L,�DΏ�ӛ�7�c�����bɆ0��f<��q\y�&�k���ߴ�J�x� ^��������ʻ4�eh��U�.���;#��Tv�bBz�*.��W��d*��Nm1��  �#�Zr�^�˩7*�3���$U�H2�N��~]h0�t"sP�(T�4y�Tj������7��d��w���TS�X�~�Sl8������&�+Z�j�<���;��=���rz �)�
E������(Z�糈�C���p�"U�"#o�;PPÆt<�r������m�otX,Uy����"IZ`E٤H��ʄ�W�"V�H�'{�+=���_~/���� �s ��,�˟+�Y��1�Lշ��\2�ٹ��㒙�Q�+��(Z�sz��Ju��$���fݸߏ����j��N;���p4H 
p{<8|� ��܎��x�6n��훨kjF�@_��8^<z-K��Ʊ�'p��u}S[԰jn+��i�w��f)⯭F4��b��"�PU�Bl(���x��¼�̩�������'�Ķ�v!�*!洞���a:��5H��MVr�I�z�
�)�\�N�c�(���ji�s�r�|�yh�����W^A�����Ӹ����|��-2�(/���$4g96�P�sX�ز�FN=A?��^D"!�\�K�v]�%��D�q{��&p���gτ�N�b<LQ=9�,�_9�p��0���'�ō����������O|��x���x�D7,u��`�$6�1�,t������<#�k6�D��h*�@ �@@K�ta5��y�.x��獩x�H �)���G(2�M���m�x]:��h�L�se��#��b�Q�3ଥ�ՐIe�8��V�Π��Z.ȘΩ�BV~��7�9M�^D��9V�¨l-�p1T�)~�~.(���JS��7�)p�Gc#�i��v�;S���7���1�P���[x����IS�U��*
s�E�����雙p���@�d�F���i
9U����7�,) 9xn9��,�ڸ�d��$���>o/��B�L��\H%�*���k�l��ҩ�cphh�p ����#:����W=���W�C�����f'��k@O&����/���OLM���g����*�~��1<4��'�b�ri?�z�����UK0o��<rUU5HD���x���`�p�����D�]"�Bov0�5J�9r�ӠPD����{�;��9�,9A/����G�*<U�<T%���L(����b�i��%�(E0�$\��4W����ݢ}2� hC����7� �#:�}�C��I���L���L�;�L��E��dGV�K�Y�vLL�9��MN�V�%��y[M���Revu�G�p�B�^�;^|i�_�<���Z����~����7�r��"���<�����!��CWWd�Jd;��f�Ԕ��\�^��e�u%,�&(Z�Adĸ�N3���dM�Ѹ����<�]��kS5�0��KϽ�Kg2u:��ج�dqr���1\����
�1e2�L&u�����C.�3��+I:Y�f��E���T6+i͈�^2p�Ak�p6I�=�dw+5
��
��T��e-��M!�iL��w8xk��k̿w��'i&B����[_"��]\O����(��E��_W�:M�XG�s�92�t���n�ʷ"*����\i���
��G��EN&�U���_M'���&G��O�<E�\t�ؐO��0qL:N?�P̥�v�#jN"K`���Ψc�gty�k0��P��`df��#3J]]ݺY���+ߧ��t㵏��۴�}C�nl�cFO}:�����᪫/E 0�mO>
��ǖ����E���CB_(�K� �d���w�(�k?qs�/$?����<����z����J��L״s	�F=�-M�e9~=ܾ:�3��ދ�#�طgwvCr�'�ftZ����c ��� #S��C�N�`��K�� ��8�������������t�L�v����{{���p,ݍ\Q�F�& �l�%2�i:���Ȩ�i�-&3�h�U��٥�0�F�!�~rc�\�R��5� �$GA��\����b`l:W�輭	L��vDJ<���p�J�F����0k.����	��R�
�N�N\V:GrN%]�����ɑ8:�뭱�wl`Ȑ��5B��f��w�=�����7tS ��0����d2Ӥ(f��*׹�>�X��>;_
�E	��ת��&������z"ea7�;���M�I����P*X���;�GR&�Ϥ��ʒ�l�
p`����se ��5t�Dl�r��X�+�����1Œ��1���t�f���FFF�	We�I1�*d�t)pD8E$��=��x�iS���E�X<0���#�Oo��Zlٲ��;�����l^S,:��LPS�BP��hJ'�4�Uѣnw�`&G¤9��'�U���ip�з�V6#0C�Iς�yM���W'
�D4^540��;�؃�E��o���巖JC_�܍�~�d�u����aZkA_Tܵ�����S�Q�Dȩȸ�ӷcFC-�~��M��[n����+
���}�`{�Up�HE	Pѵ<q��}>j��7>��=Gq��-�ډh���l�Z� ]O��B��FD"Aܳ�y����̘���~Xk����`1�����fȉɠ9,4�����l
V-[�g��z{��cú�X�n��ك�/>�Nu��WEs@A���$��t�tȕɰn	4�+�ʅ]!�>�7.���~
8��#�Y12�&�Y��x<&�UH�\�Ja:����^|�֛�`�\̙��:��d�3m���I�	x����׬�g�O��F'F�'�a�����">��2�B��W���yD���<)���xKL��D\g�Eo)����9X0r2��� �o�1���?�Usj��甘؈[������;[�	F��L�s:����,�$1�W�*���l��F�a@�T��J����UU��f	%\���\�z�I�dnL�:��}c�XI2f�S<�5����0�֧[fN;�v����eSII����ȉ��D"��P�06�>2�n��Y_Peoǩ�%===u4��oU�X���i!��t��q��
�tߙ�C�\��eE#�x�/�A'��5r2��X� ��b(J,q&=�&�d��Q�J�#z�c``hI��O�`�?9&�&7^�ݶsW�cm_P��s�6��fua���F�cW_����o�'�z�5�`\�>47m���D ����zp��~\���ii�t��zp�Л��t�R�yA"#g��)Œ��VQ4����k�h8�$1.��z���B�[�ƒ��y ��E2�H��j��="�2�U��q�A24���7s�d{�p�K,D5oWԤD1k��Ğl�0�+���X��u�0���%Z=�3l�����u1g�tcF��)� X���)�Uf�T�"K���Ͻ��|�zr�N\�E8�=�*A[w>����Dk�����W\���a�Ͽ��v׽q��L8�324���tv:g �n�A/E�%r8L���kSy+���ȑ1GB���rY߉���L*��m.�bxm���7#5��F#�i�b�K�Pb­t:qFO�"��e}�yur���<q1(sq;��K1��-M=�X(�T�vKW��p&��3��w+H��E�J �X,�)L�tlU�#J�l~AU9M7�9xӘ��=���Fk|U��F��gS�&V���r�M_����#�̒��� ���E���z�?Yv��E�������Qe�T���C	��^��eF�@��b���OW�30����Em��S���\���g����d	��2���JdZ��dV���b$�T�+�`dF�@��`�4�x��I 3��xi{,u�v�t�_�u��ż����m�`#6/_���v!�,��L��$�ޱ�׭@��V|�_�\pn������0�u�\�QAGG'v=��7o��y��T�����.��͉��QrTE�Y(LĬ�V,^�`��a:M+�=�`���(Edv��v��͊���H��Q,h�����;�Ŋ��^~��ء��A�0<<���~�>Q2�ĩS����Hy�k-���5�L��0��Y��)jf����	aX�A��%�bΉ��@���̔^��KQDi��G_F6W��C'Q�CmC5�Ο�����GF�
kh�т9M��e2�`�1szb]���C��Gl/8l$r�I*�<m_��Xk����s�|�t�	4�`�Q���/������QFK���u��4���{}.��G��J QW鄪���h�X��
"��B��Q�Q``)D����8�� ������˼cO�\NUX)�����*�;p{v�&�,�j�t�4N�s��KF�9c4�L�_$����1��!-jN5�l����3�R�LV�F�Ӯ2�]iE1Ipz�js������W��z&��?p����+�fb�?��w�3y��3�R�<wJ�$*�X4����]��>wX�:�\tH��4�"3$�{���38p:�E�H�4��ǁ?t�� Rq�D���;�,0�܅�8���kL~��������Ou����枳v�y㚕�_=� �[���q��.Dba̜;��ux��;p����<�p�]p1�?���F�>|������˻�CӴj,X�m����m��g�Ñ���uTQ ��Oep��5X�d!�>���8p�0���a*P��:6�ǎ�>r�64�4���8�,��4E��}ݨ��������Z��G���������#(x6`�?�ӧ����#�_&�9���uB7��-|>�	0ɵl�+�_c�b�x���^E����	��ఛ	E��#�|l��r��ES}��Nx����q���uǑ� ���D���9{��jl" �Fkk+~|Ϗq�UWb�E����?M��5AA�Q(�!�?�H9��4G0m)��9B��$��U�=f�'�P�"'��\����3��W��J�]S]�EC~_6�6�v��b��|���(�n����L���3�2(��!{'�#9���I�J/�$7�h+$@�
^�w6����U5��d��|�`)�L�����q�+� 5��0��� G2HY�����1�4����88�{�!���e4��JR��U�:Z04Q̗�i�Y������	��)dn�	�>�M�O�����v��R����y��>�^ԍ�͛�\bg��3��\j�1G}�(E~��P���Nͦ'[yd���=�-��
��#"E/e�����eŲ�q�'��F�����6Mr4��r��1��0a��'�Ƿ�_��s��b�Q�G��H_/�Oo}���݀���?��5t�j����'����Wq�E�q�Go�/݊��.�/� �΅Z��sG�!���������`��
��=�86Ψ��/^x�5lܼ	7n���0��2d>�+�oA�Q�U�bl�.���(l��/$�Brb�~�1t|g�['��|N͛/�c�0�V�\H��Ң��
�ВVNTq��W8�����AG�<(�Css3��0�Ir��8�k�128�b٩��	��h;uJt>\��"�`p$,�N����G0k�,����ç0}�d�9z� �5����Ͻ�&�^��t�>3��q��A�-Nr0�\^`jzD���V�X�b�ymxKO/���&7)ӫ�4*��bN#0g�u��|s\��zy)�����.�x��СC����*��U���sCd����8ً$َ♀���P�u���N���  |�ɮ��z�߈!��c�P�IyI�N�9���.�u,1m<�i�K+��L�� ����u�A�5�\h5�4����0�\�������h��L�jQs�蹖�UY_�?�gxO�W]-��jj�0A�]�%��69z|���As��ǝw�Y��W���OdԴ�Q4�����Zn�N��#{�v�}�D<*�:��@S3���1Z���dr>v�E\ e�}�������ˁ`����g~ h�_�R�� a�x�U;Ju�����l_��/���~��oc�+/����Ɗ�K���8|��0f=��5�a���ןÝ�H��p��H%���x�՗0c�J�>{9~l;�:��u�1�ۍ�^'���k����|r�O�������cl` {�3K��K�ri
�tJ����QE���/Ƭ�ٿo�@�b@04���n���h����5�` ���U�B���I�梗�C� (�ܨ��q���ĬY��L�k	�.GG�D��χX<� =�PD��˕�F��������-ق˗b��xm�1��	��854��?���>t�5X����g��=��?�֯Z����|�j�w������ŵK���g^B$�f�AK���!� T&�"�b-k2�9�b�m�+�
9�reQp�
����bK"�7��r%_�sv�ț&���H�9	M+�J���(Ŭ��&����s�QM�:�.$UĖ�1W�ar�����+���+����O�{Ǚ�h$a'`�X&F�^qadNtE��T�:Ud�ҋ�Z�.4�K4'�6���$O��c
�c�_��������H:��
�\��T6�������9��F��^�6'���P<�9z��ٯn��,�bk�bqe��2�N��<R����\����3G��H���u�[A2p�A��*
-T�E�&N�qϺ D*���7J�cn0�(����pf|l���s����\�8j��O=������'?��'o��Ӎ��'����$3<<��Ͽ�"�,���"��6�_��n؂]�=���'�X�C�}2�D�(!+��|�9��b�?�
F�ؙ�3h����+7by�����6#,�<��~�����͟�>�����U<���p�֐öA�JB1�F�X{�Zܰi�XN��>2�y����}=������"���aQC�`Jm�^�p6��qd�^���`c�u`9C����O%2 �^�cp$ɿ粚�q�h�ϙ=S\���	T�T���^߇:�U�6�s6�cit���Ğ�>l��rl�h3���BV.Y���!��g/��K�CQM��t6�]��'1m�|�C��?~z�UMtO"P8
��%焂E�]�^pt������+���D{��H(fUȴ&�yU�To��?�s��(b{���A�{�E㳋���kJ8���Z����I��*V�x�ߪ�5x;Kl;�~�TXv�e%�:�,0��}���_��j-����ȒV%�Ӵ�27��L��0�9��D�����>�՘��`Ĺ�D���'h�͖$�Qd�BIdr�2m(��b��H��2������:�����׿��}���-��$�dj�Ntt��c:K�29L�5Zhbah��/��j����h��ٸ�	�V�/�9� �.XH�s���l!�!�ϭG���lfe-�F����=mR��=��P� aX��;~�����߽��?�|�E�o|�{Hø��+0w����lni§?�?��	������<��='��k�;�U73����y���qLol@jd��	l��,���Fv���	�K6�9X2�
�\
���[����+6����1�8Չ��*r�Y������ݯ�hS+l��v�م��Z-�W�f��C8y�$�Lh�/�'I�L��H0�!/
�\4��5v�###�����u��e�Qrlp9�E�]�Upׯ�CQ,]�[��CC���GD����}�^<����K`�>��z�.�z���r,[�/�|+�,�mDNoFdt5���n8�F\�e��5m��<z�C5o5r�̠�C�9�L:8gT#ɭ�t�jD�\`��d��h������1S$���+�u%Q[#�5I��:��-�c��Y���������skj~5
g7��R鄰l�x0�&oJϋ��!38୥�*��a����t�Y���H�� C1s�k�m+�7�≚��Y}f��A��N�8�C7�0+��Mf�2��L�-6k�b��'�ןsL��wi�Z8c|Wm�s��z���z��ad���­X��0�j�@]]�xN�GZV'N���m������/|��ܭw��I&r4���e�Qq��d��\F��9�����F��ș�hT��h�D�p8F��Y1��E;�P��#������Bo��	iMS���������]\�5������{~���?��Z��[o����o|Sw����j@��9��'n�����Q|������ Zq�g>�{}�6��u�������? GdG��?�ڊ�^|.Κ偔臤��m��^�Y����1�Bn|�kwb٦��j�\�?����j\���%�O~�S4��P=�h��x�>"���>w;dU��i9sd3ٸiQ�\�^���y�g�Q�Z���!��� �l��Ћ��F^G�]%d��084���	хsÖkp����o>��@/>	Ϣ��ַ~���~4�^���qt��\�|.��&X�!�%_��-8�;��/��a�y��-�($h;r�^~	�]s��u�u���Mߑ�#_�.�<&�E:��y=LF$�a0oGIg '��ROs�Y�
\Y�u""� �$6�cZ��}4�I}� Ah���T��A�b`e�{~��U���^١2��4U(1VT\�{u�i�����y���DF����^_b�ْ�Vb���2����;j�& ,'i��d&?��ğY9�<iܩ�-߼���Gt>�MB�%'ˆ� �;c
�{#�:sFoW��)�����fa�V�X,l�6B�?>��gd��T�0h�!B?e���ջb���u�y]�`v�+eT�1Z�Y�Y�K�ѡ���β���0<�5�v9D�a<��+����,������N�D�?(^�峂�#I6�+,K�t����kVxx���Sx�������>��������k�6ϜO��WL���wu3V,Ų%0����V2�k��>�Z�-3[q���W����n���_ɱ�`��*�E�ψ�[�KV�ª�A��p��Ɂ�(��ֺ�d>2��>�����l�EüذtV,��o�����g¸`v-�'?���]v�-���?Μţ�֥��pM�e��'��d�I�557 H�0�c��G�|�9�bm6�~:G�LZ����֨ӛ�vK��#Py\}��X<.�����`f�]����`?���� j��[�p2����}�c�Es��H����u�s�Ƞ�tۯp���1�y_y�^z�Y0��Al�V����C��f�`��gw�k�N�RLH�����rKf<%��d�Z6' +Zr5}6���%Y��M���yr�����svi�!����n����JE��j��x5�*oQ��g�ފ��)T�+m��*�s��"Z7���[�z��Y\,�?K8Ï`2*Z�H��50��1�d0�6�cp�$ ��-ݦ3�,���g>���X�4���;c
�K��϶����틄"�S��� (�˕���gR��8jsz"�˵c�d�2J0��o߾�}�w��w��rv}��R����m��iL%���]W,�!����%�逋P<k;LL�D�A/@��9{���"
9��v{	]3g?����}F��J�:]^�����ή���b���I��;n�u����~翮���_�������/���ɏ�z�|��W�C[>����{��+�����F4͜���3�Bx)�	Oc�ׄ�]�kZ�h�bC��Y[�Of�[ڹTS-�� ���]3�	F�Q4~�ea�����O?��	s۟~
3gLìi306<"���`S�p"&���f����L�7�ֈz�@8$  ���wv���Uhpd�#`2��d�+���S"��վ*�CqA@��X[Zg4
q1+��M�a8p������3�����$d��t��^z��Vl>����2iH55j��r�b:�o}�h�7^���A�k/���Vc��V���Z�h^6�6��w��c'�wzQ��J��[�	��c#�s:0CG��2�8����a��dVE�l���|$uA�=���K�?�s��16���3�VY6����=�|����Pd�����a�Wa��$�d�9\~��8�H^�MF�|r��[-�E�1�r4�ˊQ�c��F^˞yb�`�ʓ���(�<d!	��2J��~owL��wq�O���L;66>�KF����"
^���0j�C�����jF}mF�ǹ���ek�;v�ᶶ����Xuu����<�=�Ne�^�b40�x�ذX�(��"b��f3�f�,65�B"�l�J��
G��X]d��昐�6R�,	��P� N�|��L$[:N�l^���ᭅ�`�e2=�ⱻ�{(�����'6]sբ��S�.�p�f'΋�����������������߿�-�V8�r�1���O]{.5Z�d&������b��9�Ӂ��C&�c%���O�­�ݎ�d�{L �{�`^m5"��Чb����6�tvvb��FMB2;����謭!Z[i.��0674��<6�ӦM��Аh?dc.�G��M�A4���؄�4�=>D��rK(��K�b�E�ɧ����s��@�ϓ;^��R�y��bչ��l�F<��M�����x�k<������B������p���;��c�?�x���VȺ�\y�r��h>����.��i�r���F����4-@�ZWa~]�;p}���a���:̓EP����sy�p'w=0��L��zR���)6��_��q͍��3@�M�j.�L�H�d���V�DݑRQT�N\��[�z��>��p�
�S�Z� 
?��P�Ken�͛BL�S�����6ȣw�̖ɪ.�ͥ��e��l��k��Ѐ�sa-Z�]�m��Ť����Θ��I�fp��S�N�8l�Z�5ը�:���r،�������h���lƘ��9r(��ة��mmmc,������o���΁�'����f�h5��r��XU��� o#��@s{/X�_��XTQ�ɂ4Ei�by��������DT6(t�/	T��F_�D-������|$b������Ҙ,R�}�'�����=���-�,Սr�p ߼�A|���в��/���1
�Gw?��Pf9�b6��&�t��j��Q�!�U��^��P����6y���ۉp�@c2����á����Ǒ���2Kxe�!�v�a.���B1��t
W+׈(6��i���!o�O�0�/�	��7��G��]v�P�.w�
]-נ��[!�K�qVf��s|������at�{��M^��SϾ��V�D� ��cd�:1M�������*��REs�-X�~=���v�JE�'͆�e"ǔ+A��㦫.���8��KX�dj�n	�pׅ�i�k`b-Rd1�e	˧��dN+�k}���F`���V�&�0Y�3C(�s�A(�&�����#�|��[�h�&���ϸ��mOeQ��>17އ �����5�l��ֿ���� ���g���íl+0FE��'�<�ʝ-
}v�WJ�?�������k6����N��?�/���tu-<��0�'���P�s��.eC�d����6�1���]�sSs[��$SΌ��
��`L��/�l���bW̂@�9�d�cل\(�Ou�\��>ƌ��xM._�f5w�r�Rr4V���Xk2]�N����C��EQ���+h�3�g��柘@��^�?��9aJ��Ġ	�Io�!��u�V�����G��}/i-�՘c�'>�dJ-Z���|����I3����>��7��i�uB*�`��躰m	U^�rV��@��#G��PDA�%8v����)\)�Quv2��u��1��}�>���A�DV��n�p`��^,�֌�G���/��a�o+Z[g"�L
�ƺ�F���:Ud�U�uFCЛY�QC2C��Z�&0X��D6�|�Y8�A%���*�<W��U�e��o|����X�f9n��r;Չh,	�х��!�b�p4��գ�!׷"U*�*�����D]N�-��N��:�μ���1���M��J��\��⋱vVbCX�`!�j(*L���
(v�hΫZ��ݡ+��J^�s��j��|��׻���c�a��`�s�T�.3�*�7:��]>��d:&��v\&��p�{xF*�]�؎�c���<7�/s�2�_j�����ݪh��E��e�m`�� �������f���Q.�XMV�%��
�Z�BDi����^��I�|��1<<l��;�3	�N�QV��E�� Zx�
�%�PV��4����{���wcL��wy���2��[�v��j�M��L:aΩ�N���MD+�Q��3�@mm=�F����x}�#�.{Ou��:x������H9�Ju�a���G6�yW���X(����r�(Ōf�$��:]6��gR83�A�����C�?�t*��Ez���8��w�#�m�DF8!l�F^ 2�jɜΨ�;:Z�:�>�Z��������;?N���꬚�5��H\70J�5W���K>�v}�])ֵ�aJ3�a�R_�=X�"�jy�=O �`��
t"�$窅��}��m=~��f�J���r���h���0�yp+n��*(�,Z��G`qXE{����0"3ę$�`��w��&`b&2b� .4U	|8�>;]L�a�XQ���ŉ,�[�K��޾X�N��w[a41���/��^?�α�Qh�̾&��y�^� �78�y��?ϲ%X�j#2!���`����p7E�z:f.0��.لKV-á]�c����� B��X,�b.��h�-3�J&r����|�����p�?ց�}cP���{(�<6�5́��4̜-`�NCӽ�ϰX����N��J��;��x��?}�W�Z�Ƕё�x��@�-�-"P�X�iem��������ʛd�*<)<��̞�Θ�z��2Dف�|�1YDM��4k4}�o;C�����z�LS֡�n,ޮ�r��/�`�1>��(�K!M�D+Y�f��q�'yZ��c
�˃���چz�sJ�ck�Q��`0�،Z���P6��YN�C��m�	��oUlU���A���38�lբ���cC��Xw޹E�ħ�n���_z�����Jz2�攧LW�!�1�k�l&��a$@�7Xɠ:�Q�(J4��xh:-E���E���C�)��k9�0/gA���A��j�ztt|a��=\'��l\P�@���߽�W��Ӄ�T\Us#:�b�Xt��(�w�a*f�������8s�T��dS*0r��E4Y2�F��fBN��}�Q�<
9	�o�Q��Y.�˖4wt�;�K����)��IFȱSl������BV B� (j� �Y�39��EĊ�f�q����`o/|�tOe����G��b4`��٘9g!�}q7�F�h{����6\�K�"�1w�R��?{�T���*ͯP8Y����8g���/���x}C'��箘��/���+Vc�9���vԐ�^<�Z*	E��a�B�:W~����
`j�Ds��3��B6O��j�2,A��/I�J-e����	���"�d���T�R>M`�
)�hBtBd���Rm�q��w֣�^�C�2�~a���m=��$������9�DX�M%nafFU�1�ɭFv�L��s��B����ذ(M�rG�LD��#���Q�LjQ0�Vk�ju���"����;�����t�"T&���r�3/��d-�"�d���gL&�G��t-��;����a̟ߘl��r`db��j�Ւ15X�8h��3�"�,M�X$L�P �u�d����AU-�Ʉ^��ݽC+�{{_,m��m��{Q��SS�(��yv�b���Lh9-;F�1�N���DF�5\N;N�]!���e��ba�C~x�^#�6+L��yߐ�C�Џ�˪jd/�I�l�pha���Cp0I��Ǉ�{�;�\>9����yv(69�N$�t��z��������\5;`v�b�D�۟�%�,-=���A�����'�w�&\��!��đ!�o��p3�7r����?N�X��t\���g0�³\���y&��vE��*�e/��rʘ����=e2�i����*2�Q�"~���O�w�a��������у	b糯���V��'���� c��,�0k¡2y���D�l���F�şL�P(`�� �y
�+,n)�8<r�,�	�H��bf�k�-C&E*!�$����N�#�J��Y�<>�	p� �(��Q��Պs�77O��j���#C�Bʹ�#���E�;B�A�s!9>7��|.��gir(V��\J���k��Nx_�������|F.���z��9�9�&p�Jf��H��56r�@��	���t��I��eGD����CYcA/��8��$�B����$�h�MYs����6gry�Dюl�uBSC�ŕ&Ϸ�	�����y=pF-M�� N�@z�ј��+q��1��)W_�����ԱT:�8�+ҥE� ��8�'#9����A��C�׃��E�J�����y}�Y+V������|��},]k����Й@Y��".���n܉P�T����PS������J�l=�|>ܲ�k�Q��ǙD�D4�"�D�/w~��)������H$:�����J���X����Ri��w��ط�/w�{�j��Y�H�4c~+>���8���a���`3�ۥ��Z�H�ƃ�g~r��k���oN��q�C��ߏ�k�E>����\{����/�F8L�-�E���դGJ��a���K�t�ăA��ݼ��`-��%pȎ_����oH�P����7�X*t.z��煦���qr7K��?D&�}�݃M�\��j7ο�_�G�V���(:bx�C�O��7��R׌��Dߝŏ4�Ę�D�3����>��_�qﶧ0ͨ����PE`��΁u$\�u8�� 75��5�˂Q):G��u^�~�Ȁ�"���jo��Np�*��8�$9u9�D^{�׸q��%�� O4�uf2yH����7&]��J��,m�p"�f`���d,��&�7�g<�5M�Zł�d*�V�xU:J(�V�8*[
�;����N勺��bE~��tˢ͐kt(��R)]�m-.������Ρ���Q�OO�'k!
����L˔�:~S�T�d��<��*����)p�g�/�4ֿ�r$9�f����P6���8��w.�1���UOQ�n�n���Š���G�:֟��ľ�wE���k�;FG�iU�H62��"&��H ����'cqXl(��}d��� C&��PI�ztl�h�"�r1���*�\4��`�4)*U�V��H����X�o߾#tZq�ǖr���K���_���{t��R�a���Vf�<z�7�?�#��xo?�ͮ��%c|�Odj�SW�����t�����y��+o��kףm(���|����9�Arr�׬C$���_��e���R� e{w/�x6�?��LO�L�\o�F�$�tAT�Wl��վ�頑��y��@��i�\�-|N���(���)<��e�'~뭟E�׬��̂P��@V��C(���ֵB3[E���ea�9���wѹ	T��!�BY�Y�=n�@�:њ�ŬR=j�sr��@X:���aR�pҼS��� ���1��n�eg�u;F�yVCu8��B�2��܆z�^\�f���w��]��J�&�ۢ��B9�^0E�z�v�F뗀�NM곩=W_un�����_|<`�'Ͳ$;�JYU��k�B=#~si���3 �;�3aȶ�{8�����:(�
��l���keE�r׀��N�$��\���`u�X���-|���W�0���փb��.	@S�k6�-�pXc��wL��?Ө�Bj��%�{���8����D�*HBXV�S��QN�0::���0��Îx���uZ�b	�+�ߵk�dD��U���&���N�T���22�HQ ��e��X2!����9z��Pp:t��͈E�uy! �-��n��\dHMh���s�^��2�	���&E��g�#��[�><*[�/��Ŀ}���ᱛ_x��ւ޼r�y����6��k��P��Q�jfPD�ENo+���kq�c��d�0.���ܫ����g^yW�p#�>�R=]ؼd6S�>�@��4��n��6��P��瞃ݒ�����JgR���X�V'_����+w2C\�R��a�fr
fB��������_F����������;�:m:6n܄�?�ކY��Cې3ۑ��Hq��Z>�����b@>��t��_s��hÃ���X�5�c1����
c0վ��.���-���~+W�G$�$K%�BZv4L�\9}������n4�6��������j���	 11��
sI��������z��P�w���Xk�����~	��ixk�p@.���rɂY_1����wn>g�����`�֭R(���ff��l�기U%�ǀ� s��3�&[�+ʋ�x3���L��6�dDf��#O�VE�jP�
9޳ &���Ga���/���V�$}`�,U�	 pAbnR��� Wt���D���Z�]6�sjK��)p�g��������{*���1SS�:��t\�d��a,p�@�hV2D5>'9f/-$�QKF�7��g�-;�m;@;���ٲeK��;�������յ��,�)���!�[�_�t\�u.��9�{G/@��b�(�R�j��.�*��=/��n�s�nn^V���&m�����Y�v�Df0�ϙ>o�0��+[�ߍ�'�_�D;s0����v�>5ECtF���6-Md\�nX-e2��]ȦT���E`2��3H�a՛����&m�l�2�$;Y΂��P���d�gtl�����~̈́�Ga�e5��W>�Ԗ���<ߵ�魽_��Mf�^���+�bq�?9ы S�+�=�	'���ѱ`{�)���a|폿��ݽ�o��n��n'���3۱l�R��������^K��d ���!l��*\{�����Q����"��?g1��H��	��̳$�7��[��⨨$h	 ��u�V�ի�	�O�Ε0<9)��_}�]�t�Kc)�jx��K�}��L�le���R:��� �4��q�B2a|��k��v��?ݎ"+*�Ϟ���^��H)0L͠����"���ݻ�r�:,6�����|7�,�ZUƩsH�"�(I�k.��A�"RɑpT�N�Y�v�	:rV'��ᠯ�*a�	LK�h��Rc�d�P\�D`چN��2vnx�봽tӆ�?{����}�����t�_��]���:���7�S��~��x�ad��Z� �)fM�˹si�>�ȋ�A}t�^v����u�r�9�Vɴ}��tjp��D�5j��^K��;$��dke��VR�=�����Lg�*��N�?�vS�[�����jnn�>��;g|��3f��%���J��ei̗D�vzj\4
Z	 x�vxD���ʖ�Xb�;��^B?t�{4&655g[��B�P���SC��6��"�D!k(0�o"��� �D>�ˎt""T3t��P�F��m�٤��dbL|�3ٴ�q��-St*�j�<cLơqb|r�a�$��G:]W��n�?=�CS��|���{����KՒtx�;��o�5P���y��05��_��C�`�:;E@ъQr�+/ۈ	�4h��k�r�􌆇Σ�q�M�p�}w�����ϼ�X��Oܼ	+7����'�	��"eU�(�����pnU�
j���������	 �z�!4:L>����t-F�a4�w`�â4�����^���l��ðhr
]YOƿB ���r�6>w�f�ȏ�h�cC_�7\�'��Í� 9�t!��o&�\��������Gp���"��"@���;{�W�9'��i�t4wu�L��f�#RL��D�����M]�xg�^��s 9��*9,9*M��j���4&ud��L���-P����/���^�n`�GL�)>7��VN�۳#eG��w�$KdfE��_�Bz�Re�xlp��@˄Cz��g��X��`�k���b0��[�\���
<]���J1�g�8���q�߯h8� @��d��S���(y�2JE��������o.s�k�8�^+��ٹk�>%�\��E̘�,l�2#n>h��g�}`y��A8dO�3��_]YI7��a�LQ���9��J���2�'�Ѯ�J�V�H� �C��C7)j�1B�
Td<�v�NBA��z�r"{��Fəit���	p`��j�*n1+	�6
����t��������g�0[�G��b������i��ơ���g��<p��+9��G�ѳU!��Wm�h4�W�z��l���<�g�M������;1<<��_}-�-�GP^��֯�?̆��Ù��:�a(8��/��n�&���}g�?Zh�X�&Ak[�ȘS"��f����BC���3=�P�/��$>�E�<xܝX�f5�^?B�4����?�2f"�d�� �j�)�`�	̒�r����;�yr�F-�a��W���ۮ^�v�CNo@٠����?~�<��6D"�����u��j��H$c�e�-�af%E�e�{�L*A�ƆT:F�1o[� l�X�Œ���!Q��Ż;��Q�@��	�g"0Z\t2eA��zL�t��d���#�_��՗?����?j���������P�G���(�V�s���|�4)����W��� @4ʚ�zIa���� ��f�W��)d[>,׀415�TU�z�Qs�|A{�GqyT�š��3b=[���~�f��M� >"�&�k���^K|ٲ�v�^k4�=�TB�T��LZ�n%m�����F��腑�5��q8s�mxll���G�oݺu��w��o�k�������7d�����ۛ�rV2ku6��V��^(F�1��y�y^�Ƅg C����K�kr�y��џ�r91���b� ��,�!K����`���x�kbb�����߅�>�b-�����g������g���=��sMw�t�v�U�pt����g����*���14@Py��OCEf����_�Ξ=�W^{]�RjZT�E�Sl�9i]Xy�F<��+x��W&�Q��!W�832�m�?�O��p�F�wPd��<N�4z _F������k��E'?� hbi�<$(��g�ln�L&�g_�sCL�8��`�M7�lk�o�o&�<��u2��w�g�U�z�d��f-&����G�@�C��67�'���U�V.��O��{�V ��X]���;,�6�[���\U�
&�F^y%�Ĉ 3p� F&�%�ZE:Gy�6�A�"`˒���t�3'0o�<x�]H�u�r-�xi����?Ad�R���˾���_��z��>�࿺N�:���l#�٩�M Tb��}G�
؎�3���O�G�Z<:�
�K��l�����h߱�f����h�	��d�:-i�*�߱c�j|x�E-kd��4�X/�5����uh�G��kr{C�\.h��1���cF��k�/v�{��9s���=��c��dt��"�z�H�&:��bA���傣�Y�2�=S���YMUIv8t������������N�g"3�����|�(�x���ȺXA2]S೓!Ցq�&/�ۅp`FD)Q�C��ҩ�14���0��z�;�%2Un��$�=U�șt����/$�å���yl�j��_�����3O���?b�O����o�\s��/�����C���ϟ�tP���'G|��|���v�:�y�<��Yt���3�o6��Q�x2�S��!E�m���g��9�K���e��>L�?���?��>~V�]����9��ɂ�
E��TU�v	���TAw�<�t���DF;��^�Q���O~��qR:�{���GNK�ی\2��y͂3�{:^�����a6�	�f�2�pjʇ��4F�L�|�rA�m��Xg��8�-������羀������/�?}�A���I����%� P����c����ʉi�*9�t�rAt��闵:3�n3�.�/E*6��N�l���!^|���m/`��QH�r�N�ߢ)���C�=�����G�*i��Hs6�m"��f�^s��\����6#�R�X�@�\_�3i
@��ʈ�_id[�?O�/�u���`�P�@��Xb��Y���Lf5g����.wps)b�L*J%JA��W*՜�`om��0�~���uي���=ǒ��H�`�+٬�L�]��Q֐1K!
#DN�J �nv�����A�"1B�r�=2:�n����_~��7n�����<��y=�����r��:O����B�D�E!�*�)�p7{av:)J2��!�r�!��g����Q̟?-�z����:��PmbB'���
 s���/���o�Ex���"������3������oE%��M�/jQ47"��`�-8|�<��?|��p�H?::�@o���=N1��͌)n����f+\�����45c~�2�v;��.3:���=����$=o=���A�3E�\��T��S�2@f�N�΄౹KeD���;o��{�BF�B�,�"@�6�l���=�`l邽��Shj���]����ba�r�~��رg?��4 ��qI� 06������נ�aM�Vu�[���W]�	iO6�=�o�Y��i5�{��y(�b
]�(������#s7���ׄ�@ ��B���nT)�\���Èc����p.�]."������C�o�]��|l��h��z���n|b󥗜��^�Ą=�Pt�Z����ld_s�*�BS!˶8k��Zpp ����d'�B�����K�>J�h��P�m�W>W(��6�V��P���S�D&����L���=��2�12��	VF4v ���-�T�JA�B_���~d���w�9p�Y�+W�E��KQ̞B� ������5$�/DT� �`S[߽��D� B1�V���=��%����6��)1n���~�g�;��J*Q,�M��z �!�ɡW�%!�ÍF,�dv�D6��t�h2!�NA�Ո�a0A �����D�MD
ܼ%R���,�N���TUk�t�>��H7�c�b(-�����L"��T:%���|8�^�YdIo��h����XI:����������C�;�� zBx�%W��iw	#�����s���L��4�����@7l�
��/�sϾ�G~�|�a,�H��>�y�tA��"dQ�g& Z �#c���݈�s�����؄�n�Ͽ����
��O���!�~�:��D����$,L�E�iz���	�̇*��7��9|���ǎ��PYК�(W�0�qn���lX��n+�z�'�&�/_���T�1�	�,^ЅӃ'���@Q�F៚�s���ϊ�����w*�h��5��J��<W"��*�&��ܞ&�����XF����y��=��AR�8y<�-7������>����o��ڳe`�����w;r���"i#�ꍆ)z�G�.w\�*"3�\�ʙ^l'���z��	�l3"_��G}��ސȶcV�3���d���57#~���ԤV���Z���ɤX�Z��~=�T`.�%�\��3�&�5kj�hl�o�����`�����3=���7蕼]Q"Z�-���	�2�}4���3E�M��"z���Te�욘�]v�ԉ�;�m�f���].�2�����cG��Ҡe^:$����H��e�����(�Y�V�7���XL�!�ry1��`!��Z�����l����aVfG�0+��2Ωd�mdr�����GH��,~��T�C�O��oӜ�+7,��TA�k�(�҈���y���Qd$g�r���
�A�D��a�?0��L`f���� ,N7���82�9e̿d	��Ե��<�����/_�'�_�D)���f@F)�sԣ��Y4�MNL��5`���v4ѽ��:�������z�#�q�$z�	ir�XDt��fX�ف�=�PSD_�G=�o~�a$�Ə�S�B��UŲ
FG3��$F&|P��_��}]�[͢P��(a	��-MN��t���=ܓS)q�@#�
r �4g�U�Q��|��5ƽ�G2B�B{��};�9h��f&��7\��#����E���r6��܋��s��/�r��sma`��W^�g|Y%�i4�u�ԋ�Z�?����.��Lu�"~ok%�������>acxB�@��#uvj2��0��7�R�j�Rɚ̖@�������w�^�������0��3�B��R�+|O�ɕ�3�&3[���)j$�p���Es͈�q́���jjBn��KN�9u�(E֋I;*��T�hF���m��x$��IQ��6�.�mmm��O#<�hJ�J���G�Z��{l˖-��qa����s==�>q�L:��Y�fQ�#� ώO�X[�"!��t��b)@��C��42��`T,�k ��v"���)Rt��B�5A��M�*����seV�UɅb���cc1.<^t�Bܤ8X����r�㏾�+{z:t����Q"ɦ�����Չ,9�bI��Ͽ�/m�7��	<�ݿG���H_�FWJ�7z��f���*��jh��p��aǡ�h&��u�)v@"�8D �y_�җ`!�}t�n$8�C���X�z%��G�,!�/(L��w��n��W�CsK;d���F���벢l4!G��/�{��`s�ڵ��	L�P,�����.]ډh"��Lz�tF����~��6��k�f��z)�k����BK@�L����E!�:����˪��t"�S�3�fDfEIB�Rc�˱��d0 �~G�2��\�YgBCs�]Kb��b(	��k�k�N�S�����Gl*�V:]u$ҩ��|�M�@����z�6��A��A�Z�{��Q��ɋD-�3gt�>0 ������c��ߗ.dxR�R�R��0�����s��i��0��&~=i6�%�j2���k��*� <�r9��'��s�
�����hqDV�z�C���=��Hj�&���p8��D��a�8D��N�=G{�H�l�2==�����u߼y�22�@a˖'g���wL��_n(�����ғ㖵z�3@r��(���=��=]���B�@�WQ:(�q�mGcYdL&,6��[�w2ƒ�,�ƻD6��F�#S^���G�I�ìŒT���m��?��+�����U��w�CN�{�VQ�k��"�D���q�����C���M��)�ew�;����Z��Nap�W�	�^�B	�����w�%���"	���u;n�r#9�r�:�v!n5[����Ǎgq��	�%l��۴�X�T�'�o�T @Qz���G���b�,�:؁DI�hOME�8x��Z� V�����s��`�b}_����{á�	U�j!�VW^�	v�);F�V�Z�Ls�
��<��#�d�D5g٘Z�y��	R%�f���4\' ��erB�2RRUW�8>8����tva&���nA� ��d.��3��ǎ�4ڌ�7]���� x��]�Tv=O���d�jA������VAݹ��ujb�<]œM��4>�� ��z#"g���ϓ
*Y6�1`��\
��/�Q�n�^o�������c�&1��0�{}*����h����bnnn_�v�ì9p�;\d��<}��a%��ţf�l�M֩a4X�TRH�ፅ#�64	�"�.0YQ<��t:�.�-GN��q��e,�|�߾��tw����SC�rI�Q�j���c����+�'�(:0I�d�4���&����Hf��'�J�H��V;,��!	�}bD�9D�5�̳��%]4�虞�l��E��/�
\bx�t��?��v[�R���ӵ�u"��@�x9S������1,h��_�2bScx�{�z�����p�݂�H��;���ܵ]�qp`�8��ƈgl.�Ke�	4��O������DR����!`�|I�-Y ٮi�q}�`o�=��H'ǦuV�㇚W��!��|yA���ir���}�-�:r�Z<h�����?�a�V�(�!�3��~n�������H&B�L�!�`�	�Ԧ�q�B^�2�i?qt�dr����`0�tj09=#�U���&��E���Kd��4:Z��$�)�^��z��z/+�V��#{�ކ'֯_����h2]3>_C:�mרuZ�q�Ι�d2.��-by�j��H-k��2g��}��gΜNX��	%W�*�4ÅkhĴ����(o�bD2�NLݨ�`
}�[R���}�y�޽���y�*5ʲA�A����i3O�B6�{���Z���6Q�f����6ό�f�X0G~�>k�#ՙ�����G_Ng�c�xo1��XMN��K�Ҧ�4##�pz\�W�j֑1mC(�#�b��25[�{��+��Γ�?��O]h�����m���ָ/��u�&��/K*�b,�Ќ�˕<re�g��q���L�|��V�]��H�J�P��w����l�a�&s��9���u޹<BF]��	�k5�R�ub|�yjj���G�J���<�wZ�}��?y�|&8q����5S-��YVZԡL�k��%��?�2<r��t|�/��?�����'�id��8WK��*-J��F85<��5W�{��;���wӳ #�4)V�4A�&�6p'����dC������6n�a�y91�	r�i	�)n<c�D�.$��ΐ����X,2scb�z���聓����X���ڀ��v�� �{01:����4�HĦň���4�CB��`d2%r��H�@��pZ���4�����$�,�����W����N�"W�vi�r3��ާ�6x�͂�d��IVW+�J�ر�o���ww/�O�࢙�y��L�����Jn�5z�<�A�U[��j�xչ��s�
��^1�@��f�/,�V{�)5��%��i�T&Q��2
=c�-�A��N���;��fkq�ɠ�ӳ�g��e��Y9r�
fx�*�d�'2%����֡���9%��Ys��w���k�<4<2����l��dl<v#�ِYb��t+�k'&Ǡ3��6PĮCs[�@�c㪬��>s��uKO��u��ÿJ��5YR���w���}��֚�&�6G�\����"�=�3�8r�$�8z���Ņtn*[�k���`|�Lb�"L,Tó�*���(���ɸrC#�r1�wFC���䤓ni�O1$��'�~����ăVwKK�,sI�����n������������h�#-��Xv%Y��V������/��P�l7]{5V�^���v�W�lē/�����9E��ңq��>����>v�*e_{�h�\����C4�}���Ĩ�����>PECش�:\�z���&��m�D�P��i�H3�<Do�<r$9�y���c�ؕ�bå����E.������?��AԳe1�I��3�'r��'7رT���Q,dɷk���c�Z#��݅:97*��F4:<�9=�:hې�(�T�J��N�Z������z���*�����1W2�Z�N+��v�D�H8nN�s!�����?��M�Wx��P�/H��B����#gu�p��Z*�4���U��Bp.��n���l�1�>P��������hy�TZ���-��X�j-���~�hk@D�\ӫ�R�IW鵳z�~����1MQ��k��ҥk"�{)�ɮ�C�X��e����������hhl��&q�(�A,Ì�O�bE�����wӽ=�|u��Ɍ(ݽ��9|�o�V���E���F�g~+U��,���x�F�n������K��O�He�$[9��7	�1۽̅~u��N�N��LO4����D� ��Z�|��mO<��f"�ˠ6t�t9����|#��X��E���4�-��������x|4�/�����_���?�D|w|�ftw6�_<���L�:��+�#AQ�ַ"_���bF$��J���܃���m?:?������~]��U�(s��w�ь�
���u���MP�y�x�yGaq8�f�)�{���9�y���,��Coo/�<Pq�,�a��,v<���Eq
J&�l*-"N���A]���Zx?��Kg�5*_��T/t�3 �n��pV�N7k�J�5Oc#�ѦϜ;�V0�ފ+����]T��UO=9OVI���*��}�P~���s"�/d�UbYd�}n&pp���]�,���$��>�qG=E�&���?+�v"�.�*u�iw�y�I_��~��S�H���쐤�i�~L�R+�
~	6��^�(F��vk8�>m�n�+)|�5~��Yʾ�扣��{lG+4g6���tഌvKQ3���4��/8<2ɔp�Vr�ұ1�  ��IDATg�}����C�'�ti1TkL|d���{���ck3��Y��5<}��h&&�qwoUbD�o
o�t��&�Y�2�$�w�"���� ����G�0X-���k�m̡�EU�ե2�����&����F�k1Q�`�zFg0>��S�UGB�{T6GgQ�J����i�x[������=��;�z�p`�.��g���X��
�{l C�Ӹu�ͰPd�¶�x��{�r�J���Yl��R����t�̌Nr�X����s)����W����/�x�ŗp|�<*"y?�n����}ظj)2*� �z�Z�lw��(�C�p��Hs�H�8�
�P�(}���X�b	�N� 9RE`d��FT�"�e�lN8���ħ�kڙ�`?�� ������W&���v]��x�Ke�a� �������*3e/9/������g�F�(y�����.s$YI�v�a1�PoR�gPg>���B%]�P�lb�����L���S
���T;d@WSz��U�w<�.�4�q��5ɲ��w��m��G���,4�MN<�PEi��)/�88a�6���d���Ȃ���tccù>��#=���ḱ���Z�h�����;�ĥ�BђW��P��G��W��F"!LOM���&��ys:/K�7�7h��B���Gonln!P0D��3�3���C�Nf�I��������4_.����5��!8��6��dFLh�(JS�䈎�8e'�/P)����5�̆[�C��}"ԅ|�qrzb���җ�[b������ǟ�������&&�MT�ض�6�z#^?;��م��Z�����)N>��7\��{�b�у���k��ra�K���u���S����� *7T� ��i�K�2����"�<�Q4���]hp8p�'�B�t�%8=z�����۸��p%FN@IDp��WѶp���>�]��Ǝ��AU��-��f+.�l#F�(%HܶZfv�
��I�os#k��7��^��A�R��,}���jxw��>�5S��[-�ck5�`�/�n9n�-N�T윜�g�屩�?|�T�<�jժ�t�.F`��dښ�d{�l���Z�)~L��ɦ��ag�#��Ě6A�=���E�p3��dο65PN�*��B0���,�đ~*��R��5Y��v�g潔f���;zb1��^
`�h$�\��tN/d�D�b1q3"�ʨ��}��xod�z����f&��h{�>̚����岍kO�>sf:�����t*&R�ܱ�Z0�qd��D�:�$�-V467#�#�W���,c>�e'O�|ݕ~�:�o}��_�ű�oþ)��r���J]&��I��42ǔD��`�9)d�%d
�������H���̃�4+�D��k�2�b�$f-�X���J�r��%�H.��Fl�7)@8�@�'���������MM�D6�fB���%�uh��z�$�����c?yG��7nB��C/��/}����>z�8��vx:��j�
<���(��7kL(���⚀'7�p�����8�/]&X�v�|w�}l^7�$N���dD���Ko��Y}M�q���ѵf=����;���3"=���&�s�R�UCM��+NZ-;��`kTr�Y�Y�F���s�>��P���0��gy��Y5S�,�^�AY�� {Y.'6r^��RUc�t��W_�9�������z������;���߯y�W;��R�,��<���f����U���sJ���
���b��ǫ��8�����^B��RwdWc�
�1�x�R,T�V���t�>P�l`�|����1�:�I��i�ehO�^P
y��%�����j3צ&(hQrQn ��=~���3����8�=-���|Չ�˖��O9�"�M�dQ&�a62�j����}Le��l��h"�(?����l�������{�oݲ���[�.���l��Yط7�Ig3����0l�S䦣���i����2�6x�[�v9ŁO�H��Lg��M65�d�͜���,X��Κ���,�R��T�sr���ܺ�f�Θ��}�OgO��<�l�lHi�l�*y�Fpj
n�9����ޓh�Z�OG�p�
�yߝxm��q��wd��^ďVѱ|�-Z��~�*�GDު%�b�kjb�1tr���B�J �ׂ-��h/axr_��g1��c�3�)�L#BN�[�����+q��
2���f���.���j��<���æ�E����g��]����aD��yYE{D]A�%��Y��\*�&\�J��޻�! �=π����h2o��W��/WY`IK��7Z]Bo�b�V��G�Oo�Ş��槯��w=�E3�����Ȉ1�L�ӝ��U,ύ��Pt��S��2˒(1�x�_�荂 5�!�oR#"�\���G]29��ɁDY��'�.�Y����h�y�e�@�R��l�j��JÄnEA����X����k��Fje��VD�5'3L�dk{��U�V�0�>К���كK7n84t~dG&��(�XX�sČ|՜�Ss��B޴вohl��P3f�J�R,4c������c�,���֭[�9U�R���3�'����KJm�\�d&��i�B���>;u�g�S��%����su*�L�@Dd*8�12�%������r:Q�V����";U^��[f��%���g/^|���Z�)�|����O��O�=-�<SH�%��3DI����&�*�����E#x�� :�[����X�v#�����O=�C�G��݅[n���=b�|�э��>�L�����s���x���/���r��+�! �W�_��?�3�Z�O<�<6T^|c'�� �Y����n��ϡ�g1�����w��/��=����+��K�P�u�C���hj+��缯Q�U�dQt��.EF^�(UK"�ōe\�{��2��b�$,�I�5e1�`uz�nh��^�3(�*���c���>�jKk��{���t��A.+��>�Ng2K�Œ���J�&�\��H��^�O*p �.�0 `�@��2��^{����h���FѦ(��Ne3Y���}�k7����|��\N����9��ko��d�F����	�֩5i�=3`��{�{"h��@CC�o��胯9p�{\�ONVC˗/ߓJ�WǢa�Uz��$��Ü����>���h��fw��t�6;fȡgSF9��z��n~缓�)����#�E{�w&��an��zc^.R$)��/�[����A0���i#�a���M�#(���œ�19S������I���ϖDR�LIN���%۔Ͽ"8|�J�]��hMʟ~�ɿ{zkv 0���3_�q��tz�e54f#R�tU#���l��%�qx�=3���ڈ�v���S���܂�7��݄�~�C�d�[7c�Cw�ǟ�5�]�L܇��q��˰�.r�V,]��<�s�a�������_��8��d���pbhL�b�^<Z2�,�4z��{�O݃@$�]o����zqɒ^���q5jj�<m�Y�2�2�uY���B�V�.��"91���#S%�uZQ��^��$�y��D�������H_7�!Iryj�}����i��x������J��۱c�nrr�/������В�5UQr�)!>U�x�,@�9G�bz�X��g�7�fC��p!�P�Ff[��Qb����4*�qw�X�降5ڭ�2�tlx�����U
��|eV[�=Q�I�Y�%$l3Y�{��tϜ餿�L��]��˖�̩0~�5~ϫ���V<���v�UJŶBN�d*�͌��"���#�"�	IT��1�1�0�G�\Х��ǎ���vOnٲ�H�9q������ht�V�t�t!�u�2\U-�[d�f:�|�y�yr|B��02g�bM|/�hf2Ԣ
.+08�d}q�xE%�j�����}�z�E88����%�Jc�g�������3�O�6u��J���sUbAN�ڠ��1���=�p��x�����ILLN��=���N8,f|�S��@F�o��u��vXqh�;p���o|�1I��q��ص�m\{�8<x#�����0I C`���oA<����/�?���	���N�����ى��B	�O��ی����֛���.	�O&T�s�a>-D�8�̲�:5ϣ��gԋ�D���1��t�.UU���c��\ږ��F��<8��q�L� F�6t��z��7tvw?��͟���P���݉D��θ�M��=�k)�fyx���#��Y\c�3�C֨U����w�Ur���:�U3�4b�x�T�L;�����}��.�/��ݙ���l���-���lT:������V��`��;S�z*6��L��e`ٲes#�b́����kά~+0�_�t{�~�./�*"�Z���f���	T�%#�u��"'�J&f݅|�6p���-�'�-_3D�����$/^����^��f��ds9� $A�[.U.�3>���F�IЎ攂 �H�"�4c�0�����D(�UTr��\�(�$�����E���Q`�����l�����ޭ������s��1���D�(E�Z�h&����ю�SQ$�~T6��p��1FX��/���8��v��[�����8޿��]�d�&�6�P���x��K����x��ǰz�Ft�wa�����/a||���	��&t5,�e+aǋ�S�hD��Ũ�XM�f��"& �ƥ+!�|�V]EJ�@,�_���=GN� ���T���E3�D���P�p�!��˂�Jeޯh��	8\A���8Y�+�R�!��g6m��MgO�q�kpI�?��7�H�����v�q��\&�$��8�u��Q�G�� �������x�ω��h�\+-�sb@`�`t<vJ ���Ȏ$I5�mn9��o=�߲�ӿ�w����p���tB����.�\��E_���Ą�٢�N�hf�%1.I�G�2m2�u/똾عV>� �6mah(u���c{'''�S�b^��UYH��� ��~Qǳ����"���4 �r�VVr����7�vt����}�O��O�-[����7��9oc�A%�YBک�U�V2���P�W�Ղь�qّ8�~��"��X�W��T"&�4��T٨g�)1�\)�Ƃ$<G�B$�]����2_������]<�MF|8����@���S��M:�U���ŀ��ӸZ��^�CUD")<���б*!�m�?���!|�(�W��L����_�E���Bgo/��:о�tG���с��.��'��M��c�"0>!��>�8V-]���lD5���V�����2�F���a^W;�'G��)p7x�q�?ҴG
y��X���H����
���-;���Oo�#T"/��f`P��"V��,(�-������H4~.�+�����Y��5z��(�����}S��Bq�wFsGģqQ6`�z�G�b,�Z�ЌX�T�����g�I�C����#��̆Zo@*��/���l<��l�~g�����?x���*q0Saif�`A�"�;&�2YL�{Ed;r^R<��*Z�&��d�jh�`n}�5�@VO�9|ŕW>�m���6�ݞ�)�����z��	,�%$�$a�E7wsc�PS�l��L��+��<��jÚ�w�����O)o6oɮ\��W^~�*��n��Z59p�S�����xM=8��̩�5�"E�|ii�=-(�q�h��zcmT�5ԪMp�Y�"����xt��?�&��C�~1@�VG��^��ȞC�K�r�٠��޲|lZp	��� ��V�T�	<��;a�}rzdk�.���3�%E�,l'O���U+15t�xN����Dsg���J���[�_�*+h!<>���w7������y-�|��xu�Sh4�p��BU* d/�CN=s-�� �1�H�}{S���e�ș)5��)��E9e�IQ���c2�R��c 3�J(WJ��s����:��������q)�HJ���hr>ks������u9)���N�+mF�Q���<�"z@��FE!Įp� �/
�u��}<9U�5g]h&��~}j�j5���ΜEޒ�x��n�z�u:��N������-ש��2[��J�{c���aSuV�(�Cyզ��B��ht�����V���I�>� �>�x���g�;��`4�(ٴ,W%֚��W�F5	#�Z��Rhu�T���I��ɘ��i�Ǐ�_�q���-ݶe�_$�,�4���o&���jY�h5�T!�JΆz�X�M�3�Aq�� �I�h��tt}pVC����եX�Z=Jd��Y��̸߀1@�,q�&��vMO�-���,3=�=�+G~3�Td�,W��jIUL��F��wʆv�K#WTH%s�
E���B�ΡScݚ%��C��8}nS�b�o�ʕb����+hkkò��� �yw�� n�|���ٺf�	*2����cO"�I`eo7��6;��+6�[M���`( ��$w��,�S�h���`��n8�$;��DQ�$�F�JU���<^���0Yd)

�2��R^��2��oa a&``�: i�,�S��b��a�K�yϑ��q����¿|���x"��>u9��;�1�o���\�����3�Y�E~�������^$�8�2�Q�`�m��M�ߩ��7U+U�G�f�Ȗ-w���﵍��_J��A&D�eulTk���l���,�e=��U�l&�T���RGW/_�H>��@�i�_�yj �I�ߙͤ��\��y��.:g��75-�^*�hN�44
Ω�b6)��l;y����)�޴��F|>��,��}{v-��W늲Q��KLQ�5���0�%��r3E�QiF�d,�8�4>Vo4jL����<G��,c]�Bsݻ(-���Ο��d��9p�ֹ��gx·� �ZY�l�X��o4i��sٞ�I$��fɑ��$�W����/?�����ޝoC�*�c�_=��_~	�D��0�ۊ��;' �$�(k���g�w�^x�y|�ڤ�C/��݋��@Q��\��3)j㚵���R��2�a�6Y��#J^ZrJ"!Z�d�RK�<R�T�ALb�.��%GS����!Kjq�:��媷�c�F.cqO��j�F��JZ���F�O���s��߮m۶�F�G���\D���L����2�x��z
�}�F����3�u�Y�`��� /(���;r��I������h���d2:��dk�7�~�|��˞wv^N��g0��D6���P�#Z�а1P�q/�<��b�̑�lW׼�ޫV�M)�k���K�N�-]�R`z���r���z�T��1����FdK�G6�h�u�i�Aii"I�C)�,6�����3�Nݴf�z(�=�ic���΍45��_X��:�jU�/�`b��QH���Y�$ H>u<2�
�1�T��X��D�o���`d_��t.jөh�IE)��������L�K�����^�ժ��~���T6�ؤ3F�5�޺�c_k�U����&z0��Ƙ�'�V�X�l�դƑ�'q��Q<F�����S"b*�I��ΟE�%�W_}��t+*��O����聗"�y=}䜁뮿��}��w����uY��W]�R.+��fr��������I�F2�LMM�A��j�|�Z������TX�ZOѩ"�^��4��>`�QIP꬈��'2,v
�j�T�d���v������Cf��{.Cx&ܫ�XhI�e��BW���� �S.4"��r�����dSlg���uev����Jd
�se��F�Y�5�D�H�S�c%%��]΃�����	���x���١�tZs��ёY�BoЈ�&�lZYO ����6�1W΢%3�
��4��Ǘ/_~~�E,��é�?�ţ��]��t�̛��Z��������F��J.��ቱQ��2\.��}������w��QI��,�N^�3�����%�%I�Y:���7:O=S�B�ĽX��h� H#K @?�x���'s�BaA��d�0�l���ͰYPҙ��k�BF��7���U"��O)���#绮>~��ԹF��X�ь���3��lZ�Ӣ?tӦ�,�i�'㦜Ƽ3�ɮ���n��D�A�@:���MH�:1�a��д���w!09�}�p���X�~��(�y��~'� �Μ�'�r����%r�Z|�3��_� "�ͷ݌}ߡ���Kנ��"O��a0��5He�z��eVMlnpC+�n�$�'�/2�l����1�N:�~�y���H;�3R�}泂����*&-�i���ݍ�;=,,�REJ*��a���^o}��4�� �{��O��_��WOw�́���{2E*��B�G��C-�[��r�l@F�8%�\sF���:Kl˵��$p����ieF T���L0��R�*�jmh����^��~�����BeqSS����ɤ̇̚-T#	s@��r¤ӊ����o8���-Ij�xSKˉK.Y0���[�9p��fGC�W\��盾���EK�P��t�|Y����tX
�I4�6�����E��>E��4TQR�D:�t����:��5}2�f�h׼�ώ-�TJ=�j�f#�Uk/��N����B�Py��C$�N��F'��z��WE��Qa�R�ϲV%:�E�5!�����1́��Xg>g���jQ�5o����=��!�(!��l>�1e��gs�F�E���V� j�-���>�J�8pF�wݲ	����8;�b�����$fؽ�]��`�=��=�@XL�����(�]�{v��I��+/AU�3��;�M���&m���a�L ��x,,<���\�΀y58��h/���&7��*���,�T�Do�8���Z�D��m4Z�1�(`VG��P)GQ��5MOZ��]t?�9`�ދk�����r���T��V�H�gq�l�j,�����J:�,�l��Ch%��"�%TjY!�U.�8��̅��K�J�L6d�9�ں:���~y�g�Ξ_�Q�ڌ�̽:�v���@�\cC4��v:P*V��'�N5�(Y�����]��\�)0��k�.����}�P,u&���xDSb�zB�:�����N�t~�e�	VW<B�L��N"�W��V�c��'O}~~w���-2�]���}3���iЪv�yr:�n6e(��(^h2�
���0;�&�6X�fe�$2:1I-Dt
�6�ј�U&�x��K�|�z���A����7_���I�Rk�k��4$滤<}�x���OO�`E��TcA�T�24:2���QPcE���3� K����>��O����?�idb	$L�dlUF#^۹�s#��S���7w㡇 �^�):[�t9Lb�$����-*(�3����3g�x�FDr8w��TW�p�9�	�^=]�"�d���Zt���!�[g�+�j��*��f6O�v���JzMo0?jW��Hfi���֣�>o�f��&:�~���qI�ވ�ٝ: ���A�u�ӳfgϣ�\6Ш~�/��?��g�p?�M0��:q�H$Rù��;�5�3����~O�8e:v��eS>�:��a�~�:��esyd�<z��G<F��<Q��Xf�Jve�j��۷�wb�1��_s��tuu9�W^}ݎ)_`i2�l)�r��xR2he!K[(�!����ES"���W@Q��
�ˎtl"�j����ў<�g�9>�����ar����k�kW��j-�-hE�,�l0����I�d�}Η�cLf<O�/���q/�����&��$B���z߻����[w�s~U�/I#�{x�i�]]u����޳�oK�4����N̙ٹ�����JY]�̝ZY��(�1X�����J���r����a6��\�`�T/Sjt�^������t�cќ�Ba�D,6��� `�����x����ܲ�����ER�H:t�b�FZ=nJ�L^(r�wS�X)&_�,/��Rv�{o6�q/\�f-}w��@��λ������oC��6�s/�r%ضc'd
e����Ѓ�b�*D,&���B����=��j��"�{x��xX��qhm�1u��^ ~�|!�VʈĈz��0"	rjU�x0���p�^b��Z"t��/��\?�Ta��W}.��=�P/���NJ.�2�i(����G�Q�2{��ja�\�+[��Y���/���:%$��YmC��'5�#J蹵V�	�x���
9���~K���k_����c���k%p��[�O�>���t���Zb���*�� n�"�Ц��D B Bx=�ӧ��]k�,�
f����1�ˊ/9s��|���R*�J���J���'igѹ�N�&�����c�~�͘!si6F��/+b��`���}���.I<8kVG_"1rftbl�S�zi5���J�V���0�jt�%D�|���5���u���P<q�����Q�I
@�T*����f��w�s`�%���+���l��4dS���*���̠t��Qs��U4(㿹Wr������U7�tJ����?
U�/��6Z���;������]{@�x�b6?�ʫ����A?���A��A������Ͼ ��~x�>�&�I�>�f�$|d) 	8:x�8
����U���-֖�T�jx��ߺ$��!��GbBbD4j�5����p��^���3��g9��i���C�a`ۿk{��_y��.�]�,D.E�999^'5+�$�8�U̑ϓ��7~'�k��L��s�\6��'fJ���E�"L4hp�^,ƚ��ε��L�{����u�����Dre ��%�#�zL���4�L:��>�+1��&C�s�/_oW~%���G�:03��92<2�R�T�BT<����,G�b| ��$�f;�^4F�P��2�X,���`�'�Y�r���tC?9s欞T&���^"�����1~�jUfH�1�I�%*U�S&�� ܴg����LA�&k�������������������0
��G�1~��!���3�H͟H�[1��I(�YE��6�bA�9ك�g9�004�4M����d@�.���x\�	w�~�5~���;w.���a$�'����P['�5��;�σ���n��ӛ`���L9�(��x6����aU/BS$
�|ښ[`Ŋ��inne����b6i�v1�-�X�X�`�9:�ɆX	�����h�[|xL��U�{�-60���p�p ��-��D/L�,%LH�����F::�ozU�m�L�L=�l��@�5U�*
�$�y�;�PE�Z�M��^�9���֛��<y��:|����2��4z��a�q��1!�]��b��w��O����l��M�����#n���֯[�'�ͬӴjTS� 	$i�A���cU�)&��pM��~mlC��
��E*74<��ֺ�1�U��p8��>}F�|�Y�� �:#�ᢩ�bga����^fՃl&�l��9
�S������TUY�ț\�:_;f1n�"z���1��ؓ����ܬi�'��^;��\�޹�g��Y�:��q	�,Z��}�"�����UL��?~�#V���B-ˁ?f�T]*	���Y��{@BD�l�*�8< ��y+�hW����y���j��O��{����	h�!�Ia�Y�����N��t�~�F8{�,~���5�?��L�XjUc32�} &S�`�	/�Z�M�;�^p���6C8ڊ�[j�,X<�_���<j���9۲e�p���6Kx�Q5� ��=�
�~X��#�$�TRd��G<S��z�u�"���*Slhhh`�L�=�N'	��\.���Owv��<���_���ر���s���f�W���s��X�uҀd���}�ɏ�ǀ�jkP��Z
&X�@�`ٲŃ,��_�lp�7�{,k�����K&s�^߂��4,$�:����ʹ4�K��x�� :�!6D#J0`P���8�X���>_���Z���3���~�"��D`}j�"Pɑ��b� G%�fz/Rt,���PS!�"x�$�
�O�*u=�:Q�""�Q,����\�p�0���O�|��Ev�;�&[RV�;���.�K��ӎ���?'rE������2^�m'zB/�����Iٝ��)����င��K{��	�'���;Ol~�x@K!���/�d�sĂ���,���-/�W�h(f�M���J2��h���QNgg':ܷoI��~"*��&W�!� 8����ج�^g�{�2?�[v�Y���ˋY��i%�z�p?� 5��\	l�Ϛ+]L/�l�v�Jұ�"��E&h�6��߶C� "��:t��OU	8F�<ŊXKP�9�������%��RU�����'���7���r-�I��v��dFH�ժ�/��Lp�{Ȳ��8�ڲ�'>Gs8䡆��+W.�I�l�����q��c��gYᾞR�(;�fbYb�99.MN���R�0&���f���a�J��L<��3gN	+W������xX�x1�>}
ʥ���W:U�.tH<p�,�� ���Uё���"ԓt{jBĎV�C4�L�@Z��� Nӌ�������0<<bY�3���m~�OGs��������k�E��E��U�~3S3#��gpp�J�˜)�� �aV\ω�`q8����;o����'a��{h���`�2~VT�
p��0(�sC�.�gN����0|�s���7
�!X#��p��;*fx�x�MV��=�����c#�����	���T+&>��Qhn�&f�*�L:w$��B���2�/a���\&������6��)�*S-A�_�:\e�4<:ExD�kdTi����ź�� pu�$���ц
���?��d<a�&Y��8>m��ӏ=��/\)�޳���o~o}��\��y4�L�';D�j�%�#N ��a�`��g��Yھ)�-�{�B���ŋ�������cbK�Fbo���m/�G#w��g�4v *f�&Q����k6c��3v���$�\��Fc$S�>{��b�RPTvSûx!ɪ��N�K�*�����~M0W�u
�V���P�X;� [}��4Rr�C��X	�J߆Uu������i���+��W���_��o�x��b�܊b�{�Y�w���� ���Id��)s�3�S���D��\��&V���b�U���2�B��!�`������d� +������>0d��,�I��̚��pȜȪ?�D�Υ!�L@��L2�2E��9W���8�8q�Ɂ�v���႖��
�ө�x?(�=n�ё���*'X�\a�����x1{�~�2F%�C{��/��ٖBmYaC�$�Ĉ����
3�SbF�S%`��?U5��P���t.#Q6kD��n��{L�&�uL|��pS������/�VbC����W݅/��t�yں�;U�À!��#�3��"�B+���@���q��h������>&F텑�����K����4U�&/{D�p1�iOÉ�y�qpx���Y{���J�<�D��c�W�@O_?xhii#���ӹ,$?t�K��ќ4�����L�[*����E�T*4�.�l�L���Z��B�
-�=��O�>}9�}��76�X�wՑ;u�boO_���d�I�jN�׬H�W@Hyxk��������������l����S\��ik����x�|$�Y<ԝ.���_�v�y���<�(��Sd�6�` E�3<�_n|HPȕ ����u"U:�}�� hs�4�j3`���np�3On�r�R8��~��%(�=����I�醦�v�{A�J��.�~}�M����KZv$뛈�i��L��+R���Q�SU�0eé� qЁ��U��S!��!. r{�/�L?�g� ��Xb@��ā���#���x9�`ޕ'�PKe���C���uC<�X�py�DlD����:��G���e��~/�v��j��gj���x���e��׬Yc�}Hf������׮;�?8�fE�v`�>G-�EQ@tO�S�� �]*9��!h@.F#�Uj� ��V�?�;��4�TG�ws�́Ç��+�Ź�>;eĹO�����|����g ��B0 �����*L�DC�g���e��}��Df��ac�ز��緁~���2�c�,�j��H��X|�)]��9��|�J��HD=|��k�r��_�����M+����|��X���PK���@��wP����{��z2cÓp��+����&��H�4Q�` ��ðe�N��W�����a476A��\:.���c��tu͘ɪK�x���=G�8�f�e����`�bE�fs;��Q	.�Uϝ?}~xtrW���BvU�1Z_<���R>��6��6O����r?�}�&�J��V����:#~�>;�Ι�B}��U�DD�&���N��=Ϗ	�l����#Ŝ����l.��ؼw֬���/���Z�o��g�ŋֺ��f/�l��#U����J:蚦b��!����J���^�W|�[}�C4|��N�_7x��Tf6���5�11\�	�2�@��?�#�vcF'����(���U�2���3p��iX�x	s~b8���=A� N�'H��%ȗvՉ+��;�.j�*�J�t:X�A�B��V��Z`H�	�Z�Vue2�����y���7c����Q��P�4����[��.�:���@����QA��˵���߅'~Ѝ�9� S%���./@5��h?L��Ц�`x��(��L՟r�3e�0߱����,������t�D�C�E0f�������ZU�|��1��x�mj�
��Z;�I��?.z�X�Od��x�'���I�~Ys$Ro��<ES硟9���8�m���d��xUM
˪���B&h�Ǝ*����g	ގ>��Z�]���!���sL�>�t:�h�޻���G+���;DJ��O������*maKs�ˍ@�$�YA�Ș�Z���$���mN�C�<$�qĜf�!9�/Y���5s��j�����cfD:>n������B��,�969)sB�U�ڨ�F�u�?NDE^���s�
����f�����ܹW�ـ��vH�2��f��� A*m4�D����&��U�(*�y��b<Ԇ%)�2�1���@�9VݰL]�m�CC��Ǖ��f�����@��?c!HӲr[�<r��%&~���㱛
�������,���翃o��^y%�����7��n��Y���z�jC��C3�pc3SG<12��'a�.@l	z�ķ�l�*:�4��U����.%K���p��h>���B����$����R���d�C�N�~y�uk_�;w���Kۅԅ&̶�k����Hl �>K@����S�Df���O�K�0�K�*��5��8�V�k�lӬ�~<��ѓ�t"���
~�㿨jpj�N��]�]�_�p:�$�&`�]N��Qe�K�]�Ωag��bt�T)� z{��.X6V��>$�����Z[��c=����сڪ�>��Uy:쩴O�� � �#sY���0ȷ0k�6#8���^,�A���� �aaV��@^:K�
F�f��!rm8�K_�2��Cd������(:� Q� S�|M�������u7c�����X(T���nt��s�rz,{�%9��ep��n\n8u�<�&�`��O��U�  ���7����O_Kv�U���@�J޽p3?�A�<xo�aB�e:������9���OC&�b��i���.lܸx<���;��&��������s�6/]��y<TΓ���Kq;pj�e��Q 0���b0�o��c��P@Wu(�Xј
U�a��dk�|��O����E�dbGnFx�����*DzT(��������"0���H4�����������q\�w���(3�j2��J%�`��$3�E��}/�O雅�J���|��C�\3�^s���S[�lv⥗�=�����.<h#�P<i.�L9��}>$��Q{�࢕��B�2f(i2h�:cw�YX�p1�
�>�z�z�h���*U 08$�I���J��|��2x}8<nƝ�u;Y	�T.@٨����3/0�C6�TLg:��;>:�<y!9�Z�j��s��#G����}���'����}�v��R�m*�������[���k b�?w����:x�NXw�Z�<�~����@����	E�4_�{V���+���Hetft���D����߂뮻>��G�t|Ũ���%K����($�1V9 @��=JbJc�����g׬Y�y���$��,�bD�*_��l����$R1����R����#��|YU��,��@4�^���lmU��@6u�&����Y�A@��Z4ѿ��&(��Bi��mګ�f���E�IC�Om��-UúJ�>���9���2mP��{��f�=H̉��t1�xR�B5�\h�D�-^�6fo<}�f�����y�u��ɱ����?��/_]�OU'2��Y�~&;yP+E%Ȧ�P��w��[�\ɂ�)�1`��������=�	C�!�J3Bs����r�D�V��I���K�
bt�&��H�2�r Ql$�Î(�'
|�\n\0;����h}��bŊ�q�ė���-�w��N���֛�B�,q�}�/@ULx��Wছ׳� CL��3�u7��Y��7@�h8<�K1�/��/��sp��٘Q��38c�q�͂k6�	9��X-����� ?�H4��1Y�~�%f:�}a����#0����b���Ry&�A��+��4���M�����#)�(@�#�%�� ���v�h(Ѭ�LU��'�5�L2�'
�����>ƃB�`#cc�/�L�\0y�����N͘�����n<vpѹ�����h�~����ID��3k:	ĞI�� i�����d6���%:|	$��EsϭY�n�$/����clD%{��������ڨT�+2��l��i|@�́����%	$�fdh�C��������J
��ip������tBkk3�R�$��M�� JN�kbJiD�L���2%?Z7��L>�fj2�:���.�:TUU����d����g]���l��V�r��q�=ǭ7�B�und��^����+�?���da"������	�!7�	�|�a�ޏ����1��}�U��/d�o���,�~�28����_��?��j!-���<�8vOP����������ϟ9�M�Ŏ��[�̙A�l�/q�ضg����8�s���\2�$�cP�^=�z�D��P����t�)�պ��V �H��� @������L��\���39]U���3g�5�c^�}���sA�Q4Z�|c睆eu!q�x����V�k��ȚLtmqJӁ��@YQT_ p����^�vŤ�P\�������iI���O�����;��C�7mFU��<DB>�z'�>j�;�΂3���pKC������)0<1�B��il�Mì��/��ar�>GR���l�(K
nj�!~�kJΚ 	���L�\b���0�2
u��8S�ʓ��{��g'�\8
68�,Fs*=)�З���Ϳ��o�G��k_���*���%xy������m7o��o���8	?z�YXy�F��_�����'x���4�a�ϳ��l���*�:��FI���} �4�s  Plp� >T �G�Ӧ�*d��!"���wr|b�7nxb�¹ݶf¯f}�'���ZUU��pXhmme�A�⊦�FdG��TV��Psc����TĘ!��2��<�Y;s� ��6Q�nb��c�/�09��X�Jery^��^�b�Um�����۶���ԋ���6�C�F��'����s]�S�$�6�<Nk_Ѓ~N����	��v��^�5W��`�!^>���������׾����f��4�<88�$W�^1��_C�S���i2����c��h#�>(e�-I�>gd|�M/Ϝ="0������!���VF��`�K����Ě�B ;E��4�Hzj]k�MES&���*JI� �<1:6�/��Ē�?�<��B
���O����������ܱ�u'&���9�g�'V.��砫�������'�'���Cl����^��D(��FC3�� Q2*8��x�(&���;���?	C�(�L�ÇK)���F٦q��&�'^��S��kWW�~E������-04e� ������iH�2m�1(�+U6HL��"Ɔ��hkkʻ�����SʫtP3ĺ`�6S]Dߗ��%3���bI5T�^�t����Ρ����
,Q;�w����C��}���-�	mQ�Mi;�Wz?�d���uA(�[0~����ֶ�w?�ٻ�?�]&���o�Q96����ǟ���[�htm!�sQ)��CZ�u$��S�i�$�j��Ⴆ��NC2��`)
��P��H�(!�DjM�z��Șq�j#�!566�ﹽ�n���UtB�T�F�&���c�J��R)y�����V]w��Ճ�b��k�x�:�������_�pq嫻v��i�{7�+��A�����{�Uˮ�e��7��]س}3���w����7!�Y��rܽ�> ���AQW =���'��ff��:�Ag:�-Њ��çN���=w���k�E{+�W���T8>_�(�t��'��Ȕ�:S`,��*f?'�sҴ������T<���h��M��,�i�0�O���H���"�K���i��T'���UˮޫL���U%�L��曟.U*+�a7�:[\�gU|S����h�"n�@(��A��A��������/�Z�條D\^���o�56rŁ��ޡ��Ȁ �С���i{��(cp�y��'�B6�����G��c���D��/���9s.\�h���bA�(R� l$�c�U5��R���8���[�d;���i
��["@IF0��7�7g��q����fKC\�B�:����Fe�S��7�f�����o���F��G��N�]��?�C��?.9 �]o;�	:�u�(D��A�Hl,K�FܨB
�!��?��Am��ç����Ͽ��K�g�����W�-[��3G��_��W���g5sS+DxF��)�u�2�?u(�v�����G��*c7���5DR>��)N�t�0I 7��B��ܙe����.N<��c?s`��������h����`���vq��B�Ez/��P��r9����Ḥ9::��cf]N׻]s����l���l68�-��Ӄ�O�y��������<1��rAC$�#��~B�=69f�!��I��H��4LE�x:���0��`$���Y��<xDа!��#��CA@D��l:�M=S��鼫�J���dj�$C�y��YO�����s��\v�ヴ>�c�}�a�����Ǐ�Z�7�M�׾�U�0-x����}�{���L������m���o�� ��7�y�L���6 
��E��<������DK?��b&��r��~��~��+&���h061�Fմ.�Rks[5fe�& ��\���"��N𠿓�ފH��"��@UE����!( �E�`&˦3���T
_R��5��5K��x䑟U^����{޾���6���F���:�0��}	0��E����J��b>�677�kooݽv�u����7�������E�WQ�[K�B�n�\�PX��%�9=����"�xp{�Ah�6�Û�Ĵ�N"9f�<8J B�¹��i�,#!+�
D�T*�j�-���q�{�����;e-D�B�֢��LǝL$�9}f�����6��e5*����z���o���������?~����(X�	[��W�d�+�̂J�kV^Oo�3V\�X�O���a�8��o��ъ+�Y���j.1ڷtF�3_���O�i����9rDzk�;����2Mբ-�-���l�A"����܊�>3-��@>�V�3#��Z��T����	.7kQ=2Ur��������}�V�z=���������S��ڵ�^��_ij�y�~&%.¥DaJ���	Sj��Πd� N,30L"��{�UK�ڄG����o��r�e��O&�*��!M��K&�~���Ke�| �(��5)�
c��R���&j���I�Ɂ�x�tpxZ�ή��l`����\'N�|�%�D��q91��L�����,����k�^7S	e��XR��ѱ������iC`�e�:@�h3Z�y�ᇕ����]��y����}�)u����WRU�ɉt̘�Y����`�2tp�C�d����A�,�"��t]-���G6���<yO[����q���������x�����9$��8[?&�� ��0"�7���8/�gjS"g��k��[u!
��FLx�&�F`��A�U$����}��t�6��<��c_��v����5��w6oH%�O#���D�D��T5 ���8Y;������.���FS%rt|ܒ�β K':fL߷q��I{���c68�-���v���l�0�&�G�O��C�L�Þ[��$"H�HZ�Rۣ��b�F��������ys�����-���i�=~(��ð8V)��.�Zp�W�X��(S����s��@�M��(��ѱkN�=����v�ƫ�`�e5*��瑰ϻ�_���{?����X�٤��) y����(�-���7o�S#��n���(��py��|e<XL�bY�X�����<��{6�p����?<�����;��^ZՌ�p8$D�5N ᵖB�U�nln��i��h��|�tX8���?���~W$VI�y\	�6��s�,;�c�$��j:[]�d�s]]��~���i?����ض�����eM�l�E��"&���8���U'h�ޛ��|ll�@����p{k���n��t{�Mx��2��ڂ���;�N�*�S'�J���T2�Ъ*G��^ '5�������"W�ܲ��)Ï+1�������U`td�͝0}�t�xTF:#C*��#�����Ä�8vhP/���֖�ߝv��^d�����Jf:��_Q4��]ｲjê��m^^�ڙ������g���֭r����y��}����pC ����޳z��������$8|aPKxa��W�4�3�8�02x�f?����¦fo��?\���x{ཥ�bi� �R_����Hi5�M1�*U �[���y�~���H"hP+�UF�g"la~������wF�'�����d*mj{c�ޘ>ݓ��k#�����v��g�%EY�t��n��%���b�Z��66�L*���I�
T�g�~���e��kٲ�o��ڔ}����ŶvѢ\yBٝN�У���t�i	��Uxf,���07��;1(@��@+��M� xRG�B�R���^P0�L���*��INb�J�t�I>S ���,�r��P�5N=���ZN7���T�8
�g��;��!���W����:/�-����}���V��=s���ǃ����՛Gᝃ�����$���xPJ
F"���hz1;՜i�?���m`p������rMYQ�54��hS#�<9i��X�����zK{������V ��TAMi�`�ʔ����-͍�ߣ���'ѿ)�/�*V&W(r��5k^�7��慄�ڶ>�D�۶�X)_��.���d�@�a2ߧX���m7�<�*J0FGG�����?g��;�X7fǀ_������=��T��ʶ�ۢ��{�{�x��[��@�U�j �+4�(;����@��%@7t���'*���8p��3�f��$�Lc ���D�Ě�1��Zd��z������)8��Q���AJ�Ԗд��	w$Y���}f�֧�t&��}Ğp���d:�Z������i�O;�~$��~?wnh�:�j�����&8A��p��@�{�-ZZ:52�|Vۏ��{6��d��a���+�;n��*+���D�� ��"ʥIΘU�M�ZgN"����p����W+D����S��IAsS}��u��gF���#pW�RY={��׼0{ƕG>����Gy��u0x饗[�yi����.�+*H�*ę@3N�~H�O�E"��Q$7
X<c]��4��|��`(�ʺu�OaR�~�f���r�]��n��R�<��s/������9C�BxEcÂS<�$�J?ڌ�4`jm����"
�(�*��V 6:��H�i��.a�N�P���ࠡF�Ϥߣ�emk��=(Z-H`��dc]N�2i�����K�?��gS6���3h��ku@�s%[~��;L�����F�w}�� �	�m�Ұ
���e�}dr���X��i�����ŧn�qq��Xb�@$On(�J�=>�LU��e,�NfҬJ������� _,�����B�>O[�L�"&�c��C4m3)(#���O@:�#?6��llV���k��歮W����ޭ{={�ܵ�����1��v�"�[k�-|K�ZՀ��>�/t]�P��Zn��8�Y�|��M���g�~f���[��� �}�̩�F�㯛����@TT����C�z�J�J�
�.���:�!&ρ�?�Tox݄��v�75F@A @�iԛ$ ��yYi��9?�3���^���&����s�[[[}����ݧeU)y�R�����1�O��Z}%��3~������ҰZ]_���Y����> �)��!��Kjyt�o��9O�كl��I���/>��K�*Jq%��?�pS�A��/������;tٖ >L|��[��|�1@Ў��>��^�� ��D?��l�h
�|4����k�n����t;a˖-����޵�~|�U��>���8h��K��NY�����Sr�8P(f`b@q�
OΜ9��믿����f��#V�'&��#��y+��U����+E�j`���  �mA�Fj�C�����A�����(�H��Ʀ����6�\C[�@аd�2�	A ���P&As�=�wN�)�0/�y�j�Jh�,���x�&b�dy����;�U�W>5>>ޏ���]6�g���z�������3�|�x��+52qɅ��hr �rU�TY=g��_��֭7�����v���P,��P��>�O�C��!���v�4F��o�;��&���)"( �NU?�Rr��k�CT5�a&V��'Ґ����bQ��^��ߝ?ca�}���p��c���Ĵ��_��ɵ�P0h���(���uB��.��w=Qp���4&I�~�t����6�|���^ye���!����@8r���?�EЪ���*K1�+%���. �@�βKb�@%�|��[gy`V�P4򠐂�a1Zf�jBυ^���BGkU�2�R��$�B�J�"7N���7:t�)F���/�*F=�0f��rEF9o"�'3]��<�+ՎT,���s���K�=��k38N����������:y������7߂���J���[���<r�om�Y��3�ly��E���qs���sM�y�a�2nk��YN�*���(7�3*b��3'���������9�D���eV�������!�b��ɛo��]��ڃ�>z��֋f�j����-��6;�~A5L@� ^m%�3%.�'&�p��9��JY�T*mz|�ɆhӫKV,z��[�%l��͙~�l���\n���I�tW��ͯHEg6��HV��w���A�%(�x�;���c�<�|�Z&��!���L�b:��ln�V�B� b����;u6�H��S�Ū��@�~�"���K������T� �����(�Q4�u`���J���w:#�W*o�����Z}�?�۟l޽o���7�2�9V�h�u�m��4�����ڹ��"�Lz���E�4�E��'���(�k?�(�aCb%ų�U8��c��B�B���ύ _C��B9��f
��T�d�зhѲ��f��4��w�V�w�z����=��z;N�L\���AR�¨*P�M6 I	ĝ@��ĐJ3u�E��p�{ﶷ��z�����o�lp�;f�~�d��ّ�d=�R"Q��$�\� A��e~�Z��h���>,�Y�T�*�+	X� �	���Q�t�Iё�;��J��j�m�*e4���͂�xƌ����6)]d�dl�����v����X,x֩�+�c����z� ~��^���G=:�4U��UW]�tWqQ�`�e��=��w���B)�JQ���jL�U(�j�G��U�L>ǸdAB� ���l�@ ZkQ /�q�녆�x>�&`���\�\M�c���_�q���K����#y��w�Ͻ���<�{�,��3�V	�j�[��@sE���v�x��<$)�=����s��77�s�M��0�Z�o����>/59�?S��f�jEr�N�g� !���P6ʠY:�4�'B#��/:'�68�m !�
�8& @LG�|�X#X���)����%{ͨ�6���%�R(~�^k���I��>��תj`b2�l�;�=�\!tm&��50������G+e��0�z{�M]]U{���e�O�����d�z]7f#(��������&&&0�>$����@�<�,Jl�����
x�)��x8Wal"�l�e���x��m�ƍ�m����c���>��۷�w����7�x�U7G�Q��v�˪��� "% ��$����$`���ѿ�T�0��x0|e�uW��a��,��7��ez��R�]o�.�������h+W5Ī���v�5�X u=T�Ztdxf�n#F����A�G�	'@Q-���(Hxh
� V��E@���0�Xղr�z@�h`��4�)� 
X�ݦ�f��g��9Pt������'O���I_�ƍ[����ڃ��[�q��ȯ�����8�}vI&�^�~A`�y�nV1dպX"���Ln��i�Z]e�g�|���<
@���Bp_5�R.���t*U&Ӆ�?}w�M�l������ =r��-�+�7��W������%��$'����fd��|����Lm�#(a��HġPf+��Ϟ5��/>t����1�[ ��+����5}rrp�I���A6f$�D�F$�=��i�@�)�Ap�|&�d35��NX��ܹs�����@��|�*�L-\�k ����HTd��+_`k�4m=�Ag�4�Q(U��v�"O�c|b|� r����ͱ��-��wfΜ���l�m0�O��o?ޚN�ע/�C��h�h�ȿb�	e��B�c��m*�68��c"1`�CP�鑪��\Q:�Gp�M`"�+�����^����8��/���!���������m�]劲��6�./OUC�?���Z*�H��cm$�9$��ڲ��C*�`|�!���"����_��S����Շ�z����?K�D�7�����Mp���� ��S@:4�@ˏ/��E$"N���������S3�ho�Vcp�C�����Zą@}J�}����_fDJ������v��� ��(�F7�8:2�Y�悅|�3�Lw�z��;��4l�!��q���u^�xqU�\X��B^������� ����j�� �k�ff��$���,���u΁�d��,T4�*�F���^�ꚿY�����?y-~�tl}��������V���~?k/�+*�+ڊ�D �!��@���f����'5
v���>��z�lN�>2f�ۦ�{�����c��O��nת�D5B�\�����<��%�b�9F����1XQ�@��d|~.�c=љ3��{Q0���j#)
Z�Jx��jE4�P�V�@�L��e�m�`xt�4�<~p�e0�"8D��`[�kz�Xȷ��j�����vŮ"��q��'f���T*�f477�n��''`bb�U�h(��$�I@���aƎ`���KL��+ҒXc;-c�O��b	2E��u��-*'V����7�q��?z�����wZ�����g/\����nE��͈��Ir�O��鶰�G$$�D���`T�i�q�t�/�
��[u��o�[�<�}���1�>_w�u�y��O?rZh�����i�JN�d�϶$���i
ـ*:���T4�Ob���v�+i������+���q�gs����Q�L��`A�2�J�i<�r165M�@:���N�����L`f"��k)W��D�4-w"��[QU!_���|f���1�%�r�m7۳g�w˓ϭ�l|Y��9�N.����k��7T�B�~G�7�.@�c�91 �v����/ɿ�'s���4�\$�j��\�rf٪՛7���ݯ<tK�����o;����>q����aI��"�|O�w���B�/�+$�	���	�ؗJ�X ڹr͊����8f�������KF$Iݪ�?=�?,��uWlr�Y�*)��;-J߁�
pU&�d�x�^�!�ʚzM��q����+�RV��U<>/x��s����T[y�~%��5(S
��09c:���Y�(<)MR����ric�Rj�羲.}��{���Q�}�����s�м)�L�4U"b#�-)"�uD:��:�(��Z��g�^?���M ۋ��2��d
ʥ�Je�!�J�l���U���u�ݯe'��~���p~{{���[n?�s�a��cp�+m��ŁC��J"�2��|�(���NgmΠ�B"�d�	�ae��M�v��x�֛��g��>�f��>`t���X'��o<QԊ��o�,�arlD,�!�\jIe��Z�V�8�qh�e6I`E4�rè��P �e˖��A�S��lu�� ��K�*l`�T�,Y�{1��>4e;���Cat|�8��q���\ID�r9�]��dS��̥K�l;��hѢ�����Q�;v�wn߹�řl�761��v��$;j�$$u.�uzr�H�j���a�����l�*��H%�hW�\���,_�̦������?{��K+��Jx�'BOo~�SǏ�x���������1P�&SY%1%2��f:�.v=�L�U���Kb%m<mj|�3��t��Hl�H�l����=='�ͯ~��bUJ��7;dw��B*S �$���d�9���\m�yJC����K�
>���)ŵh��e��l���i@ ����@ߧ�: xj�He�MB�ϩLJ}Wzm0T�,�bׂ'/q�aZ��7������&���c�/�]x�c`�mQC`�x��\��}���pG"�@�˰�੊��4Ee��������o� 	5�UjC  pP��Z5,L�����]�ܵmF�1��bJ/���+;޸���{�BK���@�=��U#ǰ434EbFk�le��e�롡!py=�$9z#��'n��η�/�����G�lp`�ϵ[f�V�9r�I���YU����E�ڂɀP��h�3x/���ٺU;�1��P`��(��ѡ_���F�DU�t*N��>
5A&F��ϫ����߳>p{���LD��*�d�m-P�!�H �� ����D�W-�VE����*�6���
�bW*�Y���?ڼtު޹��-��ɶ���<y�s���}}��Ig�.�!`k��c�UopP��yj]����N���C�g.�UP�?H�����aqV"�-�ta�ʕ߾��۷��W>�������-��>sۛo�~��.uy}�8�u����N��T����I�ɞ�w�k2�T$�O� ��J��w��]��=�\� �>�f��~��X�����}���z�P5���ܚ�O���.
N��WjbILͱ��h5�V�$h^��	i�����2���S��Bh�ZQ��]���Â��T���0�"��Pⓓ`Z��60�
Xx���E��z!�9I�=Z�\8>41>�<�7�����G���	��f�oШ�`��kϿ���B�'�����$Z��!��&��EI�T=�j�@�u��2y�f ?$#��B�Ęs$Ů��V���8~Ţ��zǭ/��ܛ�߿��ky��ǃ۷?s�[��}O�+������)��O:��t,�B���)U-���Z@`�����:��pkG�����+_�����m��-X�@���9�������Ǫ��ܙNŦ�i���`Ǵ����M�Qd��頧��n��@o,]���8�q�y�P�� �R.1&�J�ɞO��*$�7v4��Dd!�N]ڟ�*�f j}Y*�蠎l�T����b�ڦÇޛ9���V�իw:t�{�ʕ�ض߄! ��~��m�O�����R�pe�T	�x6�C�Ԫ�D��@*���.w�/�:GBJD�L��e�l{���lV'�΂��5EI�����7����Oܴ�/~)�o��|�n�~�;{�~Av:�^������d3�1Q������)����2�%��Ɇ�ש�AIA��74L6D��/Xx������`�_}l��l�m6f��Ns��G�蚮ݧsF��)br�����H|m8qj��HZ(�!�E����NEU�@"���Z)�ߡ̃�z\n(;+����]:���9s@Ȥ�����hU�Q6����k ��d�k���/�*�������������:}񭁁�Q{���_��߶����ۖ\��s�D,v�]����/xb!%�RV�Û���ZS3=��CY;�k%߁	�}�G`M�S*+ �N3�L%M���p�M���z塿��;> wN��1xi��7����/:��E�(�U|����G͗�kc��I��>��5�`!?-����\>��^�}���⏏������Qa�eu��:�,Y0�?�s�D̈Z��5�4|��I�,�ěh��
�Pe ���X,��b��l-хA�Q,���WI �\,�� �}�/�R���t-��� +�Z�΂����2fVN&S+P�e�~nq��DX�s%s�i�b!�Ng�$'SW��n��®�Br�z;��v��ȑ#RϡS͛_z��T��d2��X)G˔"+@@���-`��׬?�A���BL�&eE�L6*�c��"���T*���u�'o��uK��Ƀ~�����'�<}�޽o?���{���y}`4�`0����{/k'�^p��
��
UJ*�f��#7������=w<pt������1�����5-��_�~�}��i��}�oK��r3|�WP*��� �,���k�n������L��	���N��C�eQ6�`�*�5bD�4u�pyX��2!�x% A�M ������D�J�4�X����XU�dd9��s���'V-�J����JS"��?�۳����޳�w��u%{`Ѷ۶m��۵�����#w�O�?Q�(sKJŭ�)l�3s���Hw5������&s��3w�F�kbF��*��9H���k%�O�⑦�W6m����f�<���nQ���C��������g�wϩ��/E�^���I�y�F�dUu��$�. �w��#=#�-��P�Ԓ�b�X�1c�ᖦ��z�W�΃m+���m��Mi1|���lT��[��Ei��Ȩ��ts�^U��`�<`��ZmG[`bb��	�F���E@�,����J�f4�d���;J������U�e��}����R������	7�㍘���Ǟ����ǜ���=�����,�,,�@� /�@B�eZ�m�)_�>3����j`�b�V\)�LfFDFD}�w����m"�J��Bm� �� �Y��p���:r �	֯�J�U-�2�"���K�bԞ� �6�"��e�8sv��Bm��3�~��?=���W���n�GH�c���a�'g���=�87=}[�Ӿ��%6��က��l�q�mq��L@�ԥW��a9Y�/ҟ��V���깭v������n��G�����s��������7���m^?��$^J�g
E!W(b��	G��d�a�����)��d
�)h ^�~�FDQw|b�˃C����}
v��7��� ���YS������'m�"�/w];�h5��;]�u P���,�C�SV)X8|�ur�n!�|���y�1�`1EFj�� d�l��:d�.Fн066�كǎ�"�S@�0��H�%K�,,���D?��FB�
�,���Ut={������O=��ȩ}3���ٵ�IABj�CPp���տ��ȡ��_1�������U�vg��*&$���BfH���8���^^�ǌuȬ!&!}��$� ȿ՗�=z;ٲ�����[������q�ſ��ѻ���<��|>�Q�CV5�K�P��y�y�{13����,�5���N�i��+�+�b�����[����Y-����g�r���G�>�X0�~knf����EҠ��
H���_5<"z�>.�M�E�"�Z��6��Da�����'=
pS6ן���ck��n���O�٩�{U�كI���Z��E�Z�>vR@$,v��� ��t
\$V�f�����T�gg/93y�G�}�C'����?]ݾ�J���}�w�^��o�Wy���/;}�������jo�OeUÐ�C#_ �����P��j� �]
I7�-��F(�Ad�7����ul7vܰ#��+�m�����G׍���[ ������~�k������O���M���5���p  �%�ÿ���ry<�a�� Z-˦h[�er��֭_��k�|���č����Rp��?�8@XY��W����,K����{��R\X��4�p`�,u䦡`����m�5�:t���]���a��A�A,L�%�&�	@�(C%�Xd�u5h�B@>J���ddd<)�J���)H����@�b���S��RP Нz�Ob��$d`˾�uU��������®'N�;|��s۶�L�����I-�_`?����<��Ƴg����=V��#�JD:K�h$�b�|�~��88 �{�M0�q2��#�ޫn�
�=���ն��a>��o��ꫮyr�.���!�/>���k��[��������P�tP*-KL}��.OA8�9gZ%�n`�.�kF^�'� �w� bK�׫C�o���w<r�'o]���IjobK�Aj�,�i����ɧ��/c��Ʃ�j7�{ȶ{�HX`d�@�D�s(8����"�-Γ��
iԗp1�鎰�$���@�$'�)�����ڭj�����pc��v��ȱ����m�����`y%��`�d8���vh��x�_����Ь/]u���WN��������Z���Zb��~��U��޻0��N��.w{Dd�l]�P�P�ߥ�V� W���	�ޔ#B��ʟ� o�ؐ#���&���G������������޴m�O����Պ9	`_�����o�c?z�j�������I�̄af��7��,,,�Vž$r�e��T���Y.kY����2Ʒ���=H��\�Y{�[
R��؍�A�����{�]7"a�."���M���=�� �S�d�k�h�t��y�s�n�
����!� �
K�+��P��L��8f�ġ��U>�T�FH�ԬG�#�.�"�H}���V�A�8�%����,�D_iUđǑ&D�`�	ʎm�ﴛ��?�ܫ/���ͯ|s�5믙_{c
ުv��w�����\977��v׺���Ua�A�A���3|�(prT]�.� 
�� �q�;�~��r�1��J�R��oJn@>C9��o,mۼ��}���>T9�����.v�wf����~��S�����|y`$�A6��#����ǉ�хs�8�F�A@`��X�}
t���o]{ݕ|h:��\����~i�{������_�_�я�����Um����'�+a�.�*	��aL�F%�qa�hx
��1��g����"!Ձ
�apн h'�Mϐ��ŅH�8��	P$	Jt�cb1�4)!A1�pN��1݁ 4�.	�����B�UYj�7�:�wOO�;��ȋ?���ҫ;/�|zמ=M��0��.^B�SO=%�ffr�NLn|�{w/��������T]?4)@F/	���'�}�ez_R� �q���
��;��AA���	Y�҈�}4b��ޜ�׵�S���|�����F�������g?{�q~��_/|�K_}�+���G�lq�/
%�0e��g���t '�@��!C�"<��Y��h�vL��[(珔���sã���?9������ �_��ŁK�ْ��ֽݻ���>�J���v#z��c�\�c7DF0sa�e����	�ꫯ���$9�`YF.��&aP��2,\�V��e �����B0�"�X�!s�a��jo}��_��0 tT��"��c6�R�ࡼ�P˷��U�zc��3g����kO���+��t��}3�#�F�2$�]����Ӿ���T�=���̹+��nh4���0��ڄL
r��q�� dr�c�ĸ޶+�K\��!>O�*��	�����H��ݘn�͚�#���ڲe�3����|f���X��n�?��~�޻�;3��J��ݏI^�r���4��������/%$e8N
F�x`�	 � �L��b�on�����'oM��Ef)8H�nK������K���E���N���>T&='d�Ht����Ap ��Ry �ݮ�Q�"��K��aX��R�(&�
Eb긠��Xi�B��y$7*�~���q�.ơ��c=E��D�r�� t�R�1v^�����%��"�F){~X#'׳��z�ҩ��ǎeh�����_���\��$I�Mi�}�k�N�����GO��v�����z}w�q�z�_���8��@"xIe,)��s�!�{I�X�*�|"+	( ʈ���ri4�i��dÖ�����L.\�a��K.�z����{3��Y`�~�>��-�N���\��΋��� ŁA�Eqa���&�bW �}}��2�д��إ�`b|��j߾����w{
.JK�Aj��u���Ϟ�ǿ�=t�@��h�kq~iU��Ӏdm�Vhc��ԩS�Ci`zz��!smy�"��5vZMTa��T���^ZZ�Z(�I�����G�b�@�%>� ������Y��,.�k��� �H�(��U�m��>$`%�AS�~a+�q�c�Y\��ڝ��3�;|���U�F�lܸ�'����u��[�Zi]��a'|P;�����Ï_2y�������f�2��׸���%A�UBW�$�؁ 7�E��� �;g�Q#���Z~�+��H掀�8�&�΄��(ٰaS���G�ձ�
z��g>�?~�������~���˕�����j��M� :&�H>}3b��tT~<��d, c�S Q�7b�0�r���a�߾�|���?r6��� �_�]s͸=�/������g����Gfg.���@��	�6 +"%ҁ��Xu��,�n�ԗj$kf0��r!O��"xd�e�<K:�G�^Y Z,9��49��B.����	#�[��&8`d-X���>T�x)�B3�=�:�J�yn���L�ر���������v`����?��Ys�Pkc:.�g��wKO)������7߻uzz�ʹ��ݶe��L�&���F���$^w��c���?�/a_����}p�2Q1}�G�C PFP�r`Ji�ץ�t�\�m3)�]��Ӛbܷn�v�3��������pg���寮ط���e27�iT1�*4(�
z�2�z6�3:f�B�� Uem�2/k@)D�����6�M�-^�ƍ�~�����dv�Z
R���ZAp�s`b�\��O΋���S�3��"[p|}j�^''(@ز�RRo6H��Bg��4����>�rx>r��&
"A43Z��X����t7�t�T� �	���ɀ�1�>��B���O�& [�Ǡ��N�S���LFI0� F�A/�lO�4U� �T���Z�gN�����3��X52���������e�]�N�߬��������h���ܮ���+�jK�)�Dy؃ԉ�a	u+��� ��"�0f:�Wp����W'�@���A�H��-c��pu��\�}�4#�i5;�GGG�߼��W>�]��q����������<��bqwǃ��M��F�3��ND��)(�q�H���d�d�"�A���o]ˊ)`�������/ݴ罏���n�O3��� �_�хR�gyd�7�{�=��������K�5���k��F6mނ�V���^�	��ei���,Ҭ7H&W �A�d�&�7�,��L����"SS�c���8���a;DsR$�k0ڣ�(	y"��������f�(b�(�������n�k�|y9�D7�J�Jc��t�����o?�9���+//��y�W��s6l��U��U�V��J;~E�B����3��]����<5��{~�ma�~u���b;��=k>�%Y���|&GY-y)PF >
��6%�L9�M��M�ǐM��v�%Y7�N m�>/"�q��z,�bmɫ��O���g�������!��?�g�����ο���;��n�4���*�D�Cث��z\�C��u��jȎA��I23�DR�pl
zwGQw�ڵ�KŁ���={����4o���v�[
R��h�?{��3��y�④�l^�o^��]�����u��^�G������H��v��0$	��A� �24*"}H3WJEҩVQRd�c.U��uK<
r��[��B�0xD�k~,D�k03
.���Đe�GU��ѡ��W�R�b���z`w�h��F�
k�cQq���:�N�;����{ff~���&�������#�6l�_�nj���Z��4�)O�n�D��D�����C�����cS3g�k���/o�Z��cq��x���SzM�`Ab�%�� "��qZ#��ZB�/#����g�`��q
)�!t��0�A�S���Y'��0��#G�����kן)d����MR��m}��_V��O�l����y���_������4�Ē�/M7�t8/�@�N�}�j�ޯ�j�(��>�:@[��s Df6�za�Z��M��'����oK�Aj�v�f|�>t(>��k?�o�<��(��z��xi)w��q󥗓u�/!펍R�(�Q��<�E�i�нPo,��z�A�}�R��
�ϟ'��t�`"������lp��b�������ś:�B�}�}(�[���c�5Q�l�A�B�` FS�K��pn��X��_��6�v=�7�ѵ��u�"]}��L��'�9�Hux������'�M�~��V�S��{�n�'���ف3gΨ����cwݗ=�8�j��������Z�~i����E�X�E
��0�e�f  ���grjoiEQ���� �)�sbN6d@ �$@�!d��d��?\�pފ�{�[`��z�����}��#�L6�M���G׎��h���������uw��W�����?��e[��2�����T�%��Z�E��~ATT:T�7�K���g8���m�'��Mlz<0�<7P��
��l�d˝�|�?��;R`�V����m��.�g*��o?�Ѓ����1�U�ѭ�:yZڶm*v�-�9άDPXp��b��f6O����F��,i�sH2�(-C��HH�0>��Œ�-ig,`�'b{"j+��+��Qeee�����X;�c��LuL.�'@v��2+a�n��De^� "cdzNhڶ[�5Z�,^}��T��}�T,�8328x�4���'��|���714�n�S��C���NGo����TΝ9���l�m.5V5[�ݎ��F������C1R�(��9p���9� ���V��^{��b}� �� �L �Xd�0x�OI&��`p��C`Q����Q��K<�j��J%�e2�cC�'G��&֗��7z��^��7��=�'ϼ���IY�U
UU3��I?�� �
J���e�/�� ��hbI�����\a)_(�xǥ�������=��l���R����~c�7�U��{�ɗ_}�c�f�3�ӫ׮[� ����%�	<�����Lc�Z���Y[�K�c�iu��ET
$2f��Q�G�q	�Y{d�Y��X�5�C����U��BqE�~��.��pbY̝CRr�0��<QG��&0��<�ˣRQJ���B2�O���.5Z�5�ӳ����ƒn���ba�R��V��J�c���ݳ��`7W��t��ݻ/��B"HD���xfQot�|�{�sK�۵��F�5�:����Á��7� R��iA�y.+1� ^.Ba%F�XF����.�
��ܙ@�
b!�<0 �KN!a�"�#~?�}�ܛ�D��@�Tʃ���Β���Jb�"Z�Ã��s���ǆ��˗�G�~o��������ݬc��12�aj%Ȍ��@Aq�R�*�L���� ������ �(��4zK�������Û�m��o��K{v�i�ܗ���� �ߨ�E�I������Gy��(J0==�n�Ν���!���
�ı%QQ��p�~,�K�C��� 9� ڰ r66�E�:x?}8�L�����"�>[�è�!��)`�U� %,�|2$��w.$�v"O9\'q*��*"�Sp��|	�0@�����>��vMWuE�!��ڮ��|kT���b��ɞ��mC�k�|n���Δ+'���|�|�`tF������Z�l�ڵ+x3.�T��X���ڔ��͟����VmC��Zӱ{c��9�S�����A��OA �����A�
����],��M �'p�LE��{�#^ъ��!�� �,�Τ� ����}�vll�`Е���
\ʊ���|��K^�f��=����/>��m�"�O��	QQuM6D#�GEC�$b! j X�e؏�������cE��b�8W��ʷ��ۛ��Gv����Gߢ��������g�y���|�G�<��s��\7<:2��t�V�!�VO�&��kF,���ת�F�D�Be��+8�t�A@t�W�)T�0�d�,J4b��mX�čx9@d�Qد%G2�:�*�16U�;wQq�^Ҧ�D.���.a�u�;��B[��ۆ�K�h���t�0��T��s�� j���4!�$��4]�躶���b&���e��*�g{�������@.gg��r>�V����i�eY�V8p{kLv����A���	��R/?^� 9L�^
��ǒ�`~^my^�����^Ǩ/4������m���v�[�u����[eu����~P�]'KO�!ʂNO�R 'd-/��"k��Ӏ}���)a��+��R(�!�V!�^C:�Ā[r�XL��y�מe��!p�Ж���W*L��>�]�!��~|<y�4�W�����ҽjF=3�p~䡇^�bf���=��U�d7.k9T��]F�Q
2C�S��s�k���{���s|�-��bEQ�j�z*���u�{��W���SB�-xK[
R{C�u�m����dx⛳�_?z4����������̌b9]� �aJ1̔ouiҡDq�L��+lH��`� �r��e���Y�32]PQ`4<��#���>�1d-�8�G��� �e����i�~X��D1�F�X����?Y��{����P&�I�Z�eȔ�t����2=��K9�9��Nwu\�,�C��(}�G[Ӵz6�Y�uc:kf��w�l��7�uu�)�|U�t5ck�l�3eK$k�#?�ԢL}O� A
$��p��}�;��^�v[uEz��zJ�]W�p<��,K�Hm�Z�纪ձt۲�^��YV���uG-���9�n~��3�����A�/K�����X
,q���p�-��hcs�zV
_����K�e�c.�ɮF�dY���	Oϣ�����V���'Z�'��d���-���P��͚���O?v����ۄ(�*)�/�\%��'���3��za���'��EEZ���-d�����bI��1u��'R0r��n~�}��ĭ����}��[�Rp����t�c�=�j󅗟? 
��^���Vk���Ca���`,�縠�NTc�.��4��dp�#��Z��<t�6s��ֆ(�Y��2.��#
�~jRБ'�|m �~�2�� ���/3  ��,HWG�E0�K�&�NL ��6D�+GJCI$��%x#a�D!�#��`�g��$K��X���	����Nz���>ݶ/K�/+�K�����M���J����(JQ�;�g���H�ň�'EsKR�D��Ht߰C)�@ÂH^�ka�g�9͂(T�^AG���tz�5��T���CP膕���gSD�0�Yo��<��,�#�t>?��L�%v����A͐qC�r�`�a���� ��\ ��F�s�S�ɽÈ���H���D^j�����d��[�$�1A�3�u5h6k�V�~S�c�˪8DϙI�%kd  8��p�p�t���2 `@)@4Pj�y
<�`EE�2�|m�Z}i���=��G{��WN���Z
R{���8�qc���K��4�l�:��_�ХB�X`�0X�!E��g�{![(�b�@��P4ɳ\H=�&.�ܙ���.�2�w/O��L���f(���	��7�:38]����EQ�w��l\MQ��eu��+.G��
I����!9�BT��<pP�N�,����fE洒������'B@9��2�:
:�(�}D,�͢��GQ�O�C�lEM@���_�Z���7/�1~.��'0WG��-D �  ���B�+&��Š-��~z��8��,��!���2��Ho S�P#F�xM�u�$�|~�R�x#0������`p�1SȄ��&^��������dz(�Ӆ���)��)M�N���'��Y6KD�@:�#R(�a/B�^ϻ����5����r�P�����2Upb����(�j��'����� �C
F��!������c�l���>���ܺf!��H-����5���:c��=�KK;[�λ,�ɸ��Zv�b �r��Z�f
��+�ɒ*Ly����$)�"��ɞ�є�ɸ��B*F�@^�{��$ �d�$@	�.�����̌���=��8��9�Hf�
�m��1	Q=��J@����p�u�.3
<|���	�i�F���Z�y q���1F�	�Q�J�Xaǈ^�����Q(�HC=�X�g�?�G�
܅@�_E>s "X�Nt b6s k�t� ������I�*0 �$�gd�@G%6R[b��EC�h	�$|'l �,8w��a�!�0چlB�!e������q["�7 ����Z���^�|����AZЩ��e! %"p��)��L��	�q�F�e���3YSȘ� ��T��R3]8��(��=`AF�� (!sb[.�wh��@��)���ɗ�F���\{�u���;�{��K�)� ��������i�C�=|���� Zk[�f�� �"��<�O�6�r��LX$MC'�]tm�@i�zF2b��}%��"eq����9䈳Σ>/=������X	-e\`u�.�`q#]cK��Ɍ��/ϸ�0Xno��s�<����1َ���~��AP��}#Hd�c���?�X{�&OƼd�$��\{Ϛ�b��c��X��3,�B�N1�*�sI��["qM�2�`e&K%p� &��Z�b�5H8	�H�MKx(n$���1���b�:Wpra���E3T@��rVCR�uphr ؁�0!�$Xz�`�7��/W���C#Ě8}Ѧ�������&��~��2��J!��ԟ&���|�R
܃��4���K$p�8��w��FT������߿���i� �_d)8H�Ma۶m������7������s�uls�~�!@\X�a�>8>��H�96��ebJ�����VG���x}����E�g������CZ�����(�:���� �^a��\�Jǧ���Ls2���f.�9�'�_3��
��c�3&�܈� و`Fr$�vΜ�@�>�M��ӆ�,�s��JE��Fb�Ȁ��	{�	:���^�<��$X� cP�9�����:���������C�0 ��A�I@�y�I�Q"S��\6*�����9�����H]�͢ �2�$ʗp�����"�z�1�28X�������
�0b�Rx��X,����?�� �2�p���|?rc(�HNF�6X�2S�TE��b|���+	�������Z��g�Ž�V���>v�7]�c!���������={��8z���>���u�H+x�GI�ԨӇr@�Fo:��L�F�(T�E�}��a�[���#�MB��-�>�1���j��� @���S�%=�HU�:(�$�QK����P�ODx-��a(�8�  �	�"a܃����"*^_��8���Z
}5F�Bd)t 8�"f��pi�N$�����d��O���UP��Wpt���dc�~$,��Yv���D`;L��E���G
��PJ`��Aq��,��{��Cy��p��r�@b�Q�X�`�e��˝:l�'��~�#$*B�A���U؞H�d�H��|�^���^�����D�Ō��gY����.)����f]0�9�6X�b�t�28�ؕW\��[���C;v�Hj�������4$�W'Ǘ��lg���m�u*8w��F�auZ���� AUh�h���x�xR�1����]v����d. P: �b+�و�8��jb���k
cQ�]US�������xNP�Ql�>�{A��HR��0t$�a�"�h9=ΦP�Oء���J�q�A�Z��<!N~�X�N��xfb	�2}�@�c֮�ҩ&��	������[��|����O~Ϙ��a�_�LV��\p���B�?�0�`���"q��0�N��@X�z��@���K �`� �V��,�v�=�ԙ�K9-CѦ�Ԙ�B �|�!�� �(���eC$�ː5k�  @�l�����ld�L	� ,1$b��.2݌��%�^W�N���B�H��mv�__5���ޱ�ɫ�x�$H���R�{,���l�b����^j�6ږU�w�u]��h����nu;�A�n�� D�
]x�>�zġ���U�D#"u��L�K�q���,�� ���E���8��@��@�Iv]O24Pm�͗��O�(���H�ꮦ�WDI*P��`��(	
oq�Ҽ�s2cb+�e��&�Y�I,��L��b� 6�:�,LF7!	
���\��)�$���äe3^v�%?��ĕ�`�ujp0��ȸ�)�m��� #���e��;Ov��ǜX22���h���|�DBF�AL�AЍ��F����uNɂ��e�<�������d����v)���k����c�a3e�B���޺�bbnn��qG����٩�ke���>�?�8%T^��@0rm��Q�B�l$?�/�M�O<Y��c�������Hgp������2 O��s�,,���v.	��&�r�kхҧ74ur�3�K$�s�nB�Y(�b=D���#j���u����p�C�����)j�
��#$��PۆR� ���
 ��񘝞��A�\<86��qI���5��u�fskkDQ24%���"QoCK]�!�����W�Ӹ�Aҭ u�X�N"$��L��t����2(�����s~�y+a�B֐A�+���_x���<��#P����DI����D���+��o"?ZƇxݝ)&Q�J�"��I�P�*X��{�S#�<[*W�O��8<2<t2��7�����;�^{�ݬo�:mzٜK�l�ȗl@N����+0M�4�M�0��f���%��,��@��4��p�B4�W��}�L��9��D K��X	�).�C�:ZbQ�l3�?�qæ/ݹ�߻����6I-���� �7��(��}���ް��g��ڝ]�(�A��VD����t:-�X+Ā1��e(8(��G�Dd��5.�(�q�����U�ԐDw��c����d(���*v]H�
�ah�Y��`������3�MNNΖJ�#��?޶���s��������K۝��V�]C�7�(r��W��� *w���Q_�R2���K�B�D���F�\g!����%+4P\�;�~����u�!�;䨟�_f���2����2��) �����1J�$c�T���$�
&"�,I�=��.��C	�J�[�"�B��myӢ������l=�~Ӗ���D]�n�k��g�v����jo�Y�5�e�c�c�����Z�1�#��844���������`Y6����j��q�\��A�3X��õ�, a\�9��� ��HpP�Tb�ԣB���/�_�v�w�q�;��䇮�����p��˷����ݻ׷�}�У=�/xQ\<{��z�`�n�؍����p��Y7jK ��|@��s:����J�X.��AӘMH� ��u,�&�������������;��*���tM��Fq���(�	^e%U���U-��p��]G�>T��2:����]{�B�{fgV���^٨7/�]w�F�C�'�)LЩ����E�����.�'� ���Q�=F�fKB�������I��"$Qʲ�Z*�gWh00,����8tfXf��cP*�<��O �L��'T
�\��{6+J���]���l�"n�Vd'�Sd�ADa��A���F?�L����es�l���Ƶ��T�b��_�#}��wK���>;{��۽KzvoO�۾������\h%44��E*�2<4�e��Μ=M��6k�UTb"_E�L�/�3A@� �D��6�3p�bg��ܮ��,Lc���FDz��tG�l�.�
�������z�}7�v��k����&���O�����k��V���g�_j��َ�[sSSc�N k�BzN�3:		�� )�DQMR&�\U���E���A��vz�`��
��2#껔�E�P��P	��B?"f㗱���<���!g�tE�5������u�3���������Ucc��n��,OP�XX\�_�4��q~aq�u�	�T�E�����L�l�q$�bAdY�a�m�碃g�&el���KUՙ���'�`�����U��.�(��I��g��wP�T�ǃ`+i)䭐	'�K	�Χ$��K��pm��"�\���{�1� �z6�
B���C�hGյ�|�p�X.MV�Z��h�:6[��=������(��ϐ;�C}��{����cq썷������uV������U!4B'�|��1 uN�񁥩ZU����f�n1K�g:$8��Aa
/�s�hX�lz}e�I�rb�Pv��130Pٷq�����g>��w.�ق���������v��.,6�8=k��uo�+l��iH01хvEY#>�2�]�:�"k 8c�\�B
���T�����#}#�0�f/� �RA@5E¦�	�K~^&��cP)�����(<�.�2t/��,}� kgg�n���>��f&���#�Jyzlt��͛�����j�gg��,..�4��
�d+��5Lz�:�u�:ݖ&�#��E�v(�
:� LH�x���$p�B�@&N���Lql���Y��%NL�H�5�|~�G�,�F�ق����y
��F"��h�H���a� ��:Г�J��� u�!��<ۢ$6%I]�r�r�<_)4FFF�JC�ɱ�����BA6ڥ��~������$ 
�S����/[����;�ںV�9���V�h�@M��6D� 
Ο=�:��3A�BU���8_�GL������%��de���dzB�m��F@ �!�M���j]�dU�G�����}�;w�z��6I-�_��� �7��z����f���U�0�.��LJ��4���E��Hmq	ӻ`&���N¡!l��Z��a�R�{�s��O
%L+Ȃ`�v?�K�Qc�БaD�P\ɇ��L?G���u Qo9{~�S�'kԃs������������'w�<��Hjt�zc�QnZ�J��l��Z�^mw�U�N��ԙdY1��%�T�Ƥ���B=s�	]�i$������`�c��S���̕�
A�e��yI���%�������\�15g)���6��+�G��EA�E?O���G��ӕ�������������B�4�TU�)u����|~Ϟ�I�s��N��)7��K��oow:W�a��u�J�X2��#��g�aBZ�9{�,D������R�DT����Jbd2�:)À�dT$q����H��<��E�dd�L��c��X��ѳ��=�m���o���>��i� �_��� �7�m�Xi�pd�v�U�,�(�⮥�Ec6���E&8_ g��p�Y
�<)���U��3�x�i���@4���L��}ޅ����,jG'��� �Wt�Ё���@���L�}���tc��+X��k�O�̨��I]7����cc����.lܸ��!uNB������Z����B��*/.,UZ�ސ�8UzD���Kv�[�axIU�Q�*ı�"��D(Q����9���BL+y
I��yH��Cb����b8&@��0J��LQ �D��= l�����MQ�����MÜ*J������j��/u����g�F�hU�A7�Y�?��G���s�$�����=z�h����e�*]���K�͊,�T]���$��aaa�t{6�P@Iȭ�]Q)��k��+���/؄{�J�I��qYbbp"+�ixa@EF��Y7Yi��TUT���Ѧ��?�~���m��gv����FF�t.Bj�lK�Aj�]�eU�'?y�G]�6_y��[�®��i�8ޗ:3�:��KT�n'�1C��{�����*td3������	�#���H
{^L4�} ��҉��5	�S��Z����5 0@F#��A�At�e���b��d��c�Fkjj�>55=+I/�3�W˕ҙ5��.����;��n���QdOl��2���k7��V�^�7����F1��S� �5��Q$�H�5�:=m:=H�y��D@;�����}�!�ѧ�(���BQ b��Q �H�`i�ٓť����1!�\1�,�ˍr��,�J��+d�V�T����Ҡuv	�..Ƈ�����������#��/��/d��Q��]ܠኡ�ʮ �8�7�xnvqqA����q�^a⡦(t��Jd^N�(���@ل)&��{�=�~� 9\1k!���	�RA���g�1�/�CCգ�b��M[.y����UWm褠 �_��� �����˗�l�{�V[='��C��n�=[�( �����!��I�Q�\��Y�\!�
x�HS&7L�H�1�C���3#ԏՀ�T�:��!0%6�Q�D��ߏ�����A��y+!ԫU5�߻�+��)@���$	�\.3N�s)u>�
!u��S�gN/O��Y3wn`hhzlxt�4PYX32Q7�V�P�r��7�3���M�'7�@��)���uD۲�VӖ;��R�b�e�n(��=����LC~�F�b�c%�{@�Q
���( �cA�4͈�"9RC�4LA[���h����ǃ�Bhd
��e�bY�$���[����w�w���x��w�+���ɤN���.�q������ڝ�.z��u:֘e�ʵf#ױz
����D7aR��'?&"D*����2�(��9^X�U!^�qa�1q*�����:p��"K
��ުU�N�J��׭_��u7\w��^�����~Ֆ���.0�����}�>jJ�|���s�#�W<���A�3x�V'g�I2A�Ry�:j�i��!
T�x5"U��9��<P��d���~�ȣjq�cX��&�|;`��=�v�z��h��
H#�Y����#��;~�a������N��%Y��~���ɞ�\8\Z,�L)���K6)�^>���Jx%�?+�z�;��'�'x�[�n�X$���7��ޱW^�/*�BG�[����?g:�N�^_�#�Ns����f�R��W�z~�) ����dr�>���|6�J� ��������4�क� �!�(@|E�&d���IIVD٦a�.��[5>���_�����J��S�uY
R����8�w�|��Gʶ[�O�]iܳ:���D���8�0DR_Q<�8�OF�V�,u����0��ז����`b:��0EO
YkD�غ�1�$���ԇ��\�/�����Ȉ��A��s`?@�)k�Xy�NBTHiˑdA�F"8%�0	���:={w���R��<q�hS��y]7jf6�T5�],��K���l1����������Ɉ�$U��!ѧ�(��k������ ����9��?yJZܺ(�)"-j�te��/��ܘok?����p~a��Tq\{���T�k�gYc�k���Jy�-S�4E�AR�x��ca p�`�D.U-0.��WB�de0l7�מQ�6�*�#��YL�sI��=�Ȝ/�˯U�O��u�s��jj����fR�uZ
R��)(��N�.��̥�����`8�]��#��'��8״��M$�s!�\{�Y�y�W>Ē��H��3۲H����0�gP �:qNV��_r�֖�r�ؖ�~Vpeԙ�|@���b��JH4,�&�H�H�[��E�_��w@��_Cp�v�%�pg�M:��vEIjJ���M�chzK� �Ѝf�P��^/��?�c�����݌�qL�tEA2f&�?�����H�홽 �5�EY�$q�A��h4�3� n)�'��עTP�Q���X���{��ZN7�:^��h�v/���2~f��Vŷ�!��(B�AW9zNz�zg�^%�Q��
�s����'"��Y/O|��j�.-�$\�p��u��غ(r�f�]0��)��I ��d���:u���g^,�ϼ�mW�t�����jÆ��#/SK��k)8H�ݻrr�x��}�'��h�x�����ƒ�s�3L"����	0<+]�#���42P,&],�� ���܁
B�R��L��:ֺ����*>�mi�˅�d�?	1�����;��p"�g�+!Ip81V�4	`�/��8�y|��P8I��ƔQ~7�B?�c���������C�жa��]��Rm���Q0 �4��[���TU��w2z�kf����Őۚ��%E�eI�TA	"1BP����T�~�v�T�O�G���P�&V��"�wܢ��%?2��d�/x�����B�p�P����Ǫa`xa�Œ�� �tM5��'� !�TUY`/I6� �hA�|I·�?��w]���Df���Hp&��&L�:Pb���c���+x�$��!�/�㬙�*��a�?)�O]���n����v��C�R�MZ
R�hm�ڵγ�Ͽ��W�}�yR���O���kK]�'� S���F��:������*J�u;@�8�N�
^���"�\�`i ���C���e��A�ѩ�>�x�8d��p���������J0�X���G�l�[�<�~{���(����
�8��:_��"��s��8pr!������v#�)A�!����&�cz~�s�=y�42���$R` �Mw���FB�]����"��e�x�ѽ��odzb�8�x`�����g�`c�'�	BL�%��P'�膠"�b�{-.�G�D8/B�J�!'��N2�����)��LfG,�TX�`y�4�Ha쏻��m � $z��B���fL�|i�R�{ɖM�]�+g߻}{Z>H�a)8H�6З�;9�J D�O�z��L��p�ݔ� � A`JtԁC)�Yo02!]�@ȐR������ԁ���	$2B�e�"��'�Zc6YQ�Yt�>��sj$P� K��-�AZ�h�s�/H������kP3�.�:F}~�2=b�H��J�/�A�,������0��������D���H����PJ/4��~��c�$2�E��@�ϔy6$0̩&I��ȅ���4J��xD�07Bd-� -�j�5��A)��Q>))�$n����I �1�d)$�(��_�(x%�qQ�0(����`���%94��TmF3���|�b������]{��殹f<�����Rp��Eo7B���hP��g�~&Z�n����v���H,��!��ue�{C���J�:�@{���lA�ÐI"'�,��B��!��u�D���0	|8��~�B��ك����ȉs�8�>�� $�^+J}��tU�'=r�cr,�%p�gt$$�6� ��$4�Kb���,2vY:I�
;��UI\1�9q������TB�y/\��{��t��&
���up�0�5dEf@��i,�(�{#yƬ� DB���r�
��}%L�.N6�"(�j�1����|.�w��կ�m��N^q�xm۶mi�AjoHK�Ajo	��lrr��(���\���|�:�	������e��d�:~Ǳ�3�X��Y���A�N��81� �m��0d�2�B�j��{э�(�ms�$_⠁u8�c[I��;�d6A22�A�]���#��5��,��x -v+�m�V'�H?��M/9�lFc���E�@�SU�Q���F'>RѰR�||	�"N���ؿs������Nv�AH����.@��c(E8�:cj,e2�����S,��$p�[G�ㄝ��C3 PT���xR�6	zy|5;̤����e
6NZ�D�ERTG��v&���u}y`�ŵ�6صu㩉�w��CRK�l)8H�-c�A8q����_~яB�fm~�%�$!�,��O� ��h	dj�q<�@
E
�Y�M�܌a�V���'�٥NJ  ��]	t{�b����}�|�� =�;��R�FՆ3�#���À��(&&-�,��I���!IWE�B�8��C?J����c� ��#��}1-���Iw�ò�8QQ��r0����M��_��>�0G�rNc�U`�1�(��	֞	�''&� !��n)<�2 ��N<�x�|�E�B��}.�-`�M��(�@;a����H@�`���(hV2X&#<���^�PVTK3����ۯ�ځ���[�l=r��k��6X72���R{�[
R{K�ƍ]
���ҷ��1W�W}��T���4E��d�n�Ol�M�8�E\�&m242Nt���ɪ*i�,��l��8d����(�z��:�`�h�Y5�u��ӳS�L���%mX֍��Q�A�I�	u���]�F!�g*|b�S١�2�ٞ��� ���1�:���,�I�o�#���yZ^�����z�s � ����M�Йz^��-�)�@Τ�%�;h�G�1��������/�B ^q$1��� �{H� ��V�8)�DD���� ��d��Ь�4�;q���  "�\����,p��d�#��N�$H � ����J�}_5�N�2pNW�WI~q���/_z����.��ذa���#��f����3 ���;bdK_����K��;BM�Ա:F�,��s�4K�e�4���QZ�즙!9S��*�Q̺A�B�G�N����<p�m�Qr�����V�I&���ꪫ�|w���C'Ol>vz��^���z�J��.�[���PԦ�+c�DWT��:�υ �	���ʍ~�18meJj�A�\�cR�e{�"�r�?\��'�"p�B_&���'�� �dp��Ɍ����m%N���;������0�>�+Q�'oB�l�\ւH��ˤ͘w��,�D��k �[Ʊ�$WȽ`] v s"Ũ�I�)��2r��R�����J��v^~b瞝s{֬qӮ���̖���ޒ�{�n����$M���>Ys���&_Y[ZȐHM�@�}�����f�x6h"Xdpp��J%��((0���$�5I'k���&�N�t0�H���Q�Ѷ��j��mo?r�������ju��;/{�+w?[�8�����]@l���U�n����(0��:|Z�C���0B�G��W��!���[N�*�
��
lDrґ��Tٜ�dAgJ@F �R����숳����d���%%N��l�d߃�\�e �z>�&#�]�3n;������jD�0��+�ā%��p�0P��	��϶��LE��������v4U�+�Kg��b�������u;v�?�g��j�v�X
R{�O�.��{����v�?�i����lw0}YV�L\������F������.�暤48L�L�h�N�b��fF'fS=  p4��5�T��{���g6�>~b��Pq��m;μ�ګ�k����k��ӓ�OM혝�]��y#A��i�1hFF�� E`僤� I�G�\�fB�s�W�;k�v�[�\���ڡ}O���1RL�(�9�g�-a/�C+��5��!�?(Q��E��DD�l�A����3"f>�m���?L� �r kL����B>S�����["3������Me��S�b������5��\5<}�Ƒ6d�Hj�]d������v�m76����z�~�����wۖ=x��� a�<D����.j��g����H._$�B��fK������LK#n�H,�z 
���M_�̜�;�	�wn�/.��G]x��g����ܸq���n����v]s�e7�z�Y:wnj����湅�M����:�AMQ��4�W (�lG�f�t�#�� X�Iy̧�6>���~�!��&�h@� p�1Snį��H��r�?��j���|F�� ����h�\�aXi}���t=��4"r�a� �P����XQ?	!zD����d*��f��Ɯ�)'��G&V�?1�v|j����5�<��.fK�Aj�Q����C����^y��s�oi7[���F AL���4i� G7�N�D=�>��AB&Gr�.�>�N#lӌ(P��W{g��u����:=�}%	B�\DKVHmVb�q�T��%]^󚪔���#Y4c�")	� � 	` fzz�rϽ݃K�[�����V��������r�v�J/e����� z��(�����k/��;U��pza��ɹՉ���Wοt5�����vm�pfc�ɩ����ϛ���0���X��j�U��F9pa��U�Y��o�ͷ�˵Q���`9�Rb}�9O�W���j�����%�s���y�BiX��7��0T�EQ]�S�:
2�V��;,��G(6�H�ui�2��
�b��T*�dE�U
��ch����Ƚ���ۍ���Ϟ[�il����������
(�dii���Gŭ��T��{�?��������K���C"�i�,��}M�ҘP���.K���uۤ�9�a��6:�6Rs&H�G��:dŋ��Æ>�L��,��Q�}���N�6=4:E���W��wWV�,�l�l���X���||lf���7�'�4<��ܛ__�x~w{w�:s��� :4�ي*��)�y�Ōr�۠%]���?�̳��]q03�_�\���� �|�zc#�W�� ��E�T��  gBe��2� "��y4�{.ݒ���m�<�����"�n�X�TҌ}�V_�699qk���G�ss���Ў:ީS$EA�|Aq� }��4��݃�����c��:8�Z����I�Fu���}�y3#$�J�i��:�]��Z�Ft�$
p�*��a��ͯ,��N�}���	T(ص��]��v����1I(H�I��|���ѣ����-�4vk��6s�ģ���'/�}�zI��������t���*>N�ۇ�i�N�E1.'��$� ��"@�d%�W����t]����w@��b́:�����E�}�b@$�Y ^7p�Y8�/QG����YB��4-�<�2��"@���#�-8��Q�sfY֎����������w���t�j��IY�c�� �n�� A>�w.���`����ۺ��z����OeM�~Et1�f�(diH4I#isKah]��T$У��2�V�>Z��:	,*L�b��P����
� f�IJ]LӀ�IV�4�iqjE���J>L�8��8�k������,;�saK��.}_d�F��Իã�w��F��w��q/R�1D�����մ����e�Fo+�oEeuն�X�Ų�A�H�%�'&J�����T3*g:���[du�l��|�}+\� ��<��:��P���Ǩ։��(���گFG����wW�\� � (�P�m���[?�k��k���󶠨�Y�;�_(Q�6:)�~�#�u�6�#u;��.��VV�&&=�FlK'��i
C��0ӕ:�}_"4�s�!��̀ )fYb&ad��@L��ɜe��s��^����v��w��� �^�J�o���V�)8"���ҤV�`�N0����Yf�[�7�;!�硎�
G]��w2����h�<�V�Rok�~e�<^�[�:2�v��?pTA �� `���V��T��<˖�����|p�o���W0C� ��������J�������W�޸w��ݎ����'I��{(��,*�a/�f�U���C�!;�S� ��m��N�`�2���Og�-c�z���bB!�" & &y�
�D%!���,�U8�h�i��$rq�C`����
r���������fLp�"��a{�VAR�x���M�dèT��(q'C�uK(G����N�������-fi��'��?�	U#���9n�6�s�C�el��pN���q��
�Cz�����߾t���7.�q�^?�����Aq� _��%!���ɉ'�W������;�?�x�N��ߓeq2�B=
}�e��
K�w|* ���#!�B"S��v�,�jt�kY�L��,�İ�x�-96��>�,@d'�' ���| �(&**�`8X��`���J9�*�܈��޴ǜO�����A�X,'�	 ����1{l�
�:��*�rV�,�,�P���>APmT� pyUe*�Ǫ~�Q�N�YJ�(fߓ����న�0�{�"�=u]OfǦۖi��u��/.�� D����S$�l��iP ���f�H���˯>�y�7+�>�v������a�|�����'{�K$�J�n�Q��N����!�!���p��˶��A7,^4g�Ā�*,,*��/�B@�1�c��F)G�f����@0�R� �PN�b8CЇ��`���,���s%"���]��D(x]���l%OX&���SpU��������2�#���VN���Q=W�0aXΐ�� +R
�������14:��C�E6:�hS��ЮY�����w~��͡��I�� A�8(��H��օ��k�.�^����~t��ۇ��U_ee<
B	��sBlJ��o· ��g�#A�#�e�����D34Y��U�M���*q��l0��}�(������	��@�20W���$c� �36Ȩ� ���3u֖N��%�Cbu�w�4����&F�q�U� ��o� #`h:�~�%1�I`NEe�b�E�(3!�Y����!�����P��9�l�i��#*��_ZZz��Ko����M��}� (�Ϥ�$�ip�~y���G\��͛�����[����x�u*
�"K�$�y���4~+u���O��� `+m��[��Z�>oJ*I`h���H�>�i9Nl��4<l���<����V��X�j`s5հ���~U`Ȃ�(p#�2� 6��3 l� 
�r�Si���D��,З��0U2�0��"Q2�nlt�M�`��$*���f�~����u�N��|�pf���o���3mG##�_��)3	-8���|�|�����|i���9�k���d�����4�{��F���d�it
9�>��`���U�ي�@0�=��0�X���R!�*4@K�HT&
zu�DBR�CKC�n -x�#�N���;�;����}�Zv�y9'��-��>�,�����q)���oC�["�{��p�f�ES�������j����q���3�7Ϝ�v��W�g�n ȗ����g�ipl/�}����[7�x~�����{u�<I�_��<=�"Q��ދ|����`,4��5�tUs���ìL��?&L�Ⱥ�R�UA_�G �[�Խ�M�$���X� B�aJ�h
+��C��f`�u��R� T�vme�K1 �sl,4��`��JQ�3!����w^!��$��=H,KAʺ"Ʌ�(9D!D>=�X��`ll���_X>}��{gΌ�{�b� _.(�K�Li�h������>�y������=h�bX�~Lzݮm��z�^z_Tu&�8#�����	K�glN@�Z#��2��jEل��(�Z��Yʿ�8��ΒB�|���#��EQ�tx_^T�N�Y�c�ꏳ����^�}/Q�uI\�"�|�UP��9k}��
 
E�m��ؖ�RA����]Ǳ?>vl���������5U���� A�:P �WD������un��f���[�y�֭�6����Zs�j�� jgI����$KX����|D1���> � ��7�X�V����X�^�_����A4�$��C��{>��9!V��?���M2/k
*#�M����!�w�
$�kU�gB���,����k���n뚦,�>v�����Ϟޒgj�Sg �����)W��Sx@�e��ym�ƍ�߬���=�8���qoo��9�}"I"��%
}1�A��e�~�m@�GÉ2PT+v��:���_;PM<(�	��d����.���p�����0�P"�Dx�a�j2&h$fz�I�*F
��9)�a�i��a�͚S�4-�]�oLM��������\{a�֦�0C� _/(�k�r�^ׄ��?\����hd���;O��v;�y����t��I���4S�`�#�l՞�$�#�����h�"��d u��P���	e" �f����+�e�{4ܴf)�4ǜ���Q�p�
I�⢮�9�(��ȚѶt�P���F��v�,K�r�ݩ��OF���������	� ��uAq� E��>��q��qe��cs�`��������v�D���h*��1��Z��J�J�%"��]�&B��4����J ���@�� �T$|�_��b�O�`[b5K����"s1�d�iY�sA�rU�SYSc]3UU;�,�jVmۮ՟�굍�Fc��؟ԇ&�ǜ�;3#Ƣ8�<)�A�o(��iA��	(f�~����Z����[;pg�v[�;��I����n�7�U�H�`$�Z��zc��TγL�8�E�� �m��)���A�p���
P �E�/��R.IBNϠcQ��TQ�D���*���J-]Ӷ5�xb;��e��ѱ�F}�وS�n4��Ԕ�LLL�hN� �lP �7�ʪ���F�Px�I��ޞǾ�
�p�5���3�{^�u='�F�cQOdi�"o$YV���L�L˲La������<
�{B*v#D����$��51}i(�����+�R���C]�[�*�����ul�c5jm�vZV���O��R'����X� ���� A����)�,�0m�)!��PX_'b�)ݜ�^�i�~`$I�t<5H"�
5#5ˉ��LE�6�9��B�B&JR�(R&b,(Z��R�HJ�(j��Jd���v��1��($�����d��y���k����R߬<*`�ޭ~(�B ��{��Ow������?�s�9yA>� ��� AA�P � 2 �AA@q� � � (A �� � �8@Ad � ��� AA�P � 2 �AA@q� � � (A �� � �8@Ad � ��� AA�P � 2 �AA@q� � � (A�����}x    IEND�B`�PK
     eO�Z��[?:  ?:  /   images/b75f5fea-d559-4623-b1ce-f8cd504066c2.png�PNG

   IHDR   c   \   z�   	pHYs  �  ��+  9�IDATx��}xT���;��L&�B�P����&
F��"*�(MT@��T� H)ҤI��e�L�����������{AA�{��s�d&�Sֻ�Z���;l���/�������Cd��!����o�����B@�����b)0~:xrU��|�(5�����r$���������D�ر#|.�b�u���6}lZ="�����_
:LU��
�ӝ�P/�����:v����h��N�P�h)0�vN�/��vOK��oc�ׯn�߶��e�0��)�
6�R�5�K�ѯ_���+����ß���o�?�Z�N��z�&c9n��>�|>p�\���/�"2�O���x�S��4�y)B����]���`s&��T�A��P(��������-�C;d�4�Ñ�fee0ig3l&���3?��|�)<?��J���6�ߏ@0�-DQcB�_7�|'9�9�{-�|.a�Z!���W��$$G����n���p8���C��I�(���^��
L�:��ixa�Xl�q C�z(��C�KKuHO�7�a�nTUi����2�o��d;Z҂����Ph���\ZQs~��i��[z;v�u�7��O'��^�~�zr{�����s�.<��8�|�<9n,&lV�z
o]$ �y�}���ȉ-:vh�5j�$�8����Vt�\��QR�yΫ�4=�����s�E��+��Yѱ� �;p$�K/���g<����?��
0h��^�����+����B�j7�¹����;1~�?�8��X$�HHNN8��,.��Er��� ��1p�#}��A��	�\����(^~u��d�6�qV��ڵ�S|�d�:.qw^���fMs�@,^�^�5�Oa:+�؂��YN�A�9�E���b�蘘~=z�y��ɦ��7�
�u�����!�B(|��D�hߡ5$�wg�粚��������#�A���x^_������G�Ց�_G�ĭ�ܥ�����'�b���<���?��G/c������	Dx��W8�N{q@��#��}������S�9�x�X�0[Ⲉ�)��
M��K��y�,_.LL\���S��6f���£�����^g2 ��@bBBv��i|����'��1���+�=9vj����k��	�O�p0��ъ/ѵ{�3�_���?��3c
^��l��.'�����|.�"%��~-Ij%"�zE}K��#}$��)���=~⬠��2?R�Z�b1$a�� �$�<=�8>>q
�:._�"&.i)�`�C�Fm��}Fh�4{j�G�ݦC����ɹ3����?�ÉY��F~~����L��������]v3(�DH���C"�@&���(��[#IV&�EYZV��y�x\��'�'@��i�$%'V{=~_��<���DNz�����ı������V�EYyLf7jJzJ<�����+���'&O����S�<�O_����:z�����R��_yJ�T�^��2��TW�Y�V�fL�C] ��(eb��V�����0����sX�R*���%X��d�ec��?��ӗ!��^�`0u
Cc�d��'�BL|���A�vm�Z�y�t\Vx�
l�4m����)/ݚ����K��|z�d,[��Z�C����b�·Ah%�\�>�=2p��a[j77��6i�q�|���$���a?��?���WI�����0|У�w>X�O�pz,��� 3����I!F��qN�0�B���6m�1���6��d0.��~��BR\^�Ӆ�9�Y,���6�e�ƕӦ�  ~���������gL��P�C;�g�!<n�\��v��N��ӒѲe��6������w�&�y*xd�|��*xJ��OOf��/�ӭ[7��֓$φ��ۈ�{���S��n�����O�KĐh�ȡ���~ϑ��&.�(ùKWЮu�;Y�j�>nҤ�aÆ�ێފo7�è��>0_=P0h̝�>$2)�ݽ	zv\�v���Ԕ�b!"��@�G�]^+�g5�N���������?�5BSI�9wsޞ>��������"<N�-ě�|�N�a�E_ ��@z
���|吁=�>�jsrtT_����k�Ж� `�ի�2�F����~�h6�G>���
�W�C�V-�i�z�l��'���f��#aGB� �Sҡ��^���F��JV� ;8�?Z
yT�=]S-#��!�e�.��μ/ӯ�"��Е��E�������5[<z�?�!���J\�)F���,+V��j>9fTϋgι�|����z�/����xD����y<�VW�B�h @(Hoiݲ9�S���h�g%'�����6��=zv��w���	�"�D�T�f5� �LޚF@��L�/�8��CL"y�o�O�xj�䒊ʥ
�$�����(B}Sq�����]{_�TU,�}l�����&�����X�v��l.��t:?�h*��f���5��DBz#h�4'��G���7��j�e�7Y0�H���S��fQ� �������1�� ,�����m����6��?�p6b��v�-��t�:B���Rn~�w3�}�H�`�/�Za9Jo^CTl�6�%����~�D?�&'!�qKTTV_K�U<VVg$RC�^|�����hg�9��׷��'�N�"�3���B�9D��Yp�|ϟ>�<:�s���o�^w���r4�ʀ���d0�<y��	�ť��j��i�����Oǡ����6�Yo����!�w�����n�>SA��b��1j4k����j��K=QU�����c��S��>� <$M$#�$�.t� �'�g�=�����p ����Ek�.�R=����Q��~�V�
9�^�AÆ.;q��-�͎�m��S(9	�n�Q�k6t?�C�ˇ�_1�2T�2Η^z����W�������F��-�7�^��i��]x��A|�v#��3�PBZ��� �����gv�n�|<N��n�nrL�8A��*���p7	r'��NȢ{�-ry�kEvW�⊢'�S�B啕Od��C���8����ڔg�=r0a��_���0~��^�8r��\�C�h�ݭpXA���_�?�ʗ��6m]�E� I�zEI椁�y�Ӕϻv������B��C1�;t�8~��o�#�a]���� �#E�q�:{� �bb�V�g*����M̗�����!&	O!lt2ǝy&a\,.��Ψ�bΌ%��*o���I�B��z������<��_�{���k�w��vo��a����9p����YP���xm���gj*F��s�EQŤ�i�2� �� ���7��$O[�Tbwy���xg������l�
��' �p0��=H���@2[E?���=Ϥ��[��_�7@drLZ�`��ֲ��V$gL����Gz����c����l���y�f��ٹ˛kWm�����E"I&�'�����A��WbR�n���ȟ���{Og�աr���9
u�&]��tz���k�ӄ��N��;��1����˻n���uP�kў%D��wI�JR�5�E�z+��2��J�g	uN�+*����}��Y�-��Qs������ѫ��[�g��h-N�*�'ʫ _F��8�������nL�y/��t�B����W!�8Hv�׮}���iߍ¢���m�����jv~�a�gC_xi.���p?����":���_��_�|s��Xz��U]�
<;�1d��º5[�;�f���6���H�8���{�?�<i�e���/��h��a�`�^<q�ۊ�oU�z��*��jX/�3�.}7�ÖwO�v�h���X�VP��A�P�(�g�bQ�����zGX h����%�;��>�X<���$)�@`��'���`0,Y��¸�1a�H��k0h|��<�-o��W�����>yE��'1��q�Y�+?��`������� ��@v�&(�q뚏ϙ�c���v�틝I�_���oe�B�!�cԛ�\ۻ���dy�UEX��_��X|](�.Yd����e��Ayo���t�P^S�H���8���w��,�C,\����M,R~���3.>v��v�:�����,�sv3�<Ѽ���co�����iGii�ӓ�[���ټxq�&4�KD#�{�]��g��ѕZ�윋Y�?BN���s.��\���B	>�E(a&��#._pZ&�O�X�+ʞz�Ѥy�F��p�!`���[v�C�~R\f(����1�a��Z��I��5��{�]�{~P�H��J⻗0�J�����\�=�L��A���q���PD&�թO_W��+\6�q(��t:���[v�}�һa�6��k0�d�m�X0D���~��Ǣ����}�[�ǿ{��ea0����C{q~>�s�H,��eEt\*Jjo��.m~��X�ه��׋�D2ѳ�/���s8�� ް��Z=Xp� �����-խ�*L!O$��&��e�i�����9N3F�p!8�3��:��%Z�.�����9��٬S|�qz�EAtG�b(��/\,����}��]L7	���tw�CwY/�k/=�8F��CM<�n�������Ջ�r�������sH�c���tUDӖ��^x�'=ӊ��="	5@��|��u�/U�im ��C����Q��`S���Z	���m|��l���<��;��9���i����!��Hh���Ʋ� 5����L*�L'o���t���`�J�"�V����2{���N}���B�&�r�J1 !S�H�jZZ涱�W(���z������ɍ��8$�AzDZN1ذX��ϸI�	R.�����^�	�4��:�^�-&6�p�����Y����\�g�j��
��H�����V�fp��@��B���Ù������U�5iS�b���@g%ξ��?�����`��a1�iVTEZ����no���6	�[�qK���3_�nP� Wv������l���$r��]���OUE�U|gFyi���g<��=�2�}��ؔX&&-BjAe3Zh>��Qt�<����G���B���=�%(/���I��uQ'6����,�U$�*�q�ڵ�?<J����f^����H��Us �"/r�L8���jy�Lª� l����/<�㭡M1b喻~�L}���>,V�^*D6�Le����ܤ��I}����`&,L,�b�Y���¨�3�I����)����V�^$I
��j�������=�A��Tb��L:?�\��ߴ
/_���O�0�.��1t�����3mN\Nj���GKd*a�v�B���q�%�^�#H��aܩ�"����%���9� �y>���݁�9J�tĤ�Y����|c���V�ʅ賝�z��!�1*�zpH��^�\��[�|��v��*6�g�;KXə��O�bc�(�)�fjpP�p����.���m����rȜNɤ��ʗ'N���a���ta��z�����&�S��NԠ�~:L,y�c��a)!���i��u%�B$���n��u<��}�4#�cH|�8�{W���B�iS�V.�<Q��P�~�"�R\�Z�T&G#�ɂ ��x��:�:�$H}q�l["�%�?�|W��?EW�[�fx�A:��I�m�N��k���N�;G٭6��\�bb!��$&A��7ۭ�L(Zaq�F�^���~�m�K6~��P[c��ڽix�d\���a�������F	S�V�۸q�p-���Q6�S�$��h��K�!�ӑ�vI�Gn6��}�쿎e<!r��`x�$AK��	56�����c�x�Y:�M�`!���f�|uI^>��Ń]}��2��J�띞 %w���Ą�;�f��~,�g�#i�~Z �px��㓒od6ju��U��/7p&My�!�H2h�DE����e�Ux�Ib����>�'^_��C���{��^���[���!!3���T���W�%�h��m|bRo|�b-�N2���HX����Z?���{���>A!��R6J�1���2�b��c����d�$��իp�D�b��\��z�ǂC�"!��	j	I(2��*&��. ����	1�Z�t�ɚ����>��~�	�=��];B��/�����T��\�/z���ZÐaCw�LK���G�',�.���`0�oւPz�f��H��ۼi��O>_�_}�`���OhGϾ����lSC�i�ఄ[�`�wm;)I؄e��L*���3��\}�m	WxتT�R�~rU���*��B$e��R&W`�EZ��dXw�}��w]���j.܆J���Y-p���������B�a!�g�OP}sVke�{�m�g�X^�����^�YSU����'�#���uGu��u��П���e�>Cµ�>_������*��������	����alEyE]IE%2R��Qj���"��iq���ҝL�I
)�Fs,��IK�L*����[�;��H[w����^�(�}e��PO�4�
�x1f��@%bPmA]l��#��Bo�0U@SUb2m	X�)8�`���j�7�3H	�����M{n�F>��x匁`~s ��}�Ϙ���	�ш��˺��m�S�֭�8;d?"
£��p��.�� �m�Ʋ��z��0���B��`lIBUݕK����{c�G�!�q3Z�]��D�!	Z8x��T")�7tF	]rI	M%���b��]j���W�����Yj~�����i� �z�@���.9
�b���R=T���$I]�CuM�l&����h K_�̨u�+$a���)��Z����fU�tD����&b��ױ���'��k�.��E�,�A����!%)��`�;�{џ	)��Pg#�-��U�?1B�G��^*��={�۶zp`�P��?_�'an�8\"%��H���-��r��S���{�<�����fw��e7��1)�l��֑�e�^"���A+��]�pX�DX�4c{��V	��j	H�#I��U�^S��2���F&��vȢ�h���-��C4pPL�w����hHwiL[bd��i_l��e۾A��d��z#���g�S��p����v7�RZZ�z��&�,r?�������<���¨���/�IoR[���cG}�t�ŋ��*/�r�,g�T$Ngg�%����$z��p��$V�͌H�L�f�:Z-����a����'�ʆ�<,���4��2��'rW���n^~�R��LC�u5�z�jL���u\I�jx�lpzp�I�K�Í2+���L-��n�U��~J �8�@��(s��E��5�/�w�� 5-	b���a�L�q�]1��Uh	x�;H+b�L&KLzn�᣻��y�`�}sk�،��F��L�y���%E(�b�P��ls�j�����`�t�=��$�s^�Q�y͇�aH�����1c��O -}�s������._�XB��6�����CX1E�!�I���p"":2�4ي(l�v�!�B��Y���٢:$Hp
�IF�{c�$)����/��Q�X�X�5f�X:p��)4u�(:gPɠ�yv��Dȇ�Acb2�V�%����?Z��}�m�'����牸�P�$z҃|=����:���:���J|zx:HB��>��b��P?)�f}� ;ߺ�#H�� �b�bUR(�R�j�Йh�z�����ȄTIE4�R��+(�䐰(�U1c(����u�!�(ᗩ��"�!���.��x��h�����{z��o .J�����a�D�,.�������+a�p�l&�E�g�x�y1Ez�c�������Gyl~��v��Ji��wI�'ظB���op��;���� EE�hu������#���^��'b��<'	3V�J�]%�	)�F5�\�h!�qIⰻҊ��r!]eb-ը���Sh������8�ʊB)%���&�HhIQ
�e����x{`�����Z?�_�1J˫�-s�YI��b ������`%9Ҭ�#퉴b6�AQ���=E�{�{�N�YV��F\�]\Xh1�+c҄)Y�k���c+�C�_���@�Kh��t���pf�c��q��hk��F
!��wϕ���`��M�P�������Pcw�Q!�sB8\�MR���!$8�()+'N���������kG9ņ;Ć����Z�I\��d��a��=���:����RZ�<.�&����$����Oz�1Q�I�V�a>=�%�˙6=s��p�l3Ȥ�ͽ��Z-ƹ�ZL-xғ���Ϩu5�%�_�P7���Ev_1�py=N�R��Y�D�����	O'�:�sul|����"��DoAb�L)f�����v�� %�"�nGF��p~��|�r��p��+F�h��DX�[U(��0uV%��ѾqΛ����!�~R3���b���Gp��,�p�b�P����>�^j�l�rDGGB �x�n����j��E|<+�u�$���q��2.�|���qhra���f�^�7՗?t�MH�n�j*_�ی���њ#�#��	�)"w��jɊ��E�^���8�4�"��=�&�W}�����vo���]�Kk�:%B�"�M�V�v��b�,�"��0aN#�
uxQM�8!��:�j4�Y9�v�
�	
<>Qq�{���	љc�u�$��bG�7{��Gr%�[}�z�iL۸˟��/�u�scp� I�,f�Vo
���FD"�"��O���K�8BLn@LS����L��N���K~����j����^��w�)}��sbz�hi\�a<��.V䅠7�����K�GŢ����*��#g��l�|���ʼ���^��oﻈ-�N ]���m�A�\�vc����J0.;�a�Fl-g!M�ߪ!ɽ><U�E�  .*6?[��M���q�ԍY��C�9+NbK����R�ښ! ���"�����w�+sg���?kc0���;�$�ED�2�Q�6��Ee�m�B!M�J("�̓#'��I@�c?��*պ����l��":a�k�G+]�M=�g���PLf��:VmE��ÆǞ=�.��?�l��7�>�Z¤.iu+�G0�;'���˲��*�6 C��!�"�1�Z(ak|.l�W#c�p��Ʃ:�I���ѾQ���YV,���c%Xs�67��=Ukd�m,�������a�8r��͍��V6!.&ɕ!"��$iw��R\|�|fz0`��,�a���m����Alr�������k�R�b#[�z�g������ڠ���p��62R�tm��d�wr�=��|��:��:cю��lZDGj�l�r+c���ؖ� �nbI�j(]vp�n�#�a2����:��[0$#<��kнY#p�A��KH�n�!�r\�YPcwF���8����e��͛���yV�=�民|a%Ąh�-|~��j��M�0>�����)c��s��������|���5�Gx� �YsJZ�׺������<k��]�ǫ��c��Px�<Z���o ��za��w-�����鼯�y�Oc��Ukga���]���<�.c�Ydd4�Kc�Ir	Mq8��p����v�g�;+3�@�	���l*n�E�Fy��Ew�d��J�ޖ���Ȱ���hۋ8�� B��z>�YeӧLǶ/?�|bb� �,���)���bb�m���U �βUhٺ�QqkL���ZMmLbRb�/55ÅA�j��7�G�k�# �v�s5��=y����s�M-�������Ò�G�Ѯ��TW)�T���)-[�n���h�(A��$�"��zX�(ԣER�ݺ�a��лKgD�x�V����C &���&GR�f鞓V6s���o��Q�͛��|�7�_v�٧�N�#�;ag4|��l&��}�>��@(�+�ק{
����6$<v�wO��]`���)2�:Ԧ�g|VW[�fNl4"��\���P�A����jhh�:*�ź�s7�r\^祉�}}ܫC�❝�0{�&�5N�j"���ڶ�!�i�9Aɓ-El،NDŨ�L�}$�n.2�ӑ#A��
.����8"��������J�����=�A4��A�zx}��chܸY^��oD/����.x$G�X<o}����[����l�P �õ7N�>>�ۃ��ߖ+Ü7?A�.]����������J�RS�2��?3���}bqؿ��JMu%��-Pr�:�������O�x}6^|��_=���m���g����@��Vr��6W��&%#^�vXI\~�ȤP(���2��L>j+o�d�W����������{,3-�,Y-��S��~��=z���3g�����I�;�<2�<\K���n�<��Z���J�(u8]�a��Z�~'�������ٟ���}lAҒ%����1*.�MM�*�����f�t����/.+Fn~G�b��GΝ�����gK��������{`[���N"��)�$*g�yLo�2�R4$������B����ό�0�I� �1�w�bqI�O�I�8Z�)�ONI��o��`̰_���W�����p���}�UTԀ^��w%=C�VASW��ѾC)���D�D�XJ���Pώ�o^+�F�N�Fki��`�@,^�1��x�i�:v:�������LV��aalTt�VWy��ud�e-�z깦�����{��5F��3��b��^[H��VZ)�@�2	�.�Kf�$)�p�q٪H�� �q�����k56z�=Q��ڎ;	6�	m�r�3�&����0�R�PC/#�_�q{S��Oh����B���[��ЉX�F�k��}y_X�:�q��<�|���^�v֒���VEE��z���H@�s�����Q��W��O}��곯N�s�f����K[�sb�ݢ�����d��~��`���[T˳2�c���JtKSAt�����T�B�cK&�߾i�YP�cI���3}�|s
7/�_K�~��bB��6<�#�(����ʪ�=٩I��z�k<&��B� ,�u�RqŁv-���^8x��{��}�NT;�Ő^�h���v||�lMyɪ�7��,���.㬨�D��t���8�w����.���+���}�#~��m��~�C�C�[�X��qʡ��tO��*dX��2�HF�FrDHEfO���,�Kʆ�`��@�v���>�E��͛d��r�<B,�R�[r�n�V��d��Yb��<�9"ݒ������kX��ǿɏ�m�1Ĝ��)>,�����k�3Ԍ������bUuuȱ��P�aԵ\���v�@���k����=��_=���M@=���G� N�l��'���YCbUqߏH'�oWp�H�~bv�py��Ħ����	�б�^Fp�����bR��PH%O���6���* �����녫|��`�����(U�=�ñ=M��k�I�����&��u��>�����f �c��߮�<�l�v�UG���
<>�e%�NH��fa����C�6�/_�����|ه����J	c���_l�O�j�^/.�Z]c�s9wX��T�ǫ�e��l���h�+�q�wm{���'�AM�V�ע��J��J2ӓȽ��,)���`McJ��J(�bw8�������/������`$%���B���,���9m
n^<{��dDDF���
55��IH iU�S�?v������G�w�N��ק���󤅶����⛓�ݱڼ��5��ݿ��^�.a|�sPg>�z����~W��w�^�~�5��t@zR�c�Ed�у��++#��d�QTQ�d��ي��/J�"���x��t�<t`;��؋�?l�����;$t�k�/7����
ж}�ʸ��ᚢ��L{�R�@IE9R�Hr��̱�h�x��ė�����8� �����`�)��Z�;6��C�0q�*��e�j����𯘇���}�`l���y��{�����ܶ��QҪ��闯��du�ws L�**7<	��ǔ했��V���];��Ը0m�����-�| �U��K>�
������_��j<DSrc�,�s�l(+-AzF&# >Q�u�h�ǵ�_�����YPZQ����G`��I�>d��^kb�,>q	�:��c�6B%�mW�у�����s�W;p��Y�(��{��g��ӫ��۝N���@�Fo���6�3�DbQ�"�^@����dx���s�?�`�F���%x�h���������۔����
]���"**��tuLO�?s�]�Ur���/>0�[o�t�8���c�;K����&M�y7�6O���
*N����0d��<�-�"Z)�h��x~IEŔ ��
�f���*���l��O(�6�T*����l�h����;�̌HII��>{��M�@Lyi>>yo>���Ԭf�+�ontY��N(���������
Z�o��ux��{t�]&���å�����;����R��r�zt��+\=~���ź�����a�p��mrZ#/+��7�F��Q����M�8ಘК����p�ܣ7z���"�<��_0�1�~�������8y
���/�z����@�x�]|�h>a&�Ҷݻ�9��O+-���%�j둙�edj*K��3�4�����9]��=:t;(�J�&F�M���)�yS�Z�;w����E~~>�t�|�b��B�/W�����ؑ�z��,z�:�u��K����\
���GN���-�!&=�Jo�ŪU�6ꩻq0�#V�Ȕ*}� �e�Y��6��ӧb�s�譙��WȆ�,z����vlEy�mӥGkߡ�5O4�i��]D{4i���:��z܈P*@
���9=�t���y��E�}r���{gk"S��c!	����es�C��=����vPX\��_��~�����/خ{���˫���Aޕ�����#���cK�Oz��։�l�z�D*eӳz�@��/�Z�/�=������-��~�öR]4�l�q_��cƽ2[Lo�hs���()-k�GZx��l�T��X�&Q!�Ŗ8�d�ߟdw{�s���s���Z5oR�f���v����d�Xl]���()��U�D℈U���~�8�QA���œ^K��+y��z���W���+���O󤪮4� o���1c4���ƳS�`�'K��M���E�i=>��=�?������Ii�n4�NT�K[5�&4�!����^������N���fs�|���iL�3�<"��}��&^��.�/{�W��)T��=���A��O����t�8^����l�G��,�J�'����3�~ժ]��^8c�x�0f�� K������j��ۭ[Ǆ��Z����BZV�ki�Ysj*�>R)$hժN�	��ؘ(j���-Wy<n@���qY�(�S`19�%Bt��-'»�0~���
o�CQ�"�`�t���R H��dT�o��`�"%BxD��t�W�`pꅲ��O���::�|�շxvܨ�?mc�IG��v���wL[ޮ��&�n�Mj���۴�ɓ'��X!�K!+"�~_O�/`��e��{@=XW�BPLNIo��{@�D܇��g[�z&�]�b�ʢ"�u*��iu�F�]�,6'R��;�{$���yɆ�����^�zv�Bhj��Ѳ�ק��ɟ�/��ꎏW�����S3ߜ:o�Ј+W�k����;���'QW�I� �\!?��I�|�P �`ȯ�B�� ��C��,f(�f��&#����d68��4e��"�>3<�"n`�9.�@�G����ם@ѵ�ݷvo]>���`�o�{~�K?���y�7|��'��Y�x����ٙx�h��W�AWW��xLe|�PMB��K�2��P!V2���t�J8GЛz��X/J%����l�>xV8t1A����8��)��E;*���;�^��}f���%��n�^<��������G:`��}X��ۻ�}���';v\YXX�jl��٩u����פ���pz\,&3��f��O>�����;���]F���61��(br��
���J�<��P�;�Q��v����B<7}�i��5��9;6}����O��	��b���X��Z�=#x�Ծ�=��>Z�׼�7�lM�a���tgr|zC���`2km��f�Y~_4�w �����G~��yM��$�ELB��-�TǾ�w�Sߍ��Ѽu�kJ�`�����!�-�6�rpp��-���P�A��A}p��oU=����Ϝw|����77<�5U�<�R*E��i$C��/�����az˦7|w�֒0E1�,6�,O(Y����USY�8qx��p 7m�k�ǡI��a�ݺ��T<4`�֬ٝ�����P��?��X�Ƶ����f����l&}���(g�͈�9z���Vr� �i#ٸ���^�
����q'�|:�f�.�BV�۷~���|��6�jI�����=T`�b������װa�R�xqa��v���ן)�y
s������v�T>�����x^�Pd�GD6L�>M�<F�kߥ'�q������1������3�sfO��f%���C�߇<6�.�D�G�c��Q[[bt�lF_8<��ɚ�QtxrZ�X��
�Y�cF�Ɓ���4o�{��z�xh���ٶ�?����Z�_�П���C
�K���a�������`�_����?*�I�    IEND�B`�PK
     eO�Z�&�y`  y`  /   images/8c2f1315-cf23-4ba8-a920-becb97f13280.png�PNG

   IHDR  �  �   ��ߊ  NiCCPicc  (�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D�0գ ����d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c�%��V��h���ʢ��G`(�*x�%��(�30����s 8,�� Ě�30������n���~��@�\;b��'v$%�����)-����r�H�@=��i�F`yF'�{��Vc``����w�������w1P��y !e��?C    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs  %  %IR$�   tIME�WxG  �zTXtRaw profile type icc  8��S[n�0��)z^�8~$R��b;^eWݪ��HQb�0$|�>�� D�h`�dZ@�&F�Ąb�9��m��P=Eec������O8��`��Й�f�
�Q�A:���{�xt�k��7�����������-eP/���\!�����jS�u�mۃ��Qa;��B�["�,FدCl֤�	�����/�&�S�T�c��\���~�y�_���D6:J&�D�z����f5u�R�����Ye:�010�����?1:9�����{��5nH����^υZ�w�R��WU(5G�Ӫu2j�fo�-���)�:&c*+q�y&�"J��G��|/��d�c?&s&]����VG��^q���@����줁/0�   orNTϢw�  [5IDATx���w|e���3[�����!�XQ�	6�g׻��;�ӟ�SO�]�Slxީ��)6Գ��^C��m7����cӳ��؅|ޯ����y����S�y """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""�P �t뎇yX��s*�+��������L����>����<�r�ݵ/�ϯj>��ߌ�	�\51�;Z�w�e[�L�>��( ��R�	�NUo��W{��v��	댍
�_�f�|����Io[����7�9	s� W�>����&A����@��H��t@U���"^ n@U���^}z/[�j�[�*)9����n͚?VTV����� �*�, 4 ��{!��yLDDtX2�I�+�|���5]�dݸy����S�NMX�˯����^!"Z�SNDDDው�]8|�+LUU�S�
�n�u=&҉"""�����]bc�L������H'����ZND��fK�<�M��DDD p�ݚf���*(w��CDDD��%�$ϷX��'0���������p��a���ʓ<���#������	E��Qn������iӶ/[�lBaaAV�`�Դ48��vX�6�-fh�	�R�4J)(�L�O""":t��r�];���T�r:��'O�����z��:<7<O�����F�ۍ��*����v����"�_A��jf"��r�|��������Z�����=v�m����X5z4LZx�Ͱ�����QCrTAii)~[�+¹1k���e�E���;���^�&���� ""��:Z،m�tV��r�}^_��✕Nx�^�m�H�Q�6�5�_�6���At�z�^{�7].��#�WDDD������[u�ޤ�r9�q{"�F"""j����"b�-��t:]p{8�Q��JJK��x��.��o�\.x<,�E9�

�i*^=x@w��NDD��VPX �������}U�z<p�\�N'5C++)���r��~S�7}>*++#�F"""j� n��&"M����|��`@'""�f
�����D����>�,�E5AM	��������r��t:���(4��r� Ȉx>�N�3҉$""�������3ƌm��.�x��N%�������/ �y9�9Q���M������NDD�4 PJٍ�������(��@([�6t �z}0z������h 4��^�����(�i�ee����h�����(�iK�-W*D@�1�E=m����R�b� �Љ�����_�� t�"A��#""����+ �ϡ�ʝ��(�VZV��H�*w/D�H'����B�*�˕@LFx}>��NDD��VQY�D�Y�NDD����
��q@���;Q��*]N��!��%t�t""�h%М��J�u�h_u�8>�FDD��9�����_g/w""�h�UU���S�����G:�DDDdD��j5���~?K�DDDQK ��p�tݯCg�;Q4�b��b�W]t�)���(�i�����]��:QT�L���]ס�|
���(�i��LP�0��܉������2�fJ�r'""�j�)(���ua�;Q��bR
!:�܉���� �DD���ʝ��(�iգ�i0�OM�r'""�v͖�u]X�NDD��u*��^]B��܉����V=u��-�p`""��&uݸ�΁e������h~����*w""�����z���*w""��%���u%Ͷ���NDD�4�߯A� �+�C�)���(�i�߯��ϡE9i��5v�#""�~���J`\�.�NqDDD�N��	�)NNDD��l6[�����DDDQ�l65�`@oW�3[j^���&��Q ""#f��dX�~0�d������%سgv�؅��TTT������PJ�n�!11�������dt���D��@��!"�:��i!K�pr�V��"((,Ěu��ӏ?a�����ۊ����^�'��P�Q�4M�f��EJj*�w�#�c���5j��2a�4v":�(���fM�̡2N �ro!���b�ڵ���O���o�v�Z@��hI��� �z������ck�f,��������ӦM������b6��'�#�P\Z
�łX�#��9|Ĭ�BV�C�ϡ�I��x�d�R�=�m|�ɧض5��Q��V����TT�c�o��t����o�����_���{�]-��O7���������Wa�QG��f���x�� ��ZM�mݶ/�y�y��صk'�5�촭ܚ��-�7���Ǘ�č�wfL����/ 6j���m؀_|	�����xp�e�F:i�10�\�˄� ��n|��x�����Ͽ���"�U�&-��]��ۢ_񧫯��͛q�5� 1>�A����PXT�w�{���?�r�
��Gjj:T���d�B�*w�U����r�~�<��S((؏�L�Z���jVb��d�ɤA�4�������!�/�fK!��PX���gݏ��"�|�M蔖ƠNDQ������3�������rV�u!�a���|�8������x����sꝌ0�@n�� 33]�vEnn.�v���D���#&&�*������ �6m�m�6��
?Ȫ�ବ��g�����w/:��3�Q�Q �-[���x6oڈ��/��̀�B����F�}��nǿ��:�^�O�@�edfb�ر�:u
Ǝ���,$$$�j6n�p��(..ƪի��O�����c���5&������ks�"�S:��v8�vu"�:%�%ؿ?����p�Y X�6��҉G}���u��g��Ĥd�:}:���J�1	qq��6�|o�n�!+#Y�p�	���+0g��{�-��0�{=x���w�޸䒋�)~Y�(�(@)��ۋ �D��*wv������չs1�9�s��Q�����s�>��;	qquü����e�&3��G~�>�,r��G]{c
�Ņx���p�B��u ���B��.|l����7��ByY	�s�f2a���x��p��� !>�EA܈ ���p��31���2tx��jؼi#�{�y�UTD:눈�Q  ����]�*w���������];���t9M3��s��3�>��C��K ��f]O���z]�u�qI��g��o�e)�����.��8"�����ޚ��.@m$�q�L��Y�݋�99�3� �8�d���<1P(.*�K/����Bu"�#�D�5����EX�n^|�%���^��c�!�u�,������,7i.��bL�6-d������H��!!DBv3L�ڱK����[�0��<66�˵1l�!{LL $'&��+�D��0*�������?���9�te�:��}8��)R��ys$���~P`��f����+ ;v��']��(�O�<g�uVD��;f��8��S���/5M�����? /o+���m��������z�v���z f�6�V�f��v���G��4x?����|�=p{�����X,�Z��Y�0�L����zo��v��vCD`��`�X`�Xj�o��
��p������v�����������
Ku��6���������vC=��f��6��+_�Q�ן9p����z���`2�`�Xa�Ya�X`�~\���,=F�S�3: ������]�����f�ߚydMi��7"�^@��U�_�V�Z�S+1)_r1R����& 118k�x���QR\��H.5Kh8p� V�\�n�f��}{�b��X�n6oڄ�{������j�"..�ѣ����!''16[�>����rTVV6���dBJr2̍���/,Ě5k�d�lX��w�Fee%|>lV���е[W���#F�@�~����Т������k�d��[�{���鄈��p >>9�9:|��>�{#.6���T^Q�����u��vj����dX-���+*.����d�R�[�;w�Dee%�^o���ƢKv6r��b�0` R��[�6���k׮��ŋ�n�:�ڵ�������|��CVV6C�A߾}���|iN�M� (-+�֭[�v�Z�[�۷oGA~>\UU�z�0�͈�ۑ����]����4p z�쁄��v�ٯ��BIii��RHLH�#&&h^Wy<عs'V�\�իVa˖-�?�W�~�V�������Fnn.�����#==�6/Z���N���w�Ʉ��"��_]�QPX�������M�w8HHH`MBCR�C�r�ϡ+ e��OPU�Q�|���8��qM�Q�0t�|��(�!.>���ӷ/��!C�b�ر�r�]\R�_~]�O?�?��3�mۆ��2��kf�b��%;cǎ��iSq��ǣszzuN���:^y�U��ƛ��PA�Ν�ēO�wϞJ8�v��ǟ|�w�}�V�DaaQ��P0���ԩF�9
^x!N9eb��pj��{�|��gx�w�b�
VO��SV��;w±��/��=��9�Σw�}s^x���"���D<���Z�DFM��8����s���;X�t)
��k���43R��0b�\p��6m*R���-��������罍%K��� ��x;�iiiw�Ѹ���a' 1!�uU�G[�m���_�/���e�q����\}�j��l�Թ3����S�`ҤSЭk�6��*����#f�{����T�Z����o���hpL�UU���_���a���c�8++�)�dAJr2�)S�bƌ��ۧL��>��~̞�>��chZu�Q@iI	����$)�����nGBBB���u]�̙3q���T�� 6�M3�y)���7����DDV�Z%�{��~��i��Vy⩧#�?~]�9/�,g�s������g�Ɇ�����\��{Ӷ��p:�O>���8S��S덑�Ο��T����䤓O���������9�~�����������EV�ZU�Ϊ*y���O�-���XgBb�\vŕ�a㦠i�r{��O?�'�$�Vn'5-]���u�c��V��?�4_�R�����+���RN�<Ebbb[��������s�=_��\ix.y|>���2����kU�$&%˥�_!6mn���{��ǟ��#F��jk��^w�[m12�����?�)

DD�_�jm��x�z�.���9/6ȓ�k��5��t�Y/]-���"�ǞxR��燝��W.�����_8�9���Z<^o�cġ��������W�$&&�Đaß�L����y#�+R���_��ax�euɑ��GE���n�t��oi�t���߸Q�t�%%-�A<�">1I.��R� ~@��_��[��A�dw���V��H~a��q�ݒ�֩Z�~e�&�,�W�j��""%ee���K猬�������-r��dͺu�:���w�(ej���4��O?զ��G�̬�6c%���c�ʏ���$_*�Ny��$�k�6oGi&9a�I�h�v;�}~�|�ͷ2q�d�Z�m<v�C{L��v�Y���E��5�|s޼ꛮ���ify�ŗD�����s5zL�s�m�`���9�] �6l+�=^�\z��횏W]�'��}��|������?Q������UW�)DfBN>e�E]���b�����o����
���ߖ� �9J>��3���%��^�F��W]]�d�%��N�m;vH������n�#��n~�9���d߁�KG���Y�����n�Y���z��q�v���|)���{�%	���S&O����IgU��0�E�V�V.� ��<΁�,���x}�V�Y$t@����""��[�k���u��)S��漼f�π~hzBb��'���) ���X�|E��4�5
I���3\8�o+]�	���j����h�2�>�'PJ�j��j�C�����߭²%���k����~��#L{�R
%�������˯�����뽤�>5�9�K�����|�p&�y��g�tVɳ�o磏>ċ/�����������O<�gf?ge�i�k�O_Kҫ���O=�J�n��=�O<��#(+-#���?�v���k<��l���V���³�<�[n�۷�ե�����Vs�����f��>��Ar���5����Ǜo��nǲ�O?���|vl�Z�/�Ϥ���`�5T�����<���t����ԍe�7z�����c��
�Z.ս�Us1��d^}���طo���v���T����	۟17�p#�6oBM�4���cࠁ9r��� %%�����{����e˰r�J�߿��3X�sN��my����a��q�駵S/V�߇���:�x����n>�c��ХK6z��.�]�*W�����u�VT��:F*�~/��70}�t�\�
�̞�*���vLGl<r��W�^HOOG||<\.v�؉u��a���՝Ϥ�qW������8���o{GB����x�w�rU6�?&�YY��ݻr�� !!n�شi�l1�	@M�2����8��3P\\�G~�����=Ɓ��������HLH�����]��~�z�ܱ>��4źߋyo��̙31n�Q-��χ�^~�f݇Ғ"��:�q�ӧ/F��A�!5-q��p�\(,,D^^.\�u�֡���^fԧa��������O?��G�^�+��+V��9/4� p��!;�z�쉴�t$&&����@����!o�����=�7?�}�]L�>S&�2=�z���Q��i��z�oټ~_��ٌ�}� !>�i�8�ѣG�ꎀTK <d�ˡ�ܭ�yu�kQW�|�_""��J�R�� ��]��E�qy#"�l�
>rt3U=��N��?]#��^�
���Kc~]���b��_�o7��dee7S=	�?`����/-�[�*wM�[u�w���b���㏑'gϖ�+WIqI��=��|��z���R6m�,�ϙ#Æ�Y�e2Yd��iҳw�F���O��N?S�xk�lشY�+*l���T/]&��q���t�?&�U~��v�r�+P��0_Lf��5Z|�Y�t�KU��V�\��m�����2n�1�4S��*M�Lr�Ie����|Qu�㈓I������%kׯ�����RZ^.+V��Y�= �z�}�(��|�m���Z|ο�����_�?q����k�u��r�%��'���?�DN;��z�����������q��R&INN���uHjZ'9��d������������|�t�d�Ν��G˹�/�	I�^�:�).-5L�_MP����{���={e���7ߒ��� �TIrr�����o���g�����҈_'U��_­rOHZ��C��2�[��ʫs����楗_��fx"6\v��uD午HQq��w��m<�����O?�J���bj�""UOu��)�e����8M���v��
����j����Y��n�^�{<�>Էd�r9���͗���ӷ����\)*.iv;^�O���2h�Аy3ᤓ���(�1
���%1)E���FٴeK���˺d��[��$�kwyj�3�?���|��|���d̸�C�ˈQ�e���a狈���;��ԴN��{�!���m�\�����By��g�i�V2��0��)bЛSM4�E�?a�|��gRVQ��^RV&/��buڍ:�)霑)?���;��_~)���Azjj�|���I(��VFe@4x����^y��d`mF����;���I��������W_{Mb�/�J3ɔi�ʪ�k[��""�����s����Dd�G{\���N��E(K^z�U��x������V��s�ꐡ�F�7�~>��|�駒��E�j��v�!�W�{��z]�$����O>U{�nz��Xz����Ss���ǟ��脻��� =z�6؎�������~{��*�\w��B��Kv��2�5qU��[r�麼�����|�8y�ŗZ�
��,\��?ʖ�[�F���뺼��[ҩ�q����Ly��k�9�u>~u������8�����C-�˴��T]�;ŉ�����:nt��	�6�m��{�⥗^FeE�&��0�$<���n� �z����>���f���
��}6nl�����o���a�X��p���>}zXKgfu�=��N8����:e�D�v�ü)(����[�-W �l�⪫��UW���E�2b�p�}��P���>�)�����1c���Z0@� 8��8�����PRR�6��>�ſ�ݷ߁H��i�Ĥ�~���a�Z[tk�z1)�3�8<� :gd��5E���ܹs�s׮��Li�y�L�ݤQ�^����:�L\r�%PZ�c�������QYY����tPi����,p�W����LJr2,Cf����,]�zZ������v+���ݦ�5;��~+����k׮Ň~�E('�|.��RX�ՊI�&!>>�B���p�e�a�)���ՊSN����S�*T���eK{tcǍ��W�16[���I�p�ĉHMKCs=��=�\�}��V.��a�ē���t;^��7o�?���U�|�-�޽��wM3���/�%_sn<�	�g�v���
��֠��t�̟�em�ӑ��7�x:��55�%i�Z,8��sеk�n�桰��]RM��iF�]�H������^�Fb�#��eYE>��C��A߷Xm�����;���_#G��u�]�#�.c�ߋO>����k��� .>]t�SS[�@VV�/�:�v놙3ς�ln�vrs�"-=x��u?���ۜ#5�b����.@���V��O�>�޽[�|t��s�;���k �ٳ'��2�#(..��o�͛7�/�2X�����_	GLL���V��^z	�`�tw��~�	J��ڥ��4Κ9�n�q�>}0d�P��K��Q^V����@4MӚ-��,�+ >�����餶�>o޼K/1XBG߾}q�9g7���-���N��#G���5�VW����_�~?��6�%=-�YY!�9���ѿ�6m'%9ii��RQQVI4�|�ޣ;&L8�MkINJBN׮!�3f���)�@bB:w�l�LEE�z�!�����m��tn2Yp���!77�ݚ�@�=0��i�M���8�&��֩SgL�2fMk�Ͱ �����`�[e����+���n�t́et�������v�M�h�"�ݻ���5�<q"zT�õ�ѹ3N�~�aUdYY~���v	^�G�F�N��Plv;:g�يѣG���>�ݎ��$�������|�0�aÆ!��s`�X���a���0rԨ�Y�ZC!0�_rrJ�|q���1�� 2?��#��`������ĉk�@m/&MÄ	�����7������Ö�����>�+jJ�k׮0����|>����5���DS��b��9}��d��zz�`D�6�Jm�>�-[fp�$��`ʔɭjwn�0q����%���t,Y�eeem*i��V4���`2�[=�i��JHH@�v���b� 6�a����m��3�L8hP��6[B�4����h�a�Á�i�@����.��y�73���}��r�*���>}z�)�F��h���<X��o��xڼ�A�!11��n�SRS`���	H?����%���xU��HE�{ȥ������
@iY6n�h��]�tA�~�Z�w��}���m�6��o�1z����j�����$''#�Kv۷c���tٶ2��j��w�^mi�v�a����ѭ[ז��`;m팚��{��Q�����Ў��� �d�\ߴiS�o^�2�W�ۯ1..��fXD���F��@��r�4MCL��4�i��RXX��;w�߳WO����l����ܾF���cZ;w�j�V���;����iƗ۸��fn��N��:m�v:��m�-�)���X8���(_��~õ%/�e���f�w�.��c��{�n0��ٻg/���߆���vdfd�9��X���ۤ@��TbVJi!�H��J)$��#T�����6�5�G�����W��Ē����؃�̽�d�`2Yj'f���҉��m�F|\<�����q8���9 �)�@�MHH8��c�=D3V������m[�3���Lطw��vA�� JKK���ڪPR\��6m�j�"9%�]�n6��B��v�8m��T�w��)�.���Lf�����t�x��hTPPgee��Lf3����Ih�tɂ�b����$
~���-�;b�i�bs����j|��������l�Z�'���<��~ط��MK�^�O<�8fϞ��-Q�݆�U�ۍ�¶t����G����6��A%f���n ''6�.��N���p:�H	��pQVVVݩ��~
L��z ����d[Uմ)C�u������j6[`1�@��:%��c2���RZ��mP <^o�APD�(5M����P\ܶAZ4�`��5��2�B���9�+ ddd">DUdQQ
�x'-�n�a�f2��#�Q݋�)A��m�Ř�&�ڱ�Б�d2�|�^�V^OscL ����+8]U����J)��C7k��nGm��f�~�m� ������xRTT���o�]�K�1w�*@����]v����9�`>��M碦��E�p�iLGؘ
���>x=��E�"At�vxl�:i��;�q��;���O߾�FGZ�fmTݙn����+QT\]��(Tk���_�W����Y��Pe{�T�����zЎ���@�����G��e�h~������.���?�Ƞ���ʕ+�t���=�����SO>�?���r1l�0�9@NN`2��f����_�QYQ����r��	>8��4�cbjg�"j��M���x���;�<s�O6�f2�K�.�%:�����r��G:��� �>qqq�(����+�}�h���ښ�����_�k�v�ڵ�|���t��@��}0b��u֙8jԨ&�)���i@��������"�t�������QS�z���1��!+���s_������f�s�7� $�znC���#'�+֭]��]Î۱h�t X�~=���P����ʅ���}[�[���郣F�j�ل��m6Tx=h�Ș�������������mSi�Z?8P=�Պ�x�N�U.bc�پ��&�D-��U�!���`����wW�������rE�u֯��n�w().F「�1�2220|����OMI5|F���b���}�m;vT�����l6dtj��̨c3��HO7��N���E����$�/��f[:n@ v��'MBl\��f�-X�e˗G,�
��m��駟AĨ3�`��a�ݫW�w�;�W�����P�t���ׇ���A׃����S�N=/��g�n�6S���;w�t2�ZLucu,��ƌ9
��r��$�iؽk7��{��ko��9֭]���M�7[l�x�)HLH�SSS��c<�Hޖ-(*j�`F�Ôb��͆�$%%��8�D�޽z�f��������o���\�լ1��҉�&��Ն�1�_��.]0i�$(ͨ׫�?��.\tȿ�
���7�xOU]���G�8���1!!}g�Rؽk76���v۶m���[`ti�ѣRSSbNRGҳW/���� ��%%%��}�Y_޶mX�b�nۆ��b������ܩMj&
���a�4�}�L������ְs�v<��c؟�Ⱦ�
�����9/b�0�7�0u�T���ǰm�j6c��Q�XlA�TTT�/�����m��W_c�޽~:j>b���ٶH�{�n�e8߹���k�j��v�n�Tŷ�z�N��3N�g���/�7��x��G�漷QTT��N-"�hh�U�w�*w0h�@�y֙P���_|�^xa\n�!�2~��Wx��W��U������9g�k3�{�1�32��E�W_}��۶��) �������/t�}���aԨ����$
� HMI��1c�&X�����7o�m�/���|�}{�`������x��yx��'q��7�GCE���!Ҵc�:v��b"�Й���z���O���SO>��^zn���u���q���`�>��- e�̙ga��ͮ�o�>}�h�w5l\���|�8� ���ϰl�2�}���aÆ�ܤ�Ƥi8�	HI1�Y�g�~�%K����X��t����7
���!��W`KcƎAff��L&4��XE�9�zˉ&�t�:�s�u�(�_����fw x9�������栢��u��E���K/��=�����/���)^@B\�O�{L�q�=�*<������e����Vᩧ�Fee��{�2aڴi���>�/pth�5
�F�B���a�x��Ǳw��6������W_ᓏ?6\2>!	'Nl�6�H��Ï��5d��i�pJ�S �Ʉ�.��N��C��� ?���|˭؜��n]m�n���G��O�`ѯ��X� 6.��_0hР���ĉ'W_��ض5�� �mk�>) ���C=�իV!xէ��ݻaƌ�T��UM��y�Gl�:�}��'x�٨t�~������u������� F�Q����C�{q$�ڬ0�-���'����9�L��@zj*n����ۯ?�= �P^V���'.��b�2�5�;�ߪ�^���<�}�?p�����K~�6�L8��p޹���, ���p饗��Y澜?7�p#6l�ܪ���k��r�mx��wO0�ɂ/�C�a��iӦ�㏇ѹ��z�ܳ����BQ+{�+z��q�X��Q�UABb2.��rtJK��{�#6[�!x<-Z���΁-��7�_¶�z�����u'2�d�8�+躎_�	�^s-.�݅x~΋X�n=���-�����+1��q��s��#�"����8�N��[n����P�8�t̘1��}]��>�5�_/X �����Ѷj������E���ÿ_��M����
Ǝ�+.�V���$ux�SZ���/��2�.+����ч�M7݌�k�A�0�58�u]���~ß��>��Ð���S&c�ē#�-�L\|b�1�
�}�̛7e�+~]���g���>_�8?3�M)�}��pV:q�m�#��>�zd��t⛯��?���ݻ㨣�°�Cѯ_dee������NTVVb��}X�b%�/[��K�b��mգ�5׏Q0v�8<���գG��� HIN7ހ�k�b�eA�MAD��W_a��u8��p�93�۷/����҉-y[�чa�k�a떼�u5��[�����н{�QZ�șp≸��k0��Y�r9���T��rᕗ_������/�ӦMC�n]g0\���
y[����c�ܹؼqS��<t����IhR������aÆ`�*�ٳ��z����0` ���PU�B~~�?����Zx�_C 1�|�fo6}>�9��!��_|�Ep{<���b��=]j���x�i�zlڸo�a���@bR�6t�\.8�NT�������P�a��`�1������#Z}����1�Y����my0z�g��]x��G��o`���}�hdee!55&MCaQ��ۇ�K�b���عc'�~o�}ё��	����4q�8�ԁ	 �ł���
�v��K/�T�hӠ.��5�W��nǜ9s0|�p�1�3����Ʉ��r�ܹ+W��o�-�֭���y�|�;�#G�0�Y��=z��g�T���G���>� Ji���ǟp".���%%u�<�����}3j�\���
t��	��+VT�*�_l]�QQQ���2��j*��i�-VL;�T�{�=<p`���S�L���p�-�`[�u���;�g�N|�駰X,�X-PJ�������DGVv�����.�I��e��N �$%���^��z�MA�^/�lڈ-�6��wޅ�j��b�����v�ü��93w�uN�1#�W&ҙq��l;v,�5>�a�� O[ri��(,,DrRR�w#z����yUs����eO� j��̳��+�����<�����	��^��=	w������sϴ[0 M�0s�Y�={6F��y>�h�u.��ge%*+*��x�*ԅ-��!C��SO��/�����ړ �����܇��+���{\s><n*+*QYQ��*Wu�i�|��={��G��W\���!��I�N��aC�5 
�����H'?�h��;����Ç���O>�����b�"p��|\�q�2�T���+���;�����[Ӕ©S���W_��.��	�a�W��*���HLJ�e�_��_g�y&,&Z��[�P�+�j:��}�]x��'0t�(MC�`��@5�K�|���<�T�y�E��y��ͭ;އ��.L�s󭷠KvW�$�WTT`ǎ�ޅhn:zs@��4�����)���{������5kQ\T���Z�խ���̒�����1c������ɓjs9XGH <�<3�'O�+���E�����%ψ��GRr
�=�X\tх�4i��ڶ�n<�t�i��� ����4���vj�_�01�N��K]�������X�����¬�z��rI��o�V@lL.��b�;��}|��6o����=?Z�y��5�����_r1.��|dt�Ԧ�]D�=��ů��~=	<�l{��ߪ���f̀���+W���>_+ۨ�ra˖�����ݙux]g@oV�i�='���:\x��X�r%���{���ö��P\T��e0�w0
���I�ջƍ;�L:�F�DjJ2���
s�p��c�ē��w���>ǢE�k�.8t�N�̈��C�^�0��q�2e
�9f<��{���S
�9�2tX�1�u���ܾ0�ZYj����l2��HW�_G��}`j�H_�@�G��1x�Ph����޽{u	�y�6|x�s]ב��[��v���:lx��뺎~���j��b��(���9��_�ѫWO�Z]�S�f@n.f��\x���������`��U(�/���Fs%Jbbc��)Ç����N�	'��ݻäT����d6UUU. "���T8z�V||���Ғ��/8b㐐�ت�6�L�y֙0` ޚ����%��塬��6�( J�`�48bc�������sЩ:�2��w�ݳ;+��_r)^x�y�m6��@M��"(,,Į]��c�l޼�7oF~~>�N'\�@�v��M�`�ِ��Դ4dgg#77����ӻR��`�>�#u,j����Ǝ;�n�:�^�[�n���P^V��
����@\\,233�77���b�����̄�:��~�ʊ
8�Π�[,$&%Ak�ޝ��p��o�j�"!!�p���G���vv����\�W�t���"�{f�III��p�Dee%*&1�-HJJl�픗���r}/��I+_�Q����Rlٲ�ׯ�ڵ�k׮�w��n���!6.q��HLLD�޽1`�@���=�wG|\��;߫�n����=�4�II�߱���xQVVt\�a����M!P�p�@>��m�Ν�p����N@)���!11	����YY����n{}D�_�7<�ԓh�&4&&f����ڳo���P���]��^z1v;z+��]A���x<�z��z���|��|Д����
{LlVk��F��g���������J�l6�b�"�no�6~����/w{m�p����hَ�6u ^�.�^�70��R�X,�Z��Z�������<8X�>(��ߏd-�fa�! ��o�4���p���~���9�4>#�&���b�u����3�Ѳ�m* V�VKBȠ}0��<8�ېF?��z���ЯlCoo��k?�N^�)ԑ�|?��kᡦ��|	��:Q4-�����p�""��$ 4�ërg	���(J�Hӧ2�E9	���e�8""�(&�.͏3�6t""�������Q4-�����:�E�:�5_B�u�����(-�)�D�˝���;���0¿�h�DDD�>�.��V��0�E%DCm�::QTif��z2�E-�$�6tv�#""�Zv/wщ���VJ��DDDQIDD����Љ����ha������(���;#:Q4����3�E)��{�����(j�7�+{�E��&g�s�DDD�K­rg	���(��`�5��E��̶�Q0"��Љ��� ����ֈ���Z�Я�U���;Q��yl��`�XNDD�D��|l���(���Y�NDD�D���NDDtؓ�Oe('""�ja��V�E�0��Y�NDD���ǡ_����[���8�+Q���H�����Ba�;��#�8Rё ���,�E�p��YB'""�b��rg	����c,�j-X�����Vؽ�Չ���V���Y�NDD�X�NDDt`Fu""��ő∈���2s""�(��ʝ����NqDDD�?ζFDDt�p,w""�#B�m��DDD�,��eX�NDD�Z0�E+�GDDt��ќ��(J���;�Љ���Xx%t�r""��֒��։���T�c�3�E%�!"":"�߆.�r'""�V�V�3�E��*�棵��E��c��Z�)�����Yx%t�C'""�R�oF��Z5�ADDD�R-��>s8K�u���()-�����C�D:J!���h]ס (��4�]���������*�]�+@s�	���jE������U�HD�Q�y����>x<(M�b��d6!PFm�밴�����ػ{ws�U���J ��W�1J�DDD�C!�[�* W�߆v�'""�B���Eo""�Ù���G:%DDD�j���tJ�����t@y5�ie�N	�� ���v��H�����ZGӴ����2-%%�q�Ų������#�aK)����φ��F@Ff�q���wy<�" ���j�U�{N�p0:�%@��iͶ�����pD�g?��������9ETM)��R�V��}gm\�a�:����F�~�w��ի��2"V f��b���1&�ɪ�4��4��4�R�T��`B৪��R5WE�T��k�U�f�.�PX�v����RhxW����x9.����R�<\(T�]�R��ԀR����u�V���o5�k���^�=�:Z���Y�~Ԧ���������j��d}J��u�������4��Z��p�	��ʂޠ��^��u��c�o�5��b�x��/=��WD�H�����9��:{�~���������nHBi�{ͪ��R�4����k?���F��w���'��f�!��`geI��5�|M^�~�������4�	��t�cP��V�p��Vw\��n�f�'�z}���`����~i�'|�P������e��e��FK׻�68�W� ۯ9$���dݵ��p����u?t����������K�Y_��]�j�GR/���\�dX �5ikt\��*e�R�p��I�ɋz���ͯ?��ڹ};�~x�W��]��E��O�����FGT},�4��o
 �t]����߯ ݯ+]~�_��D �_W��t%"�~��s��oP՗]��^W�i� ՜ "�7H"XMŊ��>���]���>k��כ����}{��m�9��g���_y�7���4������]�78�J)���x���q�I'��^O���_��5oIݽj��O ��V��b��Ҡ���"5�RR�����R��$5W��;_���U_���BW_]�҅�r��ȁ?���M��r��7�R����d����/U�=}��Li��i
J��MдڿiJA�(/nKE�c}+M� Д��Ai�mk�Mi  ���;�ݨ�j�,��Q{JNIE~�<�쫇q1� ��)[�fʼ^�}>8u14��4��~�AY4(� ~?4ѠC�I5z�_�h�P ���\����k�R
���5��=�j���5�^[k�ª��5�)S��/uWߠ�cG��ɧLz������-���+��s�|6��0٘PRZ��n�/��r�������#F�87--}魷��ߏ�1���d�l����&��-W�ƥd�hT�Qu�T����7��n+�ꭣ�i�h=5�u ́�Oլ\I��������R��ڂQuU��K����[����_�D�N�	�ʹ�p`E���Hmy]�4����P��nOS
�i]��L�u@��lF �X`����*������t�	�v#..J)j|����Kv6X/�y	&�����D|B��v�G�7p9�� Æ��m;v���."�Ꟈ�����?"1�Xi����*���?�㳟�[��E�05�ک���L8�$�������M�Pغu֮] Hk�a꣏?�?���`��������'���Y看��6�sύtr����w��w��[o뒙���a���Lr�=�8"J�""�,\$	tMh��q�ۏ=q¸�YY�>,DD�XB��23�0c�i11��A?.\��Ҳút� l۱w�u֬^��_	������~�o����[o�S�<�$ŀNA���`��1n�ñ�d2]f͚�ض}[���j
@IY|�!|��Wh�p�RSS�>��c^�~��k�N\w�5�N6Q����[t꜉�cƞc�����ݭ�ye��ڎq������#�=.��xi��O�ظ���=�8�#.҇���Y,�SP����٫���7[,֢`�x�.��˯p{�	�>��3<��cpV��q��d6{323������7�Ήtr��Bb@���:�����:u�e�Z����l�2���V��
��U�qｳ�o�n4�(�����G5�I���6nğ��C��MDD�:�>����k猬7��t����N���?6��""���Η���ILL���#G���8"}���ڮ� ��={�]��A���d�'��}��*�G�w��l1A��M&�;;��"���.�sϽ�>DDaa�;��q���d6W[���b��%�r��j�O?��>�,�n����aC_7�Xٳg���H'��(,�d���>Đ��Щs�-��Ш}���8����T�n~߬�p`�^;��11�srr������G�?yB��MDD�>f�s..�������_�UQJRR���oDm���ȁ����f��٭[ϫ����/��F�����EXB��F�����,��>0�}c
%%%X�|y��j�������G|�}�)$%'�w������S&cǎ���D:�DDD�G����?`Ѝ&�E^�����rE])]D��>�N�A�i4��KX5���t���&"":8���[d�tØqGO���F}��a�u���	���`�|�J>r�a0�X�e}r�] ��}���NpDDt�:u��8�̳�&$&m1z=)9U��u������!�͕f����go����s��_o�!�YMD�jlC�f%�$#77woLL���K(���bٲe�Njuj �׋�_��?�F���0��~�j���x��"�t""���G���={?��I����9�|�p:#^Jy��s�vs��Q0hȰ �~c,X�l&"":�j:�6��f��g�"[�n�h@�����#Gs��������w?��r���]wϊt|_|���O�p��Wh�<zbb������v��ϛ����u�ge�?�x�4qR������й�Kq�Eg''��
�5Q�$�=�`Ăys���8�v�=�x(3���"�Ý9�	��CRb"����6
���˖.���D�ÁC*?��x���vW!�8�f�ٓ�����E��p�ݳP�*�R���DD�c/w
Kf�,\q٥����U�f|ڬ]���8�iS V�]������A�`��BrJ��G;��S�L����x��q.E�� �KF�;�j����GOLJ���y���ED
���/(�v󸸄���3<�s& ��>�t�z_|�N�p��:}P|B��P��<��#�$���x�^y��G�k�nn������� j6Q#�#��),�'O�裎����8�-'�K�.���:$����xꩧQ�D��vMӐ����i�Ϙw���`���8��#��DDD�ܜ� "Z�^}�`f�a������^3N���e���>o�IbRʢ�&��k��!����,$":hXB����J���V��f=�R
�v�Ė͛Z:4 %eex��G��/���4���]�u���W_nY�|n��o��B""���>j,N�xʉ�ظ�6kM3�#�=~�J�^�_�|z�8b���M&��[���������\�;�~O������s����GϞ���o����묬L��^ݎB��ޮϣ+ �}�=�x�	8+��txD��Qc�z殿�����>�L�����(z<�������]�u��xxUȰ�#dێ�ZJ�ۺUN8�$�vsh��m��㏱�c  o��v�����(��߸ 0pА�4�,Fϣ����7�k��."RVQ!�\�g1ޮ&��շ_������{���#�eDD�;�Q��ر		IHNN^n�Z���R(--��+�m�~��ƛ�׿^����oUӐ�)��S&M�{�Y3e�M����t�E��3N�̳�����ۨS ��K�UU��R���?�$��䆬jOLJYq�)����,"":�XB���������p�n�ܚ�kPPXئm) ;w��}�fa�0|D�n/�޽�_9͇}�����HgQt{� "澹�_2`FIZz'��ZUB�W��t����ILf�a�\3Y�n�{>�ҫsmW��Z<=��HgQ��UU �3�:�ŦZ��*��}��U�~y��Krr�W�k�����3g��3���0y�4�qNDD����
#G�i�Θ�P���+/UO�K�""�M�����=c�>�d �DDD-u�5��ڿ\ףS�����Qc�ɞ���.�׌Ӿg�>�q�!K��͓�o�-"��v�x���"�-DD�Nq�*��;��O��!�U۾}�n��z�*��>�>����S
��>�0�9g�9S߱s'�v�u��""���[�[3���&�%T)Z��R����󎤥wY:OLJ�8q�Q�9�  �/�t�~D=z���i��pĹC{՟�������V����G�l7����G��= |2�K����HgQ�qrj�-[�`��G#..n���(v:+;U��^���%蜞f8Q��_X��+�-�Qk��i�ҥ�[����7F��5�V�9-*Q�=��l�~{���[��qY]rdђ%!����̺���cBV�wꜱ����;�����@���������7ބ��G�>�ߡ&j��b���n�ED>������jW���P|܉���7��>�t����{ ��S��d�;ĸ]�u��M�>_�`�f�:9j̸����M<t�c?.��z�?f��g8�9Q��vƙ��UW����^���ēN�����t�������J偗R&�ֽ���xc��睏��^�]'"":r�����Y���G��ޣ׶P=�kwY�|E�������ǟ�G\�vs%)�i�Κy�$ p�uk�ϵQ��v~[�,��1�~0�r��~�?�Ou����_~%9]���jWb���{�	w��魷����|�]&"":򔔕AD���N�b��hG�t��]���{ٴe�{�	!{�k&�<􋧞y���7܈y$һKDDtd��変�\i��xC��%3N?CV�['��j1�X6;���k�������W����G��Y����}��l��\@��8d����h��<!1�s����$"�_~����#��DDDG�5k� �Sgddgǚ��OB�������Ymr�	'~4��S�}�y�:�_��M""�#ߥ� ���z�����u�׀���=����:�\ �眈��8q�46�;>#>!��s%�]���DD��nl޶-һGDD�q|�� ���g���[��f�L�>��=���~��7X�zu�w����c���7��~������̬�ו2�8��cbw�vƙ�fv���v""�����G{܈ظ��-
�J�9b���õ֦�:>�/һBDD�1=?w.�="��=z]g2[��	��"i靾0hp����b��a��""��������N8��8-)!1�悹R&;n�޻��Ǥc�;"ªv""�H[�`  ����{7[�뫫ԃt�-��w]|��h�N'�{��H���o��S�L �쎋�L%]w8�^�<uZ����GT:��N:���@$%�"%5�j����i�FU��j?5�Sv�,t��k6l�t�����1�dA�Ι8pprFf������Ė����LIM�ӳOߞv� p��wG:�DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDG���Nþ�C   xeXIfMM *                  J       R(       �i       Z       �      �    �      o�           ����   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��    IEND�B`�PK
     eO�Z�����  �  /   images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.png�PNG

   IHDR   d   d   p�T   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     eO�ZYQ���  ��                   cirkitFile.jsonPK 
     eO�Z                        �  jsons/PK 
     eO�Z�o�r*  *               2�  jsons/user_defined.jsonPK 
     eO�Z                        l  images/PK 
     eO�Z~`�	� � /             �  images/5de4bec6-ccea-4571-acb8-2cf876e4e4fc.pngPK 
     eO�ZN�ɴ<  <  /             �� images/f4826ebb-d8ab-4c3e-8d6e-ffd2265d28af.pngPK 
     eO�Zj���� �� /             P images/3281a32a-bb08-42cb-a591-9481e2c9eb0d.pngPK 
     eO�Z��I2\k  \k  /             @� images/35c60fd9-1fb3-48b8-b3d7-7968b0279531.pngPK 
     eO�Z	��} } /             �S images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     eO�Zd��   �   /             H�	 images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
     eO�Z�Xw�s� s� /              �	 images/49baae61-cb81-429b-96a1-6cfb8f124b59.pngPK 
     eO�Z��X��&  �&  /             �� images/9c69fbd4-c376-47ca-8b4c-793dd402431a.pngPK 
     eO�Z�Lz��L �L /             � images/256658b1-ffe9-46c3-9f0b-70052a8fe00d.pngPK 
     eO�Z9?B��  �  /             �� images/d18021d8-4522-4af4-a3c6-358ee97fa8ad.pngPK 
     eO�Z���*6 *6 /             3 images/a1588c66-a70c-44df-b30c-55fdbd854069.pngPK 
     eO�ZIRP4#  4#  /             �P images/2dd92824-eee5-446a-82e5-cb3be823b6e8.pngPK 
     eO�Z�IQ�H� H� /             +t images/a05d3615-68b8-4f26-98d6-1aedf7f6d878.pngPK 
     eO�Z��[?:  ?:  /             �T images/b75f5fea-d559-4623-b1ce-f8cd504066c2.pngPK 
     eO�Z�&�y`  y`  /             L� images/8c2f1315-cf23-4ba8-a920-becb97f13280.pngPK 
     eO�Z�����  �  /             � images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.pngPK      �  L   